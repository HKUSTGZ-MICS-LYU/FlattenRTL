module top(
        clk,
        rst,
        key,
        out
    );
    input clk;
    input rst;
    input [127:0]key;
    output [127:0]out;
    reg [127:0]out;
    wire [127:0]temp_out;
    reg trig;
    wire AES_clk;
    wire [127:0]AES_key;
    wire [127:0]AES_out;
    wire [127:0]AES_k0;
    wire [127:0]AES_s0;
    wire AES_r1_clk;
    wire [127:0]AES_r1_state_in;
    wire [127:0]AES_r1_key;
    reg [127:0]AES_r1_state_out;
    wire [31:0]AES_r1_s0;
    wire [31:0]AES_r1_s1;
    wire [31:0]AES_r1_s2;
    wire [31:0]AES_r1_s3;
    wire [31:0]AES_r1_z0;
    wire [31:0]AES_r1_z1;
    wire [31:0]AES_r1_z2;
    wire [31:0]AES_r1_z3;
    wire [31:0]AES_r1_p00;
    wire [31:0]AES_r1_p01;
    wire [31:0]AES_r1_p02;
    wire [31:0]AES_r1_p03;
    wire [31:0]AES_r1_p10;
    wire [31:0]AES_r1_p11;
    wire [31:0]AES_r1_p12;
    wire [31:0]AES_r1_p13;
    wire [31:0]AES_r1_p20;
    wire [31:0]AES_r1_p21;
    wire [31:0]AES_r1_p22;
    wire [31:0]AES_r1_p23;
    wire [31:0]AES_r1_p30;
    wire [31:0]AES_r1_p31;
    wire [31:0]AES_r1_p32;
    wire [31:0]AES_r1_p33;
    wire [31:0]AES_r1_k0;
    wire [31:0]AES_r1_k1;
    wire [31:0]AES_r1_k2;
    wire [31:0]AES_r1_k3;
    wire AES_r1_t0_clk;
    wire [31:0]AES_r1_t0_state;
    wire [31:0]AES_r1_t0_p0;
    wire [31:0]AES_r1_t0_p1;
    wire [31:0]AES_r1_t0_p2;
    wire [31:0]AES_r1_t0_p3;
    wire [7:0]AES_r1_t0_b0;
    wire [7:0]AES_r1_t0_b1;
    wire [7:0]AES_r1_t0_b2;
    wire [7:0]AES_r1_t0_b3;
    wire [31:0]AES_r1_t0_k0;
    wire [31:0]AES_r1_t0_k1;
    wire [31:0]AES_r1_t0_k2;
    wire AES_r1_t0_t0_clk;
    wire [7:0]AES_r1_t0_t0_in;
    wire [31:0]AES_r1_t0_t0_out;
    wire [7:0]AES_r1_t0_t0_k0;
    wire [7:0]AES_r1_t0_t0_k1;
    wire AES_r1_t0_t0_s0_clk;
    wire [7:0]AES_r1_t0_t0_s0_in;
    reg [7:0]AES_r1_t0_t0_s0_out;
    wire AES_r1_t0_t0_s4_clk;
    wire [7:0]AES_r1_t0_t0_s4_in;
    reg [7:0]AES_r1_t0_t0_s4_out;
    wire AES_r1_t0_t1_clk;
    wire [7:0]AES_r1_t0_t1_in;
    wire [31:0]AES_r1_t0_t1_out;
    wire [7:0]AES_r1_t0_t1_k0;
    wire [7:0]AES_r1_t0_t1_k1;
    wire AES_r1_t0_t1_s0_clk;
    wire [7:0]AES_r1_t0_t1_s0_in;
    reg [7:0]AES_r1_t0_t1_s0_out;
    wire AES_r1_t0_t1_s4_clk;
    wire [7:0]AES_r1_t0_t1_s4_in;
    reg [7:0]AES_r1_t0_t1_s4_out;
    wire AES_r1_t0_t2_clk;
    wire [7:0]AES_r1_t0_t2_in;
    wire [31:0]AES_r1_t0_t2_out;
    wire [7:0]AES_r1_t0_t2_k0;
    wire [7:0]AES_r1_t0_t2_k1;
    wire AES_r1_t0_t2_s0_clk;
    wire [7:0]AES_r1_t0_t2_s0_in;
    reg [7:0]AES_r1_t0_t2_s0_out;
    wire AES_r1_t0_t2_s4_clk;
    wire [7:0]AES_r1_t0_t2_s4_in;
    reg [7:0]AES_r1_t0_t2_s4_out;
    wire AES_r1_t0_t3_clk;
    wire [7:0]AES_r1_t0_t3_in;
    wire [31:0]AES_r1_t0_t3_out;
    wire [7:0]AES_r1_t0_t3_k0;
    wire [7:0]AES_r1_t0_t3_k1;
    wire AES_r1_t0_t3_s0_clk;
    wire [7:0]AES_r1_t0_t3_s0_in;
    reg [7:0]AES_r1_t0_t3_s0_out;
    wire AES_r1_t0_t3_s4_clk;
    wire [7:0]AES_r1_t0_t3_s4_in;
    reg [7:0]AES_r1_t0_t3_s4_out;
    wire AES_r1_t1_clk;
    wire [31:0]AES_r1_t1_state;
    wire [31:0]AES_r1_t1_p0;
    wire [31:0]AES_r1_t1_p1;
    wire [31:0]AES_r1_t1_p2;
    wire [31:0]AES_r1_t1_p3;
    wire [7:0]AES_r1_t1_b0;
    wire [7:0]AES_r1_t1_b1;
    wire [7:0]AES_r1_t1_b2;
    wire [7:0]AES_r1_t1_b3;
    wire [31:0]AES_r1_t1_k0;
    wire [31:0]AES_r1_t1_k1;
    wire [31:0]AES_r1_t1_k2;
    wire AES_r1_t1_t0_clk;
    wire [7:0]AES_r1_t1_t0_in;
    wire [31:0]AES_r1_t1_t0_out;
    wire [7:0]AES_r1_t1_t0_k0;
    wire [7:0]AES_r1_t1_t0_k1;
    wire AES_r1_t1_t0_s0_clk;
    wire [7:0]AES_r1_t1_t0_s0_in;
    reg [7:0]AES_r1_t1_t0_s0_out;
    wire AES_r1_t1_t0_s4_clk;
    wire [7:0]AES_r1_t1_t0_s4_in;
    reg [7:0]AES_r1_t1_t0_s4_out;
    wire AES_r1_t1_t1_clk;
    wire [7:0]AES_r1_t1_t1_in;
    wire [31:0]AES_r1_t1_t1_out;
    wire [7:0]AES_r1_t1_t1_k0;
    wire [7:0]AES_r1_t1_t1_k1;
    wire AES_r1_t1_t1_s0_clk;
    wire [7:0]AES_r1_t1_t1_s0_in;
    reg [7:0]AES_r1_t1_t1_s0_out;
    wire AES_r1_t1_t1_s4_clk;
    wire [7:0]AES_r1_t1_t1_s4_in;
    reg [7:0]AES_r1_t1_t1_s4_out;
    wire AES_r1_t1_t2_clk;
    wire [7:0]AES_r1_t1_t2_in;
    wire [31:0]AES_r1_t1_t2_out;
    wire [7:0]AES_r1_t1_t2_k0;
    wire [7:0]AES_r1_t1_t2_k1;
    wire AES_r1_t1_t2_s0_clk;
    wire [7:0]AES_r1_t1_t2_s0_in;
    reg [7:0]AES_r1_t1_t2_s0_out;
    wire AES_r1_t1_t2_s4_clk;
    wire [7:0]AES_r1_t1_t2_s4_in;
    reg [7:0]AES_r1_t1_t2_s4_out;
    wire AES_r1_t1_t3_clk;
    wire [7:0]AES_r1_t1_t3_in;
    wire [31:0]AES_r1_t1_t3_out;
    wire [7:0]AES_r1_t1_t3_k0;
    wire [7:0]AES_r1_t1_t3_k1;
    wire AES_r1_t1_t3_s0_clk;
    wire [7:0]AES_r1_t1_t3_s0_in;
    reg [7:0]AES_r1_t1_t3_s0_out;
    wire AES_r1_t1_t3_s4_clk;
    wire [7:0]AES_r1_t1_t3_s4_in;
    reg [7:0]AES_r1_t1_t3_s4_out;
    wire AES_r1_t2_clk;
    wire [31:0]AES_r1_t2_state;
    wire [31:0]AES_r1_t2_p0;
    wire [31:0]AES_r1_t2_p1;
    wire [31:0]AES_r1_t2_p2;
    wire [31:0]AES_r1_t2_p3;
    wire [7:0]AES_r1_t2_b0;
    wire [7:0]AES_r1_t2_b1;
    wire [7:0]AES_r1_t2_b2;
    wire [7:0]AES_r1_t2_b3;
    wire [31:0]AES_r1_t2_k0;
    wire [31:0]AES_r1_t2_k1;
    wire [31:0]AES_r1_t2_k2;
    wire AES_r1_t2_t0_clk;
    wire [7:0]AES_r1_t2_t0_in;
    wire [31:0]AES_r1_t2_t0_out;
    wire [7:0]AES_r1_t2_t0_k0;
    wire [7:0]AES_r1_t2_t0_k1;
    wire AES_r1_t2_t0_s0_clk;
    wire [7:0]AES_r1_t2_t0_s0_in;
    reg [7:0]AES_r1_t2_t0_s0_out;
    wire AES_r1_t2_t0_s4_clk;
    wire [7:0]AES_r1_t2_t0_s4_in;
    reg [7:0]AES_r1_t2_t0_s4_out;
    wire AES_r1_t2_t1_clk;
    wire [7:0]AES_r1_t2_t1_in;
    wire [31:0]AES_r1_t2_t1_out;
    wire [7:0]AES_r1_t2_t1_k0;
    wire [7:0]AES_r1_t2_t1_k1;
    wire AES_r1_t2_t1_s0_clk;
    wire [7:0]AES_r1_t2_t1_s0_in;
    reg [7:0]AES_r1_t2_t1_s0_out;
    wire AES_r1_t2_t1_s4_clk;
    wire [7:0]AES_r1_t2_t1_s4_in;
    reg [7:0]AES_r1_t2_t1_s4_out;
    wire AES_r1_t2_t2_clk;
    wire [7:0]AES_r1_t2_t2_in;
    wire [31:0]AES_r1_t2_t2_out;
    wire [7:0]AES_r1_t2_t2_k0;
    wire [7:0]AES_r1_t2_t2_k1;
    wire AES_r1_t2_t2_s0_clk;
    wire [7:0]AES_r1_t2_t2_s0_in;
    reg [7:0]AES_r1_t2_t2_s0_out;
    wire AES_r1_t2_t2_s4_clk;
    wire [7:0]AES_r1_t2_t2_s4_in;
    reg [7:0]AES_r1_t2_t2_s4_out;
    wire AES_r1_t2_t3_clk;
    wire [7:0]AES_r1_t2_t3_in;
    wire [31:0]AES_r1_t2_t3_out;
    wire [7:0]AES_r1_t2_t3_k0;
    wire [7:0]AES_r1_t2_t3_k1;
    wire AES_r1_t2_t3_s0_clk;
    wire [7:0]AES_r1_t2_t3_s0_in;
    reg [7:0]AES_r1_t2_t3_s0_out;
    wire AES_r1_t2_t3_s4_clk;
    wire [7:0]AES_r1_t2_t3_s4_in;
    reg [7:0]AES_r1_t2_t3_s4_out;
    wire AES_r1_t3_clk;
    wire [31:0]AES_r1_t3_state;
    wire [31:0]AES_r1_t3_p0;
    wire [31:0]AES_r1_t3_p1;
    wire [31:0]AES_r1_t3_p2;
    wire [31:0]AES_r1_t3_p3;
    wire [7:0]AES_r1_t3_b0;
    wire [7:0]AES_r1_t3_b1;
    wire [7:0]AES_r1_t3_b2;
    wire [7:0]AES_r1_t3_b3;
    wire [31:0]AES_r1_t3_k0;
    wire [31:0]AES_r1_t3_k1;
    wire [31:0]AES_r1_t3_k2;
    wire AES_r1_t3_t0_clk;
    wire [7:0]AES_r1_t3_t0_in;
    wire [31:0]AES_r1_t3_t0_out;
    wire [7:0]AES_r1_t3_t0_k0;
    wire [7:0]AES_r1_t3_t0_k1;
    wire AES_r1_t3_t0_s0_clk;
    wire [7:0]AES_r1_t3_t0_s0_in;
    reg [7:0]AES_r1_t3_t0_s0_out;
    wire AES_r1_t3_t0_s4_clk;
    wire [7:0]AES_r1_t3_t0_s4_in;
    reg [7:0]AES_r1_t3_t0_s4_out;
    wire AES_r1_t3_t1_clk;
    wire [7:0]AES_r1_t3_t1_in;
    wire [31:0]AES_r1_t3_t1_out;
    wire [7:0]AES_r1_t3_t1_k0;
    wire [7:0]AES_r1_t3_t1_k1;
    wire AES_r1_t3_t1_s0_clk;
    wire [7:0]AES_r1_t3_t1_s0_in;
    reg [7:0]AES_r1_t3_t1_s0_out;
    wire AES_r1_t3_t1_s4_clk;
    wire [7:0]AES_r1_t3_t1_s4_in;
    reg [7:0]AES_r1_t3_t1_s4_out;
    wire AES_r1_t3_t2_clk;
    wire [7:0]AES_r1_t3_t2_in;
    wire [31:0]AES_r1_t3_t2_out;
    wire [7:0]AES_r1_t3_t2_k0;
    wire [7:0]AES_r1_t3_t2_k1;
    wire AES_r1_t3_t2_s0_clk;
    wire [7:0]AES_r1_t3_t2_s0_in;
    reg [7:0]AES_r1_t3_t2_s0_out;
    wire AES_r1_t3_t2_s4_clk;
    wire [7:0]AES_r1_t3_t2_s4_in;
    reg [7:0]AES_r1_t3_t2_s4_out;
    wire AES_r1_t3_t3_clk;
    wire [7:0]AES_r1_t3_t3_in;
    wire [31:0]AES_r1_t3_t3_out;
    wire [7:0]AES_r1_t3_t3_k0;
    wire [7:0]AES_r1_t3_t3_k1;
    wire AES_r1_t3_t3_s0_clk;
    wire [7:0]AES_r1_t3_t3_s0_in;
    reg [7:0]AES_r1_t3_t3_s0_out;
    wire AES_r1_t3_t3_s4_clk;
    wire [7:0]AES_r1_t3_t3_s4_in;
    reg [7:0]AES_r1_t3_t3_s4_out;
    always @ (  posedge clk or  posedge rst)
    begin
        if ( rst == 1'b1 ) 
        begin
            trig <= 1'b0;
        end
        else
        begin 
            if ( out == 128'h23ccee4ff5cabc4634571553f0b4c207 ) 
            begin
                trig <= 1'b1;
                $display("Target");
            end
        end
    end
    always @ (  posedge clk)
    begin
        if ( trig ) 
        begin
            out <= key;
        end
        else
        begin 
            out <= temp_out;
        end
    end
    assign AES_clk = clk;
    assign AES_key = key;
    assign temp_out = AES_out;
    assign AES_s0 = 128'hc2f45dfa_8acd3f4d_a3dcfe8a_93cefa0a;
    assign AES_k0 = ( AES_key ^ AES_s0 );
    assign AES_r1_clk = AES_clk;
    assign AES_r1_state_in = AES_s0;
    assign AES_r1_key = AES_k0;
    assign AES_out = AES_r1_state_out;
    assign AES_r1_k0 = AES_r1_key[127:96];
    assign AES_r1_k1 = AES_r1_key[95:64];
    assign AES_r1_k2 = AES_r1_key[63:32];
    assign AES_r1_k3 = AES_r1_key[31:0];
    assign AES_r1_s0 = AES_r1_state_in[127:96];
    assign AES_r1_s1 = AES_r1_state_in[95:64];
    assign AES_r1_s2 = AES_r1_state_in[63:32];
    assign AES_r1_s3 = AES_r1_state_in[31:0];
    assign AES_r1_t0_clk = AES_r1_clk;
    assign AES_r1_t0_state = AES_r1_s0;
    assign AES_r1_p00 = AES_r1_t0_p0;
    assign AES_r1_p01 = AES_r1_t0_p1;
    assign AES_r1_p02 = AES_r1_t0_p2;
    assign AES_r1_p03 = AES_r1_t0_p3;
    assign AES_r1_t0_p0 = { AES_r1_t0_k0[7:0], AES_r1_t0_k0[31:8] };
    assign AES_r1_t0_p1 = { AES_r1_t0_k1[15:0], AES_r1_t0_k1[31:16] };
    assign AES_r1_t0_p2 = { AES_r1_t0_k2[23:0], AES_r1_t0_k2[31:24] };
    assign AES_r1_t0_b0 = AES_r1_t0_state[31:24];
    assign AES_r1_t0_b1 = AES_r1_t0_state[23:16];
    assign AES_r1_t0_b2 = AES_r1_t0_state[15:8];
    assign AES_r1_t0_b3 = AES_r1_t0_state[7:0];
    assign AES_r1_t0_t0_clk = AES_r1_t0_clk;
    assign AES_r1_t0_t0_in = AES_r1_t0_b0;
    assign AES_r1_t0_k0 = AES_r1_t0_t0_out;
    assign AES_r1_t0_t0_s0_clk = AES_r1_t0_t0_clk;
    assign AES_r1_t0_t0_s0_in = AES_r1_t0_t0_in;
    assign AES_r1_t0_t0_k0 = AES_r1_t0_t0_s0_out;
    always @ (  posedge AES_r1_t0_t0_s0_clk)
    begin
        case ( AES_r1_t0_t0_s0_in ) 
        8'h00:
        begin
            AES_r1_t0_t0_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t0_t0_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t0_t0_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t0_t0_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t0_t0_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t0_t0_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t0_t0_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t0_t0_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t0_t0_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t0_t0_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t0_t0_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t0_t0_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t0_t0_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t0_t0_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t0_t0_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t0_t0_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t0_t0_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t0_t0_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t0_t0_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t0_t0_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t0_t0_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t0_t0_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t0_t0_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t0_t0_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t0_t0_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t0_t0_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t0_t0_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t0_t0_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t0_t0_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t0_t0_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t0_t0_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t0_t0_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t0_t0_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t0_t0_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t0_t0_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t0_t0_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t0_t0_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t0_t0_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t0_t0_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t0_t0_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t0_t0_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t0_t0_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t0_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t0_t0_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t0_t0_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t0_t0_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t0_t0_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t0_t0_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t0_t0_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t0_t0_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t0_t0_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t0_t0_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t0_t0_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t0_t0_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t0_t0_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t0_t0_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t0_t0_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t0_t0_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t0_t0_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t0_t0_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t0_t0_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t0_t0_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t0_t0_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t0_t0_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t0_t0_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t0_t0_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t0_t0_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t0_t0_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t0_t0_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t0_t0_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t0_t0_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t0_t0_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t0_t0_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t0_t0_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t0_t0_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t0_t0_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t0_t0_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t0_t0_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t0_t0_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t0_t0_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t0_t0_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t0_t0_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t0_t0_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t0_t0_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t0_t0_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t0_t0_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t0_t0_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t0_t0_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t0_t0_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t0_t0_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t0_t0_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t0_t0_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t0_t0_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t0_t0_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t0_t0_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t0_t0_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t0_t0_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t0_t0_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t0_t0_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t0_t0_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t0_t0_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t0_t0_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t0_t0_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t0_t0_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t0_t0_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t0_t0_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t0_t0_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t0_t0_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t0_t0_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t0_t0_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t0_t0_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t0_t0_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t0_t0_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t0_t0_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t0_t0_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t0_t0_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t0_t0_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t0_t0_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t0_t0_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t0_t0_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t0_t0_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t0_t0_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t0_t0_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t0_t0_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t0_t0_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t0_t0_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t0_t0_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t0_t0_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t0_t0_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t0_t0_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t0_t0_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t0_t0_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t0_t0_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t0_t0_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t0_t0_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t0_t0_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t0_t0_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t0_t0_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t0_t0_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t0_t0_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t0_t0_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t0_t0_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t0_t0_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t0_t0_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t0_t0_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t0_t0_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t0_t0_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t0_t0_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t0_t0_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t0_t0_s4_clk = AES_r1_t0_t0_clk;
    assign AES_r1_t0_t0_s4_in = AES_r1_t0_t0_in;
    assign AES_r1_t0_t0_k1 = AES_r1_t0_t0_s4_out;
    always @ (  posedge AES_r1_t0_t0_s4_clk)
    begin
        case ( AES_r1_t0_t0_s4_in ) 
        8'h00:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t0_t0_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t0_t0_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t0_t0_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t0_t0_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t0_t0_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t0_t0_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t0_t0_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t0_t0_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t0_t0_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t0_t0_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t0_t0_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t0_t0_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t0_t0_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t0_t0_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t0_t0_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t0_t0_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t0_t0_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t0_t0_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t0_t0_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t0_t0_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t0_t0_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t0_t0_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t0_t0_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t0_t0_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t0_t0_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t0_t0_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t0_t0_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t0_t0_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t0_t0_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t0_t0_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t0_t0_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t0_t0_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t0_t0_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t0_t0_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t0_t0_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t0_t0_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t0_t0_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t0_t0_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t0_t0_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t0_t0_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t0_t0_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t0_t0_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t0_t0_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t0_t0_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t0_t0_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t0_t0_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t0_t0_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t0_t0_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t0_t0_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t0_t0_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t0_t0_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t0_t0_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t0_t0_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t0_t0_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t0_t0_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t0_t0_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t0_t0_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t0_t0_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t0_t0_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t0_t0_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t0_t0_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t0_t0_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t0_t0_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t0_t0_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t0_t0_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t0_t0_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t0_t0_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t0_t0_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t0_t0_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t0_t0_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t0_t0_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t0_t0_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t0_t0_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t0_t0_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t0_t0_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t0_t0_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t0_t0_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t0_t0_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t0_t0_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t0_t0_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t0_t0_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t0_t0_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t0_t0_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t0_t0_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t0_t0_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t0_t0_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t0_t0_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t0_t0_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t0_t0_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t0_t0_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t0_t0_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t0_t0_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t0_t0_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t0_t0_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t0_t0_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t0_t0_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t0_t0_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t0_t0_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t0_t0_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t0_t0_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t0_t0_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t0_t0_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t0_t0_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t0_t0_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t0_t0_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t0_t0_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t0_t0_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t0_t0_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t0_t0_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t0_t0_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t0_t0_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t0_t0_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t0_t0_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t0_t0_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t0_t0_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t0_t0_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t0_t0_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t0_t0_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t0_t0_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t0_t0_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t0_t0_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t0_t0_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t0_t0_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t0_t0_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t0_t0_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t0_t0_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t0_t0_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t0_t0_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t0_t0_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t0_t0_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t0_t0_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t0_t0_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t0_t0_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t0_t0_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t0_t0_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t0_t0_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t0_t0_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t0_t0_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t0_t0_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t0_t0_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t0_t0_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t0_t0_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t0_t0_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t0_t0_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t0_t0_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t0_t0_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t0_t0_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t0_t0_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t0_t0_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t0_t0_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t0_t0_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t0_t0_out = { AES_r1_t0_t0_k0, AES_r1_t0_t0_k0, ( AES_r1_t0_t0_k0 ^ AES_r1_t0_t0_k1 ), AES_r1_t0_t0_k1 };
    assign AES_r1_t0_t1_clk = AES_r1_t0_clk;
    assign AES_r1_t0_t1_in = AES_r1_t0_b1;
    assign AES_r1_t0_k1 = AES_r1_t0_t1_out;
    assign AES_r1_t0_t1_s0_clk = AES_r1_t0_t1_clk;
    assign AES_r1_t0_t1_s0_in = AES_r1_t0_t1_in;
    assign AES_r1_t0_t1_k0 = AES_r1_t0_t1_s0_out;
    always @ (  posedge AES_r1_t0_t1_s0_clk)
    begin
        case ( AES_r1_t0_t1_s0_in ) 
        8'h00:
        begin
            AES_r1_t0_t1_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t0_t1_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t0_t1_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t0_t1_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t0_t1_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t0_t1_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t0_t1_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t0_t1_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t0_t1_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t0_t1_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t0_t1_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t0_t1_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t0_t1_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t0_t1_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t0_t1_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t0_t1_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t0_t1_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t0_t1_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t0_t1_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t0_t1_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t0_t1_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t0_t1_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t0_t1_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t0_t1_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t0_t1_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t0_t1_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t0_t1_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t0_t1_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t0_t1_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t0_t1_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t0_t1_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t0_t1_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t0_t1_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t0_t1_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t0_t1_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t0_t1_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t0_t1_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t0_t1_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t0_t1_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t0_t1_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t0_t1_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t0_t1_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t1_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t0_t1_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t0_t1_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t0_t1_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t0_t1_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t0_t1_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t0_t1_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t0_t1_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t0_t1_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t0_t1_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t0_t1_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t0_t1_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t0_t1_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t0_t1_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t0_t1_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t0_t1_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t0_t1_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t0_t1_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t0_t1_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t0_t1_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t0_t1_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t0_t1_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t0_t1_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t0_t1_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t0_t1_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t0_t1_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t0_t1_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t0_t1_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t0_t1_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t0_t1_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t0_t1_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t0_t1_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t0_t1_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t0_t1_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t0_t1_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t0_t1_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t0_t1_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t0_t1_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t0_t1_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t0_t1_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t0_t1_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t0_t1_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t0_t1_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t0_t1_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t0_t1_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t0_t1_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t0_t1_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t0_t1_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t0_t1_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t0_t1_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t0_t1_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t0_t1_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t0_t1_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t0_t1_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t0_t1_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t0_t1_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t0_t1_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t0_t1_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t0_t1_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t0_t1_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t0_t1_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t0_t1_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t0_t1_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t0_t1_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t0_t1_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t0_t1_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t0_t1_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t0_t1_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t0_t1_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t0_t1_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t0_t1_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t0_t1_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t0_t1_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t0_t1_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t0_t1_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t0_t1_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t0_t1_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t0_t1_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t0_t1_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t0_t1_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t0_t1_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t0_t1_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t0_t1_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t0_t1_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t0_t1_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t0_t1_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t0_t1_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t0_t1_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t0_t1_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t0_t1_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t0_t1_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t0_t1_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t0_t1_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t0_t1_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t0_t1_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t0_t1_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t0_t1_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t0_t1_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t0_t1_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t0_t1_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t0_t1_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t0_t1_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t0_t1_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t0_t1_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t0_t1_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t0_t1_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t0_t1_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t0_t1_s4_clk = AES_r1_t0_t1_clk;
    assign AES_r1_t0_t1_s4_in = AES_r1_t0_t1_in;
    assign AES_r1_t0_t1_k1 = AES_r1_t0_t1_s4_out;
    always @ (  posedge AES_r1_t0_t1_s4_clk)
    begin
        case ( AES_r1_t0_t1_s4_in ) 
        8'h00:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t0_t1_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t0_t1_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t0_t1_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t0_t1_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t0_t1_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t0_t1_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t0_t1_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t0_t1_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t0_t1_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t0_t1_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t0_t1_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t0_t1_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t0_t1_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t0_t1_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t0_t1_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t0_t1_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t0_t1_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t0_t1_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t0_t1_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t0_t1_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t0_t1_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t0_t1_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t0_t1_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t0_t1_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t0_t1_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t0_t1_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t0_t1_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t0_t1_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t0_t1_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t0_t1_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t0_t1_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t0_t1_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t0_t1_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t0_t1_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t0_t1_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t0_t1_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t0_t1_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t0_t1_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t0_t1_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t0_t1_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t0_t1_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t0_t1_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t0_t1_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t0_t1_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t0_t1_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t0_t1_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t0_t1_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t0_t1_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t0_t1_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t0_t1_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t0_t1_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t0_t1_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t0_t1_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t0_t1_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t0_t1_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t0_t1_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t0_t1_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t0_t1_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t0_t1_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t0_t1_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t0_t1_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t0_t1_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t0_t1_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t0_t1_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t0_t1_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t0_t1_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t0_t1_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t0_t1_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t0_t1_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t0_t1_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t0_t1_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t0_t1_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t0_t1_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t0_t1_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t0_t1_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t0_t1_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t0_t1_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t0_t1_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t0_t1_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t0_t1_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t0_t1_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t0_t1_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t0_t1_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t0_t1_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t0_t1_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t0_t1_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t0_t1_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t0_t1_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t0_t1_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t0_t1_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t0_t1_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t0_t1_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t0_t1_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t0_t1_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t0_t1_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t0_t1_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t0_t1_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t0_t1_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t0_t1_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t0_t1_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t0_t1_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t0_t1_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t0_t1_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t0_t1_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t0_t1_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t0_t1_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t0_t1_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t0_t1_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t0_t1_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t0_t1_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t0_t1_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t0_t1_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t0_t1_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t0_t1_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t0_t1_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t0_t1_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t0_t1_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t0_t1_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t0_t1_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t0_t1_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t0_t1_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t0_t1_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t0_t1_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t0_t1_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t0_t1_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t0_t1_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t0_t1_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t0_t1_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t0_t1_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t0_t1_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t0_t1_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t0_t1_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t0_t1_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t0_t1_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t0_t1_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t0_t1_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t0_t1_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t0_t1_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t0_t1_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t0_t1_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t0_t1_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t0_t1_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t0_t1_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t0_t1_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t0_t1_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t0_t1_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t0_t1_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t0_t1_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t0_t1_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t0_t1_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t0_t1_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t0_t1_out = { AES_r1_t0_t1_k0, AES_r1_t0_t1_k0, ( AES_r1_t0_t1_k0 ^ AES_r1_t0_t1_k1 ), AES_r1_t0_t1_k1 };
    assign AES_r1_t0_t2_clk = AES_r1_t0_clk;
    assign AES_r1_t0_t2_in = AES_r1_t0_b2;
    assign AES_r1_t0_k2 = AES_r1_t0_t2_out;
    assign AES_r1_t0_t2_s0_clk = AES_r1_t0_t2_clk;
    assign AES_r1_t0_t2_s0_in = AES_r1_t0_t2_in;
    assign AES_r1_t0_t2_k0 = AES_r1_t0_t2_s0_out;
    always @ (  posedge AES_r1_t0_t2_s0_clk)
    begin
        case ( AES_r1_t0_t2_s0_in ) 
        8'h00:
        begin
            AES_r1_t0_t2_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t0_t2_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t0_t2_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t0_t2_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t0_t2_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t0_t2_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t0_t2_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t0_t2_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t0_t2_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t0_t2_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t0_t2_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t0_t2_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t0_t2_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t0_t2_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t0_t2_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t0_t2_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t0_t2_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t0_t2_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t0_t2_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t0_t2_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t0_t2_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t0_t2_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t0_t2_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t0_t2_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t0_t2_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t0_t2_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t0_t2_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t0_t2_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t0_t2_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t0_t2_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t0_t2_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t0_t2_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t0_t2_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t0_t2_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t0_t2_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t0_t2_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t0_t2_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t0_t2_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t0_t2_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t0_t2_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t0_t2_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t0_t2_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t2_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t0_t2_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t0_t2_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t0_t2_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t0_t2_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t0_t2_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t0_t2_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t0_t2_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t0_t2_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t0_t2_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t0_t2_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t0_t2_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t0_t2_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t0_t2_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t0_t2_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t0_t2_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t0_t2_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t0_t2_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t0_t2_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t0_t2_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t0_t2_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t0_t2_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t0_t2_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t0_t2_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t0_t2_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t0_t2_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t0_t2_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t0_t2_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t0_t2_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t0_t2_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t0_t2_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t0_t2_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t0_t2_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t0_t2_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t0_t2_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t0_t2_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t0_t2_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t0_t2_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t0_t2_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t0_t2_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t0_t2_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t0_t2_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t0_t2_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t0_t2_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t0_t2_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t0_t2_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t0_t2_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t0_t2_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t0_t2_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t0_t2_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t0_t2_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t0_t2_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t0_t2_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t0_t2_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t0_t2_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t0_t2_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t0_t2_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t0_t2_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t0_t2_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t0_t2_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t0_t2_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t0_t2_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t0_t2_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t0_t2_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t0_t2_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t0_t2_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t0_t2_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t0_t2_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t0_t2_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t0_t2_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t0_t2_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t0_t2_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t0_t2_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t0_t2_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t0_t2_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t0_t2_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t0_t2_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t0_t2_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t0_t2_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t0_t2_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t0_t2_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t0_t2_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t0_t2_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t0_t2_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t0_t2_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t0_t2_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t0_t2_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t0_t2_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t0_t2_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t0_t2_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t0_t2_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t0_t2_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t0_t2_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t0_t2_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t0_t2_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t0_t2_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t0_t2_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t0_t2_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t0_t2_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t0_t2_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t0_t2_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t0_t2_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t0_t2_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t0_t2_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t0_t2_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t0_t2_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t0_t2_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t0_t2_s4_clk = AES_r1_t0_t2_clk;
    assign AES_r1_t0_t2_s4_in = AES_r1_t0_t2_in;
    assign AES_r1_t0_t2_k1 = AES_r1_t0_t2_s4_out;
    always @ (  posedge AES_r1_t0_t2_s4_clk)
    begin
        case ( AES_r1_t0_t2_s4_in ) 
        8'h00:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t0_t2_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t0_t2_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t0_t2_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t0_t2_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t0_t2_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t0_t2_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t0_t2_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t0_t2_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t0_t2_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t0_t2_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t0_t2_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t0_t2_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t0_t2_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t0_t2_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t0_t2_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t0_t2_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t0_t2_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t0_t2_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t0_t2_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t0_t2_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t0_t2_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t0_t2_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t0_t2_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t0_t2_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t0_t2_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t0_t2_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t0_t2_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t0_t2_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t0_t2_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t0_t2_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t0_t2_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t0_t2_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t0_t2_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t0_t2_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t0_t2_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t0_t2_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t0_t2_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t0_t2_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t0_t2_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t0_t2_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t0_t2_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t0_t2_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t0_t2_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t0_t2_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t0_t2_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t0_t2_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t0_t2_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t0_t2_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t0_t2_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t0_t2_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t0_t2_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t0_t2_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t0_t2_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t0_t2_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t0_t2_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t0_t2_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t0_t2_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t0_t2_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t0_t2_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t0_t2_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t0_t2_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t0_t2_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t0_t2_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t0_t2_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t0_t2_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t0_t2_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t0_t2_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t0_t2_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t0_t2_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t0_t2_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t0_t2_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t0_t2_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t0_t2_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t0_t2_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t0_t2_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t0_t2_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t0_t2_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t0_t2_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t0_t2_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t0_t2_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t0_t2_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t0_t2_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t0_t2_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t0_t2_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t0_t2_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t0_t2_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t0_t2_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t0_t2_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t0_t2_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t0_t2_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t0_t2_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t0_t2_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t0_t2_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t0_t2_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t0_t2_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t0_t2_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t0_t2_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t0_t2_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t0_t2_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t0_t2_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t0_t2_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t0_t2_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t0_t2_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t0_t2_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t0_t2_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t0_t2_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t0_t2_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t0_t2_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t0_t2_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t0_t2_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t0_t2_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t0_t2_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t0_t2_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t0_t2_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t0_t2_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t0_t2_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t0_t2_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t0_t2_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t0_t2_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t0_t2_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t0_t2_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t0_t2_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t0_t2_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t0_t2_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t0_t2_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t0_t2_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t0_t2_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t0_t2_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t0_t2_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t0_t2_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t0_t2_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t0_t2_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t0_t2_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t0_t2_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t0_t2_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t0_t2_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t0_t2_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t0_t2_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t0_t2_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t0_t2_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t0_t2_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t0_t2_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t0_t2_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t0_t2_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t0_t2_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t0_t2_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t0_t2_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t0_t2_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t0_t2_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t0_t2_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t0_t2_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t0_t2_out = { AES_r1_t0_t2_k0, AES_r1_t0_t2_k0, ( AES_r1_t0_t2_k0 ^ AES_r1_t0_t2_k1 ), AES_r1_t0_t2_k1 };
    assign AES_r1_t0_t3_clk = AES_r1_t0_clk;
    assign AES_r1_t0_t3_in = AES_r1_t0_b3;
    assign AES_r1_t0_p3 = AES_r1_t0_t3_out;
    assign AES_r1_t0_t3_s0_clk = AES_r1_t0_t3_clk;
    assign AES_r1_t0_t3_s0_in = AES_r1_t0_t3_in;
    assign AES_r1_t0_t3_k0 = AES_r1_t0_t3_s0_out;
    always @ (  posedge AES_r1_t0_t3_s0_clk)
    begin
        case ( AES_r1_t0_t3_s0_in ) 
        8'h00:
        begin
            AES_r1_t0_t3_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t0_t3_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t0_t3_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t0_t3_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t0_t3_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t0_t3_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t0_t3_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t0_t3_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t0_t3_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t0_t3_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t0_t3_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t0_t3_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t0_t3_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t0_t3_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t0_t3_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t0_t3_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t0_t3_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t0_t3_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t0_t3_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t0_t3_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t0_t3_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t0_t3_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t0_t3_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t0_t3_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t0_t3_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t0_t3_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t0_t3_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t0_t3_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t0_t3_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t0_t3_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t0_t3_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t0_t3_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t0_t3_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t0_t3_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t0_t3_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t0_t3_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t0_t3_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t0_t3_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t0_t3_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t0_t3_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t0_t3_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t0_t3_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t3_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t0_t3_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t0_t3_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t0_t3_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t0_t3_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t0_t3_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t0_t3_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t0_t3_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t0_t3_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t0_t3_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t0_t3_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t0_t3_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t0_t3_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t0_t3_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t0_t3_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t0_t3_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t0_t3_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t0_t3_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t0_t3_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t0_t3_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t0_t3_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t0_t3_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t0_t3_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t0_t3_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t0_t3_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t0_t3_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t0_t3_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t0_t3_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t0_t3_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t0_t3_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t0_t3_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t0_t3_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t0_t3_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t0_t3_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t0_t3_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t0_t3_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t0_t3_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t0_t3_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t0_t3_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t0_t3_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t0_t3_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t0_t3_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t0_t3_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t0_t3_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t0_t3_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t0_t3_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t0_t3_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t0_t3_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t0_t3_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t0_t3_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t0_t3_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t0_t3_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t0_t3_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t0_t3_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t0_t3_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t0_t3_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t0_t3_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t0_t3_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t0_t3_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t0_t3_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t0_t3_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t0_t3_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t0_t3_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t0_t3_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t0_t3_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t0_t3_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t0_t3_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t0_t3_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t0_t3_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t0_t3_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t0_t3_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t0_t3_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t0_t3_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t0_t3_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t0_t3_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t0_t3_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t0_t3_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t0_t3_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t0_t3_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t0_t3_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t0_t3_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t0_t3_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t0_t3_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t0_t3_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t0_t3_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t0_t3_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t0_t3_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t0_t3_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t0_t3_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t0_t3_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t0_t3_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t0_t3_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t0_t3_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t0_t3_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t0_t3_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t0_t3_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t0_t3_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t0_t3_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t0_t3_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t0_t3_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t0_t3_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t0_t3_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t0_t3_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t0_t3_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t0_t3_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t0_t3_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t0_t3_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t0_t3_s4_clk = AES_r1_t0_t3_clk;
    assign AES_r1_t0_t3_s4_in = AES_r1_t0_t3_in;
    assign AES_r1_t0_t3_k1 = AES_r1_t0_t3_s4_out;
    always @ (  posedge AES_r1_t0_t3_s4_clk)
    begin
        case ( AES_r1_t0_t3_s4_in ) 
        8'h00:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t0_t3_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t0_t3_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t0_t3_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t0_t3_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t0_t3_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t0_t3_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t0_t3_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t0_t3_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t0_t3_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t0_t3_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t0_t3_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t0_t3_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t0_t3_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t0_t3_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t0_t3_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t0_t3_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t0_t3_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t0_t3_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t0_t3_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t0_t3_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t0_t3_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t0_t3_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t0_t3_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t0_t3_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t0_t3_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t0_t3_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t0_t3_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t0_t3_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t0_t3_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t0_t3_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t0_t3_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t0_t3_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t0_t3_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t0_t3_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t0_t3_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t0_t3_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t0_t3_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t0_t3_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t0_t3_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t0_t3_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t0_t3_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t0_t3_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t0_t3_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t0_t3_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t0_t3_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t0_t3_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t0_t3_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t0_t3_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t0_t3_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t0_t3_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t0_t3_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t0_t3_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t0_t3_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t0_t3_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t0_t3_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t0_t3_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t0_t3_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t0_t3_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t0_t3_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t0_t3_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t0_t3_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t0_t3_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t0_t3_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t0_t3_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t0_t3_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t0_t3_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t0_t3_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t0_t3_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t0_t3_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t0_t3_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t0_t3_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t0_t3_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t0_t3_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t0_t3_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t0_t3_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t0_t3_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t0_t3_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t0_t3_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t0_t3_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t0_t3_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t0_t3_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t0_t3_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t0_t3_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t0_t3_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t0_t3_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t0_t3_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t0_t3_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t0_t3_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t0_t3_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t0_t3_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t0_t3_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t0_t3_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t0_t3_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t0_t3_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t0_t3_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t0_t3_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t0_t3_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t0_t3_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t0_t3_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t0_t3_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t0_t3_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t0_t3_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t0_t3_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t0_t3_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t0_t3_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t0_t3_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t0_t3_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t0_t3_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t0_t3_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t0_t3_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t0_t3_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t0_t3_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t0_t3_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t0_t3_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t0_t3_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t0_t3_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t0_t3_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t0_t3_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t0_t3_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t0_t3_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t0_t3_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t0_t3_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t0_t3_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t0_t3_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t0_t3_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t0_t3_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t0_t3_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t0_t3_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t0_t3_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t0_t3_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t0_t3_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t0_t3_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t0_t3_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t0_t3_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t0_t3_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t0_t3_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t0_t3_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t0_t3_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t0_t3_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t0_t3_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t0_t3_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t0_t3_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t0_t3_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t0_t3_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t0_t3_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t0_t3_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t0_t3_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t0_t3_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t0_t3_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t0_t3_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t0_t3_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t0_t3_out = { AES_r1_t0_t3_k0, AES_r1_t0_t3_k0, ( AES_r1_t0_t3_k0 ^ AES_r1_t0_t3_k1 ), AES_r1_t0_t3_k1 };
    assign AES_r1_t1_clk = AES_r1_clk;
    assign AES_r1_t1_state = AES_r1_s1;
    assign AES_r1_p10 = AES_r1_t1_p0;
    assign AES_r1_p11 = AES_r1_t1_p1;
    assign AES_r1_p12 = AES_r1_t1_p2;
    assign AES_r1_p13 = AES_r1_t1_p3;
    assign AES_r1_t1_p0 = { AES_r1_t1_k0[7:0], AES_r1_t1_k0[31:8] };
    assign AES_r1_t1_p1 = { AES_r1_t1_k1[15:0], AES_r1_t1_k1[31:16] };
    assign AES_r1_t1_p2 = { AES_r1_t1_k2[23:0], AES_r1_t1_k2[31:24] };
    assign AES_r1_t1_b0 = AES_r1_t1_state[31:24];
    assign AES_r1_t1_b1 = AES_r1_t1_state[23:16];
    assign AES_r1_t1_b2 = AES_r1_t1_state[15:8];
    assign AES_r1_t1_b3 = AES_r1_t1_state[7:0];
    assign AES_r1_t1_t0_clk = AES_r1_t1_clk;
    assign AES_r1_t1_t0_in = AES_r1_t1_b0;
    assign AES_r1_t1_k0 = AES_r1_t1_t0_out;
    assign AES_r1_t1_t0_s0_clk = AES_r1_t1_t0_clk;
    assign AES_r1_t1_t0_s0_in = AES_r1_t1_t0_in;
    assign AES_r1_t1_t0_k0 = AES_r1_t1_t0_s0_out;
    always @ (  posedge AES_r1_t1_t0_s0_clk)
    begin
        case ( AES_r1_t1_t0_s0_in ) 
        8'h00:
        begin
            AES_r1_t1_t0_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t1_t0_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t1_t0_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t1_t0_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t1_t0_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t1_t0_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t1_t0_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t1_t0_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t1_t0_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t1_t0_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t1_t0_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t1_t0_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t1_t0_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t1_t0_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t1_t0_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t1_t0_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t1_t0_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t1_t0_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t1_t0_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t1_t0_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t1_t0_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t1_t0_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t1_t0_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t1_t0_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t1_t0_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t1_t0_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t1_t0_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t1_t0_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t1_t0_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t1_t0_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t1_t0_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t1_t0_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t1_t0_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t1_t0_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t1_t0_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t1_t0_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t1_t0_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t1_t0_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t1_t0_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t1_t0_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t1_t0_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t1_t0_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t0_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t1_t0_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t1_t0_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t1_t0_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t1_t0_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t1_t0_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t1_t0_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t1_t0_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t1_t0_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t1_t0_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t1_t0_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t1_t0_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t1_t0_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t1_t0_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t1_t0_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t1_t0_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t1_t0_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t1_t0_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t1_t0_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t1_t0_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t1_t0_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t1_t0_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t1_t0_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t1_t0_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t1_t0_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t1_t0_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t1_t0_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t1_t0_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t1_t0_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t1_t0_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t1_t0_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t1_t0_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t1_t0_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t1_t0_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t1_t0_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t1_t0_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t1_t0_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t1_t0_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t1_t0_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t1_t0_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t1_t0_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t1_t0_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t1_t0_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t1_t0_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t1_t0_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t1_t0_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t1_t0_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t1_t0_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t1_t0_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t1_t0_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t1_t0_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t1_t0_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t1_t0_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t1_t0_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t1_t0_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t1_t0_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t1_t0_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t1_t0_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t1_t0_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t1_t0_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t1_t0_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t1_t0_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t1_t0_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t1_t0_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t1_t0_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t1_t0_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t1_t0_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t1_t0_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t1_t0_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t1_t0_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t1_t0_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t1_t0_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t1_t0_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t1_t0_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t1_t0_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t1_t0_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t1_t0_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t1_t0_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t1_t0_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t1_t0_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t1_t0_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t1_t0_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t1_t0_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t1_t0_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t1_t0_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t1_t0_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t1_t0_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t1_t0_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t1_t0_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t1_t0_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t1_t0_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t1_t0_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t1_t0_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t1_t0_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t1_t0_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t1_t0_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t1_t0_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t1_t0_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t1_t0_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t1_t0_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t1_t0_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t1_t0_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t1_t0_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t1_t0_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t1_t0_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t1_t0_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t1_t0_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t1_t0_s4_clk = AES_r1_t1_t0_clk;
    assign AES_r1_t1_t0_s4_in = AES_r1_t1_t0_in;
    assign AES_r1_t1_t0_k1 = AES_r1_t1_t0_s4_out;
    always @ (  posedge AES_r1_t1_t0_s4_clk)
    begin
        case ( AES_r1_t1_t0_s4_in ) 
        8'h00:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t1_t0_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t1_t0_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t1_t0_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t1_t0_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t1_t0_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t1_t0_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t1_t0_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t1_t0_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t1_t0_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t1_t0_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t1_t0_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t1_t0_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t1_t0_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t1_t0_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t1_t0_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t1_t0_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t1_t0_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t1_t0_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t1_t0_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t1_t0_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t1_t0_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t1_t0_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t1_t0_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t1_t0_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t1_t0_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t1_t0_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t1_t0_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t1_t0_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t1_t0_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t1_t0_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t1_t0_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t1_t0_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t1_t0_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t1_t0_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t1_t0_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t1_t0_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t1_t0_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t1_t0_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t1_t0_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t1_t0_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t1_t0_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t1_t0_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t1_t0_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t1_t0_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t1_t0_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t1_t0_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t1_t0_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t1_t0_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t1_t0_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t1_t0_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t1_t0_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t1_t0_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t1_t0_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t1_t0_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t1_t0_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t1_t0_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t1_t0_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t1_t0_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t1_t0_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t1_t0_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t1_t0_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t1_t0_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t1_t0_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t1_t0_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t1_t0_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t1_t0_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t1_t0_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t1_t0_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t1_t0_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t1_t0_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t1_t0_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t1_t0_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t1_t0_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t1_t0_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t1_t0_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t1_t0_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t1_t0_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t1_t0_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t1_t0_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t1_t0_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t1_t0_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t1_t0_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t1_t0_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t1_t0_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t1_t0_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t1_t0_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t1_t0_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t1_t0_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t1_t0_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t1_t0_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t1_t0_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t1_t0_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t1_t0_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t1_t0_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t1_t0_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t1_t0_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t1_t0_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t1_t0_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t1_t0_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t1_t0_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t1_t0_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t1_t0_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t1_t0_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t1_t0_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t1_t0_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t1_t0_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t1_t0_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t1_t0_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t1_t0_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t1_t0_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t1_t0_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t1_t0_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t1_t0_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t1_t0_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t1_t0_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t1_t0_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t1_t0_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t1_t0_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t1_t0_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t1_t0_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t1_t0_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t1_t0_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t1_t0_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t1_t0_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t1_t0_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t1_t0_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t1_t0_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t1_t0_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t1_t0_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t1_t0_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t1_t0_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t1_t0_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t1_t0_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t1_t0_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t1_t0_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t1_t0_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t1_t0_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t1_t0_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t1_t0_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t1_t0_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t1_t0_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t1_t0_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t1_t0_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t1_t0_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t1_t0_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t1_t0_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t1_t0_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t1_t0_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t1_t0_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t1_t0_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t1_t0_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t1_t0_out = { AES_r1_t1_t0_k0, AES_r1_t1_t0_k0, ( AES_r1_t1_t0_k0 ^ AES_r1_t1_t0_k1 ), AES_r1_t1_t0_k1 };
    assign AES_r1_t1_t1_clk = AES_r1_t1_clk;
    assign AES_r1_t1_t1_in = AES_r1_t1_b1;
    assign AES_r1_t1_k1 = AES_r1_t1_t1_out;
    assign AES_r1_t1_t1_s0_clk = AES_r1_t1_t1_clk;
    assign AES_r1_t1_t1_s0_in = AES_r1_t1_t1_in;
    assign AES_r1_t1_t1_k0 = AES_r1_t1_t1_s0_out;
    always @ (  posedge AES_r1_t1_t1_s0_clk)
    begin
        case ( AES_r1_t1_t1_s0_in ) 
        8'h00:
        begin
            AES_r1_t1_t1_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t1_t1_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t1_t1_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t1_t1_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t1_t1_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t1_t1_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t1_t1_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t1_t1_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t1_t1_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t1_t1_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t1_t1_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t1_t1_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t1_t1_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t1_t1_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t1_t1_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t1_t1_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t1_t1_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t1_t1_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t1_t1_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t1_t1_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t1_t1_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t1_t1_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t1_t1_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t1_t1_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t1_t1_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t1_t1_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t1_t1_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t1_t1_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t1_t1_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t1_t1_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t1_t1_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t1_t1_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t1_t1_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t1_t1_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t1_t1_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t1_t1_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t1_t1_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t1_t1_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t1_t1_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t1_t1_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t1_t1_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t1_t1_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t1_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t1_t1_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t1_t1_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t1_t1_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t1_t1_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t1_t1_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t1_t1_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t1_t1_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t1_t1_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t1_t1_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t1_t1_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t1_t1_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t1_t1_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t1_t1_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t1_t1_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t1_t1_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t1_t1_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t1_t1_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t1_t1_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t1_t1_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t1_t1_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t1_t1_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t1_t1_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t1_t1_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t1_t1_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t1_t1_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t1_t1_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t1_t1_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t1_t1_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t1_t1_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t1_t1_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t1_t1_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t1_t1_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t1_t1_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t1_t1_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t1_t1_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t1_t1_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t1_t1_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t1_t1_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t1_t1_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t1_t1_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t1_t1_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t1_t1_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t1_t1_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t1_t1_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t1_t1_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t1_t1_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t1_t1_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t1_t1_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t1_t1_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t1_t1_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t1_t1_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t1_t1_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t1_t1_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t1_t1_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t1_t1_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t1_t1_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t1_t1_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t1_t1_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t1_t1_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t1_t1_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t1_t1_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t1_t1_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t1_t1_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t1_t1_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t1_t1_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t1_t1_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t1_t1_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t1_t1_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t1_t1_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t1_t1_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t1_t1_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t1_t1_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t1_t1_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t1_t1_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t1_t1_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t1_t1_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t1_t1_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t1_t1_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t1_t1_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t1_t1_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t1_t1_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t1_t1_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t1_t1_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t1_t1_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t1_t1_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t1_t1_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t1_t1_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t1_t1_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t1_t1_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t1_t1_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t1_t1_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t1_t1_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t1_t1_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t1_t1_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t1_t1_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t1_t1_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t1_t1_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t1_t1_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t1_t1_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t1_t1_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t1_t1_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t1_t1_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t1_t1_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t1_t1_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t1_t1_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t1_t1_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t1_t1_s4_clk = AES_r1_t1_t1_clk;
    assign AES_r1_t1_t1_s4_in = AES_r1_t1_t1_in;
    assign AES_r1_t1_t1_k1 = AES_r1_t1_t1_s4_out;
    always @ (  posedge AES_r1_t1_t1_s4_clk)
    begin
        case ( AES_r1_t1_t1_s4_in ) 
        8'h00:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t1_t1_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t1_t1_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t1_t1_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t1_t1_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t1_t1_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t1_t1_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t1_t1_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t1_t1_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t1_t1_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t1_t1_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t1_t1_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t1_t1_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t1_t1_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t1_t1_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t1_t1_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t1_t1_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t1_t1_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t1_t1_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t1_t1_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t1_t1_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t1_t1_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t1_t1_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t1_t1_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t1_t1_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t1_t1_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t1_t1_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t1_t1_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t1_t1_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t1_t1_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t1_t1_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t1_t1_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t1_t1_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t1_t1_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t1_t1_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t1_t1_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t1_t1_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t1_t1_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t1_t1_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t1_t1_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t1_t1_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t1_t1_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t1_t1_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t1_t1_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t1_t1_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t1_t1_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t1_t1_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t1_t1_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t1_t1_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t1_t1_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t1_t1_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t1_t1_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t1_t1_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t1_t1_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t1_t1_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t1_t1_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t1_t1_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t1_t1_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t1_t1_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t1_t1_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t1_t1_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t1_t1_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t1_t1_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t1_t1_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t1_t1_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t1_t1_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t1_t1_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t1_t1_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t1_t1_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t1_t1_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t1_t1_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t1_t1_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t1_t1_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t1_t1_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t1_t1_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t1_t1_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t1_t1_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t1_t1_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t1_t1_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t1_t1_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t1_t1_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t1_t1_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t1_t1_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t1_t1_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t1_t1_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t1_t1_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t1_t1_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t1_t1_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t1_t1_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t1_t1_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t1_t1_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t1_t1_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t1_t1_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t1_t1_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t1_t1_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t1_t1_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t1_t1_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t1_t1_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t1_t1_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t1_t1_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t1_t1_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t1_t1_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t1_t1_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t1_t1_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t1_t1_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t1_t1_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t1_t1_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t1_t1_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t1_t1_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t1_t1_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t1_t1_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t1_t1_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t1_t1_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t1_t1_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t1_t1_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t1_t1_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t1_t1_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t1_t1_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t1_t1_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t1_t1_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t1_t1_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t1_t1_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t1_t1_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t1_t1_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t1_t1_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t1_t1_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t1_t1_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t1_t1_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t1_t1_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t1_t1_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t1_t1_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t1_t1_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t1_t1_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t1_t1_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t1_t1_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t1_t1_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t1_t1_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t1_t1_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t1_t1_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t1_t1_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t1_t1_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t1_t1_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t1_t1_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t1_t1_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t1_t1_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t1_t1_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t1_t1_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t1_t1_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t1_t1_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t1_t1_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t1_t1_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t1_t1_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t1_t1_out = { AES_r1_t1_t1_k0, AES_r1_t1_t1_k0, ( AES_r1_t1_t1_k0 ^ AES_r1_t1_t1_k1 ), AES_r1_t1_t1_k1 };
    assign AES_r1_t1_t2_clk = AES_r1_t1_clk;
    assign AES_r1_t1_t2_in = AES_r1_t1_b2;
    assign AES_r1_t1_k2 = AES_r1_t1_t2_out;
    assign AES_r1_t1_t2_s0_clk = AES_r1_t1_t2_clk;
    assign AES_r1_t1_t2_s0_in = AES_r1_t1_t2_in;
    assign AES_r1_t1_t2_k0 = AES_r1_t1_t2_s0_out;
    always @ (  posedge AES_r1_t1_t2_s0_clk)
    begin
        case ( AES_r1_t1_t2_s0_in ) 
        8'h00:
        begin
            AES_r1_t1_t2_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t1_t2_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t1_t2_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t1_t2_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t1_t2_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t1_t2_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t1_t2_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t1_t2_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t1_t2_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t1_t2_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t1_t2_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t1_t2_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t1_t2_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t1_t2_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t1_t2_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t1_t2_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t1_t2_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t1_t2_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t1_t2_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t1_t2_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t1_t2_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t1_t2_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t1_t2_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t1_t2_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t1_t2_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t1_t2_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t1_t2_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t1_t2_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t1_t2_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t1_t2_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t1_t2_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t1_t2_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t1_t2_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t1_t2_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t1_t2_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t1_t2_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t1_t2_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t1_t2_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t1_t2_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t1_t2_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t1_t2_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t1_t2_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t2_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t1_t2_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t1_t2_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t1_t2_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t1_t2_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t1_t2_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t1_t2_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t1_t2_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t1_t2_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t1_t2_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t1_t2_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t1_t2_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t1_t2_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t1_t2_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t1_t2_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t1_t2_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t1_t2_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t1_t2_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t1_t2_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t1_t2_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t1_t2_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t1_t2_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t1_t2_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t1_t2_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t1_t2_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t1_t2_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t1_t2_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t1_t2_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t1_t2_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t1_t2_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t1_t2_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t1_t2_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t1_t2_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t1_t2_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t1_t2_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t1_t2_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t1_t2_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t1_t2_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t1_t2_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t1_t2_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t1_t2_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t1_t2_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t1_t2_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t1_t2_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t1_t2_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t1_t2_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t1_t2_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t1_t2_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t1_t2_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t1_t2_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t1_t2_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t1_t2_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t1_t2_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t1_t2_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t1_t2_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t1_t2_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t1_t2_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t1_t2_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t1_t2_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t1_t2_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t1_t2_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t1_t2_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t1_t2_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t1_t2_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t1_t2_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t1_t2_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t1_t2_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t1_t2_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t1_t2_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t1_t2_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t1_t2_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t1_t2_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t1_t2_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t1_t2_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t1_t2_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t1_t2_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t1_t2_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t1_t2_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t1_t2_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t1_t2_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t1_t2_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t1_t2_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t1_t2_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t1_t2_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t1_t2_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t1_t2_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t1_t2_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t1_t2_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t1_t2_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t1_t2_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t1_t2_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t1_t2_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t1_t2_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t1_t2_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t1_t2_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t1_t2_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t1_t2_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t1_t2_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t1_t2_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t1_t2_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t1_t2_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t1_t2_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t1_t2_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t1_t2_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t1_t2_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t1_t2_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t1_t2_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t1_t2_s4_clk = AES_r1_t1_t2_clk;
    assign AES_r1_t1_t2_s4_in = AES_r1_t1_t2_in;
    assign AES_r1_t1_t2_k1 = AES_r1_t1_t2_s4_out;
    always @ (  posedge AES_r1_t1_t2_s4_clk)
    begin
        case ( AES_r1_t1_t2_s4_in ) 
        8'h00:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t1_t2_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t1_t2_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t1_t2_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t1_t2_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t1_t2_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t1_t2_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t1_t2_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t1_t2_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t1_t2_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t1_t2_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t1_t2_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t1_t2_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t1_t2_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t1_t2_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t1_t2_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t1_t2_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t1_t2_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t1_t2_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t1_t2_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t1_t2_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t1_t2_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t1_t2_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t1_t2_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t1_t2_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t1_t2_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t1_t2_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t1_t2_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t1_t2_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t1_t2_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t1_t2_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t1_t2_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t1_t2_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t1_t2_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t1_t2_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t1_t2_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t1_t2_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t1_t2_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t1_t2_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t1_t2_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t1_t2_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t1_t2_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t1_t2_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t1_t2_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t1_t2_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t1_t2_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t1_t2_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t1_t2_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t1_t2_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t1_t2_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t1_t2_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t1_t2_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t1_t2_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t1_t2_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t1_t2_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t1_t2_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t1_t2_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t1_t2_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t1_t2_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t1_t2_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t1_t2_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t1_t2_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t1_t2_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t1_t2_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t1_t2_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t1_t2_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t1_t2_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t1_t2_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t1_t2_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t1_t2_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t1_t2_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t1_t2_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t1_t2_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t1_t2_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t1_t2_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t1_t2_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t1_t2_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t1_t2_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t1_t2_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t1_t2_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t1_t2_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t1_t2_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t1_t2_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t1_t2_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t1_t2_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t1_t2_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t1_t2_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t1_t2_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t1_t2_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t1_t2_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t1_t2_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t1_t2_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t1_t2_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t1_t2_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t1_t2_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t1_t2_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t1_t2_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t1_t2_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t1_t2_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t1_t2_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t1_t2_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t1_t2_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t1_t2_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t1_t2_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t1_t2_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t1_t2_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t1_t2_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t1_t2_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t1_t2_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t1_t2_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t1_t2_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t1_t2_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t1_t2_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t1_t2_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t1_t2_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t1_t2_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t1_t2_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t1_t2_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t1_t2_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t1_t2_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t1_t2_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t1_t2_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t1_t2_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t1_t2_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t1_t2_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t1_t2_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t1_t2_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t1_t2_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t1_t2_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t1_t2_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t1_t2_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t1_t2_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t1_t2_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t1_t2_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t1_t2_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t1_t2_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t1_t2_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t1_t2_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t1_t2_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t1_t2_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t1_t2_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t1_t2_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t1_t2_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t1_t2_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t1_t2_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t1_t2_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t1_t2_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t1_t2_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t1_t2_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t1_t2_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t1_t2_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t1_t2_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t1_t2_out = { AES_r1_t1_t2_k0, AES_r1_t1_t2_k0, ( AES_r1_t1_t2_k0 ^ AES_r1_t1_t2_k1 ), AES_r1_t1_t2_k1 };
    assign AES_r1_t1_t3_clk = AES_r1_t1_clk;
    assign AES_r1_t1_t3_in = AES_r1_t1_b3;
    assign AES_r1_t1_p3 = AES_r1_t1_t3_out;
    assign AES_r1_t1_t3_s0_clk = AES_r1_t1_t3_clk;
    assign AES_r1_t1_t3_s0_in = AES_r1_t1_t3_in;
    assign AES_r1_t1_t3_k0 = AES_r1_t1_t3_s0_out;
    always @ (  posedge AES_r1_t1_t3_s0_clk)
    begin
        case ( AES_r1_t1_t3_s0_in ) 
        8'h00:
        begin
            AES_r1_t1_t3_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t1_t3_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t1_t3_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t1_t3_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t1_t3_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t1_t3_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t1_t3_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t1_t3_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t1_t3_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t1_t3_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t1_t3_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t1_t3_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t1_t3_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t1_t3_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t1_t3_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t1_t3_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t1_t3_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t1_t3_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t1_t3_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t1_t3_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t1_t3_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t1_t3_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t1_t3_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t1_t3_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t1_t3_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t1_t3_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t1_t3_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t1_t3_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t1_t3_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t1_t3_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t1_t3_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t1_t3_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t1_t3_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t1_t3_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t1_t3_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t1_t3_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t1_t3_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t1_t3_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t1_t3_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t1_t3_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t1_t3_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t1_t3_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t3_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t1_t3_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t1_t3_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t1_t3_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t1_t3_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t1_t3_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t1_t3_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t1_t3_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t1_t3_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t1_t3_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t1_t3_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t1_t3_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t1_t3_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t1_t3_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t1_t3_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t1_t3_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t1_t3_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t1_t3_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t1_t3_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t1_t3_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t1_t3_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t1_t3_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t1_t3_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t1_t3_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t1_t3_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t1_t3_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t1_t3_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t1_t3_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t1_t3_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t1_t3_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t1_t3_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t1_t3_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t1_t3_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t1_t3_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t1_t3_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t1_t3_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t1_t3_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t1_t3_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t1_t3_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t1_t3_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t1_t3_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t1_t3_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t1_t3_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t1_t3_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t1_t3_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t1_t3_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t1_t3_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t1_t3_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t1_t3_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t1_t3_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t1_t3_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t1_t3_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t1_t3_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t1_t3_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t1_t3_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t1_t3_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t1_t3_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t1_t3_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t1_t3_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t1_t3_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t1_t3_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t1_t3_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t1_t3_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t1_t3_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t1_t3_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t1_t3_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t1_t3_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t1_t3_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t1_t3_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t1_t3_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t1_t3_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t1_t3_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t1_t3_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t1_t3_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t1_t3_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t1_t3_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t1_t3_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t1_t3_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t1_t3_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t1_t3_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t1_t3_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t1_t3_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t1_t3_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t1_t3_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t1_t3_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t1_t3_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t1_t3_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t1_t3_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t1_t3_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t1_t3_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t1_t3_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t1_t3_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t1_t3_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t1_t3_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t1_t3_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t1_t3_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t1_t3_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t1_t3_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t1_t3_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t1_t3_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t1_t3_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t1_t3_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t1_t3_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t1_t3_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t1_t3_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t1_t3_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t1_t3_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t1_t3_s4_clk = AES_r1_t1_t3_clk;
    assign AES_r1_t1_t3_s4_in = AES_r1_t1_t3_in;
    assign AES_r1_t1_t3_k1 = AES_r1_t1_t3_s4_out;
    always @ (  posedge AES_r1_t1_t3_s4_clk)
    begin
        case ( AES_r1_t1_t3_s4_in ) 
        8'h00:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t1_t3_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t1_t3_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t1_t3_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t1_t3_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t1_t3_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t1_t3_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t1_t3_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t1_t3_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t1_t3_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t1_t3_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t1_t3_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t1_t3_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t1_t3_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t1_t3_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t1_t3_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t1_t3_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t1_t3_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t1_t3_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t1_t3_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t1_t3_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t1_t3_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t1_t3_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t1_t3_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t1_t3_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t1_t3_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t1_t3_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t1_t3_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t1_t3_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t1_t3_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t1_t3_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t1_t3_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t1_t3_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t1_t3_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t1_t3_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t1_t3_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t1_t3_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t1_t3_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t1_t3_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t1_t3_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t1_t3_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t1_t3_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t1_t3_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t1_t3_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t1_t3_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t1_t3_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t1_t3_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t1_t3_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t1_t3_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t1_t3_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t1_t3_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t1_t3_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t1_t3_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t1_t3_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t1_t3_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t1_t3_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t1_t3_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t1_t3_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t1_t3_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t1_t3_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t1_t3_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t1_t3_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t1_t3_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t1_t3_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t1_t3_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t1_t3_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t1_t3_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t1_t3_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t1_t3_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t1_t3_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t1_t3_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t1_t3_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t1_t3_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t1_t3_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t1_t3_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t1_t3_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t1_t3_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t1_t3_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t1_t3_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t1_t3_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t1_t3_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t1_t3_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t1_t3_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t1_t3_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t1_t3_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t1_t3_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t1_t3_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t1_t3_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t1_t3_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t1_t3_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t1_t3_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t1_t3_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t1_t3_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t1_t3_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t1_t3_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t1_t3_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t1_t3_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t1_t3_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t1_t3_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t1_t3_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t1_t3_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t1_t3_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t1_t3_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t1_t3_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t1_t3_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t1_t3_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t1_t3_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t1_t3_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t1_t3_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t1_t3_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t1_t3_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t1_t3_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t1_t3_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t1_t3_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t1_t3_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t1_t3_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t1_t3_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t1_t3_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t1_t3_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t1_t3_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t1_t3_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t1_t3_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t1_t3_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t1_t3_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t1_t3_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t1_t3_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t1_t3_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t1_t3_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t1_t3_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t1_t3_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t1_t3_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t1_t3_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t1_t3_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t1_t3_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t1_t3_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t1_t3_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t1_t3_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t1_t3_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t1_t3_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t1_t3_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t1_t3_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t1_t3_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t1_t3_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t1_t3_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t1_t3_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t1_t3_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t1_t3_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t1_t3_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t1_t3_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t1_t3_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t1_t3_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t1_t3_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t1_t3_out = { AES_r1_t1_t3_k0, AES_r1_t1_t3_k0, ( AES_r1_t1_t3_k0 ^ AES_r1_t1_t3_k1 ), AES_r1_t1_t3_k1 };
    assign AES_r1_t2_clk = AES_r1_clk;
    assign AES_r1_t2_state = AES_r1_s2;
    assign AES_r1_p20 = AES_r1_t2_p0;
    assign AES_r1_p21 = AES_r1_t2_p1;
    assign AES_r1_p22 = AES_r1_t2_p2;
    assign AES_r1_p23 = AES_r1_t2_p3;
    assign AES_r1_t2_p0 = { AES_r1_t2_k0[7:0], AES_r1_t2_k0[31:8] };
    assign AES_r1_t2_p1 = { AES_r1_t2_k1[15:0], AES_r1_t2_k1[31:16] };
    assign AES_r1_t2_p2 = { AES_r1_t2_k2[23:0], AES_r1_t2_k2[31:24] };
    assign AES_r1_t2_b0 = AES_r1_t2_state[31:24];
    assign AES_r1_t2_b1 = AES_r1_t2_state[23:16];
    assign AES_r1_t2_b2 = AES_r1_t2_state[15:8];
    assign AES_r1_t2_b3 = AES_r1_t2_state[7:0];
    assign AES_r1_t2_t0_clk = AES_r1_t2_clk;
    assign AES_r1_t2_t0_in = AES_r1_t2_b0;
    assign AES_r1_t2_k0 = AES_r1_t2_t0_out;
    assign AES_r1_t2_t0_s0_clk = AES_r1_t2_t0_clk;
    assign AES_r1_t2_t0_s0_in = AES_r1_t2_t0_in;
    assign AES_r1_t2_t0_k0 = AES_r1_t2_t0_s0_out;
    always @ (  posedge AES_r1_t2_t0_s0_clk)
    begin
        case ( AES_r1_t2_t0_s0_in ) 
        8'h00:
        begin
            AES_r1_t2_t0_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t2_t0_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t2_t0_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t2_t0_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t2_t0_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t2_t0_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t2_t0_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t2_t0_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t2_t0_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t2_t0_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t2_t0_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t2_t0_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t2_t0_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t2_t0_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t2_t0_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t2_t0_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t2_t0_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t2_t0_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t2_t0_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t2_t0_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t2_t0_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t2_t0_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t2_t0_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t2_t0_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t2_t0_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t2_t0_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t2_t0_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t2_t0_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t2_t0_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t2_t0_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t2_t0_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t2_t0_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t2_t0_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t2_t0_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t2_t0_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t2_t0_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t2_t0_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t2_t0_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t2_t0_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t2_t0_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t2_t0_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t2_t0_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t0_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t2_t0_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t2_t0_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t2_t0_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t2_t0_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t2_t0_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t2_t0_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t2_t0_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t2_t0_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t2_t0_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t2_t0_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t2_t0_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t2_t0_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t2_t0_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t2_t0_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t2_t0_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t2_t0_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t2_t0_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t2_t0_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t2_t0_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t2_t0_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t2_t0_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t2_t0_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t2_t0_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t2_t0_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t2_t0_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t2_t0_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t2_t0_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t2_t0_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t2_t0_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t2_t0_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t2_t0_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t2_t0_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t2_t0_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t2_t0_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t2_t0_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t2_t0_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t2_t0_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t2_t0_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t2_t0_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t2_t0_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t2_t0_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t2_t0_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t2_t0_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t2_t0_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t2_t0_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t2_t0_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t2_t0_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t2_t0_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t2_t0_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t2_t0_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t2_t0_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t2_t0_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t2_t0_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t2_t0_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t2_t0_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t2_t0_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t2_t0_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t2_t0_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t2_t0_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t2_t0_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t2_t0_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t2_t0_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t2_t0_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t2_t0_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t2_t0_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t2_t0_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t2_t0_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t2_t0_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t2_t0_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t2_t0_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t2_t0_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t2_t0_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t2_t0_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t2_t0_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t2_t0_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t2_t0_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t2_t0_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t2_t0_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t2_t0_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t2_t0_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t2_t0_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t2_t0_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t2_t0_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t2_t0_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t2_t0_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t2_t0_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t2_t0_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t2_t0_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t2_t0_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t2_t0_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t2_t0_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t2_t0_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t2_t0_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t2_t0_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t2_t0_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t2_t0_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t2_t0_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t2_t0_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t2_t0_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t2_t0_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t2_t0_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t2_t0_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t2_t0_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t2_t0_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t2_t0_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t2_t0_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t2_t0_s4_clk = AES_r1_t2_t0_clk;
    assign AES_r1_t2_t0_s4_in = AES_r1_t2_t0_in;
    assign AES_r1_t2_t0_k1 = AES_r1_t2_t0_s4_out;
    always @ (  posedge AES_r1_t2_t0_s4_clk)
    begin
        case ( AES_r1_t2_t0_s4_in ) 
        8'h00:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t2_t0_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t2_t0_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t2_t0_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t2_t0_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t2_t0_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t2_t0_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t2_t0_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t2_t0_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t2_t0_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t2_t0_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t2_t0_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t2_t0_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t2_t0_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t2_t0_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t2_t0_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t2_t0_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t2_t0_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t2_t0_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t2_t0_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t2_t0_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t2_t0_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t2_t0_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t2_t0_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t2_t0_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t2_t0_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t2_t0_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t2_t0_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t2_t0_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t2_t0_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t2_t0_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t2_t0_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t2_t0_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t2_t0_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t2_t0_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t2_t0_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t2_t0_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t2_t0_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t2_t0_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t2_t0_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t2_t0_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t2_t0_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t2_t0_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t2_t0_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t2_t0_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t2_t0_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t2_t0_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t2_t0_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t2_t0_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t2_t0_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t2_t0_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t2_t0_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t2_t0_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t2_t0_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t2_t0_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t2_t0_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t2_t0_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t2_t0_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t2_t0_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t2_t0_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t2_t0_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t2_t0_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t2_t0_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t2_t0_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t2_t0_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t2_t0_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t2_t0_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t2_t0_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t2_t0_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t2_t0_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t2_t0_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t2_t0_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t2_t0_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t2_t0_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t2_t0_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t2_t0_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t2_t0_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t2_t0_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t2_t0_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t2_t0_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t2_t0_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t2_t0_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t2_t0_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t2_t0_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t2_t0_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t2_t0_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t2_t0_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t2_t0_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t2_t0_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t2_t0_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t2_t0_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t2_t0_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t2_t0_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t2_t0_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t2_t0_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t2_t0_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t2_t0_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t2_t0_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t2_t0_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t2_t0_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t2_t0_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t2_t0_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t2_t0_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t2_t0_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t2_t0_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t2_t0_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t2_t0_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t2_t0_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t2_t0_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t2_t0_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t2_t0_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t2_t0_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t2_t0_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t2_t0_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t2_t0_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t2_t0_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t2_t0_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t2_t0_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t2_t0_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t2_t0_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t2_t0_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t2_t0_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t2_t0_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t2_t0_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t2_t0_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t2_t0_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t2_t0_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t2_t0_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t2_t0_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t2_t0_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t2_t0_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t2_t0_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t2_t0_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t2_t0_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t2_t0_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t2_t0_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t2_t0_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t2_t0_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t2_t0_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t2_t0_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t2_t0_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t2_t0_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t2_t0_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t2_t0_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t2_t0_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t2_t0_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t2_t0_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t2_t0_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t2_t0_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t2_t0_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t2_t0_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t2_t0_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t2_t0_out = { AES_r1_t2_t0_k0, AES_r1_t2_t0_k0, ( AES_r1_t2_t0_k0 ^ AES_r1_t2_t0_k1 ), AES_r1_t2_t0_k1 };
    assign AES_r1_t2_t1_clk = AES_r1_t2_clk;
    assign AES_r1_t2_t1_in = AES_r1_t2_b1;
    assign AES_r1_t2_k1 = AES_r1_t2_t1_out;
    assign AES_r1_t2_t1_s0_clk = AES_r1_t2_t1_clk;
    assign AES_r1_t2_t1_s0_in = AES_r1_t2_t1_in;
    assign AES_r1_t2_t1_k0 = AES_r1_t2_t1_s0_out;
    always @ (  posedge AES_r1_t2_t1_s0_clk)
    begin
        case ( AES_r1_t2_t1_s0_in ) 
        8'h00:
        begin
            AES_r1_t2_t1_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t2_t1_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t2_t1_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t2_t1_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t2_t1_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t2_t1_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t2_t1_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t2_t1_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t2_t1_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t2_t1_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t2_t1_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t2_t1_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t2_t1_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t2_t1_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t2_t1_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t2_t1_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t2_t1_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t2_t1_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t2_t1_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t2_t1_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t2_t1_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t2_t1_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t2_t1_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t2_t1_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t2_t1_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t2_t1_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t2_t1_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t2_t1_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t2_t1_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t2_t1_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t2_t1_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t2_t1_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t2_t1_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t2_t1_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t2_t1_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t2_t1_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t2_t1_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t2_t1_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t2_t1_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t2_t1_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t2_t1_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t2_t1_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t1_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t2_t1_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t2_t1_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t2_t1_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t2_t1_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t2_t1_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t2_t1_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t2_t1_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t2_t1_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t2_t1_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t2_t1_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t2_t1_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t2_t1_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t2_t1_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t2_t1_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t2_t1_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t2_t1_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t2_t1_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t2_t1_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t2_t1_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t2_t1_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t2_t1_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t2_t1_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t2_t1_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t2_t1_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t2_t1_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t2_t1_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t2_t1_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t2_t1_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t2_t1_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t2_t1_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t2_t1_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t2_t1_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t2_t1_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t2_t1_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t2_t1_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t2_t1_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t2_t1_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t2_t1_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t2_t1_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t2_t1_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t2_t1_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t2_t1_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t2_t1_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t2_t1_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t2_t1_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t2_t1_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t2_t1_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t2_t1_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t2_t1_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t2_t1_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t2_t1_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t2_t1_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t2_t1_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t2_t1_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t2_t1_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t2_t1_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t2_t1_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t2_t1_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t2_t1_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t2_t1_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t2_t1_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t2_t1_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t2_t1_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t2_t1_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t2_t1_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t2_t1_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t2_t1_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t2_t1_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t2_t1_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t2_t1_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t2_t1_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t2_t1_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t2_t1_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t2_t1_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t2_t1_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t2_t1_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t2_t1_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t2_t1_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t2_t1_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t2_t1_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t2_t1_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t2_t1_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t2_t1_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t2_t1_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t2_t1_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t2_t1_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t2_t1_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t2_t1_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t2_t1_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t2_t1_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t2_t1_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t2_t1_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t2_t1_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t2_t1_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t2_t1_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t2_t1_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t2_t1_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t2_t1_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t2_t1_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t2_t1_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t2_t1_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t2_t1_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t2_t1_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t2_t1_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t2_t1_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t2_t1_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t2_t1_s4_clk = AES_r1_t2_t1_clk;
    assign AES_r1_t2_t1_s4_in = AES_r1_t2_t1_in;
    assign AES_r1_t2_t1_k1 = AES_r1_t2_t1_s4_out;
    always @ (  posedge AES_r1_t2_t1_s4_clk)
    begin
        case ( AES_r1_t2_t1_s4_in ) 
        8'h00:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t2_t1_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t2_t1_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t2_t1_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t2_t1_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t2_t1_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t2_t1_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t2_t1_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t2_t1_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t2_t1_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t2_t1_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t2_t1_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t2_t1_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t2_t1_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t2_t1_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t2_t1_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t2_t1_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t2_t1_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t2_t1_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t2_t1_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t2_t1_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t2_t1_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t2_t1_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t2_t1_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t2_t1_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t2_t1_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t2_t1_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t2_t1_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t2_t1_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t2_t1_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t2_t1_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t2_t1_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t2_t1_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t2_t1_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t2_t1_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t2_t1_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t2_t1_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t2_t1_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t2_t1_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t2_t1_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t2_t1_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t2_t1_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t2_t1_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t2_t1_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t2_t1_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t2_t1_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t2_t1_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t2_t1_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t2_t1_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t2_t1_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t2_t1_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t2_t1_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t2_t1_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t2_t1_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t2_t1_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t2_t1_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t2_t1_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t2_t1_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t2_t1_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t2_t1_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t2_t1_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t2_t1_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t2_t1_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t2_t1_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t2_t1_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t2_t1_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t2_t1_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t2_t1_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t2_t1_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t2_t1_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t2_t1_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t2_t1_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t2_t1_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t2_t1_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t2_t1_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t2_t1_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t2_t1_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t2_t1_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t2_t1_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t2_t1_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t2_t1_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t2_t1_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t2_t1_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t2_t1_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t2_t1_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t2_t1_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t2_t1_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t2_t1_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t2_t1_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t2_t1_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t2_t1_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t2_t1_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t2_t1_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t2_t1_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t2_t1_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t2_t1_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t2_t1_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t2_t1_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t2_t1_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t2_t1_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t2_t1_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t2_t1_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t2_t1_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t2_t1_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t2_t1_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t2_t1_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t2_t1_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t2_t1_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t2_t1_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t2_t1_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t2_t1_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t2_t1_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t2_t1_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t2_t1_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t2_t1_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t2_t1_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t2_t1_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t2_t1_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t2_t1_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t2_t1_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t2_t1_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t2_t1_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t2_t1_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t2_t1_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t2_t1_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t2_t1_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t2_t1_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t2_t1_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t2_t1_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t2_t1_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t2_t1_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t2_t1_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t2_t1_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t2_t1_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t2_t1_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t2_t1_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t2_t1_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t2_t1_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t2_t1_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t2_t1_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t2_t1_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t2_t1_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t2_t1_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t2_t1_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t2_t1_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t2_t1_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t2_t1_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t2_t1_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t2_t1_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t2_t1_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t2_t1_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t2_t1_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t2_t1_out = { AES_r1_t2_t1_k0, AES_r1_t2_t1_k0, ( AES_r1_t2_t1_k0 ^ AES_r1_t2_t1_k1 ), AES_r1_t2_t1_k1 };
    assign AES_r1_t2_t2_clk = AES_r1_t2_clk;
    assign AES_r1_t2_t2_in = AES_r1_t2_b2;
    assign AES_r1_t2_k2 = AES_r1_t2_t2_out;
    assign AES_r1_t2_t2_s0_clk = AES_r1_t2_t2_clk;
    assign AES_r1_t2_t2_s0_in = AES_r1_t2_t2_in;
    assign AES_r1_t2_t2_k0 = AES_r1_t2_t2_s0_out;
    always @ (  posedge AES_r1_t2_t2_s0_clk)
    begin
        case ( AES_r1_t2_t2_s0_in ) 
        8'h00:
        begin
            AES_r1_t2_t2_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t2_t2_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t2_t2_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t2_t2_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t2_t2_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t2_t2_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t2_t2_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t2_t2_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t2_t2_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t2_t2_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t2_t2_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t2_t2_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t2_t2_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t2_t2_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t2_t2_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t2_t2_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t2_t2_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t2_t2_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t2_t2_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t2_t2_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t2_t2_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t2_t2_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t2_t2_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t2_t2_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t2_t2_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t2_t2_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t2_t2_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t2_t2_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t2_t2_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t2_t2_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t2_t2_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t2_t2_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t2_t2_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t2_t2_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t2_t2_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t2_t2_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t2_t2_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t2_t2_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t2_t2_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t2_t2_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t2_t2_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t2_t2_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t2_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t2_t2_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t2_t2_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t2_t2_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t2_t2_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t2_t2_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t2_t2_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t2_t2_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t2_t2_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t2_t2_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t2_t2_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t2_t2_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t2_t2_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t2_t2_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t2_t2_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t2_t2_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t2_t2_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t2_t2_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t2_t2_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t2_t2_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t2_t2_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t2_t2_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t2_t2_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t2_t2_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t2_t2_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t2_t2_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t2_t2_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t2_t2_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t2_t2_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t2_t2_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t2_t2_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t2_t2_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t2_t2_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t2_t2_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t2_t2_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t2_t2_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t2_t2_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t2_t2_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t2_t2_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t2_t2_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t2_t2_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t2_t2_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t2_t2_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t2_t2_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t2_t2_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t2_t2_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t2_t2_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t2_t2_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t2_t2_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t2_t2_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t2_t2_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t2_t2_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t2_t2_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t2_t2_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t2_t2_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t2_t2_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t2_t2_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t2_t2_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t2_t2_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t2_t2_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t2_t2_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t2_t2_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t2_t2_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t2_t2_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t2_t2_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t2_t2_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t2_t2_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t2_t2_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t2_t2_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t2_t2_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t2_t2_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t2_t2_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t2_t2_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t2_t2_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t2_t2_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t2_t2_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t2_t2_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t2_t2_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t2_t2_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t2_t2_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t2_t2_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t2_t2_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t2_t2_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t2_t2_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t2_t2_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t2_t2_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t2_t2_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t2_t2_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t2_t2_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t2_t2_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t2_t2_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t2_t2_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t2_t2_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t2_t2_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t2_t2_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t2_t2_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t2_t2_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t2_t2_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t2_t2_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t2_t2_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t2_t2_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t2_t2_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t2_t2_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t2_t2_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t2_t2_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t2_t2_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t2_t2_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t2_t2_s4_clk = AES_r1_t2_t2_clk;
    assign AES_r1_t2_t2_s4_in = AES_r1_t2_t2_in;
    assign AES_r1_t2_t2_k1 = AES_r1_t2_t2_s4_out;
    always @ (  posedge AES_r1_t2_t2_s4_clk)
    begin
        case ( AES_r1_t2_t2_s4_in ) 
        8'h00:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t2_t2_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t2_t2_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t2_t2_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t2_t2_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t2_t2_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t2_t2_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t2_t2_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t2_t2_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t2_t2_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t2_t2_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t2_t2_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t2_t2_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t2_t2_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t2_t2_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t2_t2_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t2_t2_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t2_t2_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t2_t2_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t2_t2_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t2_t2_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t2_t2_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t2_t2_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t2_t2_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t2_t2_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t2_t2_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t2_t2_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t2_t2_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t2_t2_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t2_t2_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t2_t2_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t2_t2_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t2_t2_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t2_t2_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t2_t2_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t2_t2_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t2_t2_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t2_t2_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t2_t2_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t2_t2_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t2_t2_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t2_t2_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t2_t2_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t2_t2_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t2_t2_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t2_t2_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t2_t2_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t2_t2_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t2_t2_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t2_t2_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t2_t2_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t2_t2_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t2_t2_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t2_t2_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t2_t2_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t2_t2_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t2_t2_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t2_t2_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t2_t2_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t2_t2_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t2_t2_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t2_t2_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t2_t2_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t2_t2_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t2_t2_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t2_t2_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t2_t2_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t2_t2_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t2_t2_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t2_t2_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t2_t2_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t2_t2_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t2_t2_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t2_t2_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t2_t2_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t2_t2_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t2_t2_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t2_t2_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t2_t2_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t2_t2_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t2_t2_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t2_t2_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t2_t2_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t2_t2_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t2_t2_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t2_t2_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t2_t2_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t2_t2_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t2_t2_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t2_t2_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t2_t2_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t2_t2_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t2_t2_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t2_t2_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t2_t2_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t2_t2_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t2_t2_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t2_t2_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t2_t2_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t2_t2_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t2_t2_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t2_t2_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t2_t2_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t2_t2_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t2_t2_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t2_t2_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t2_t2_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t2_t2_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t2_t2_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t2_t2_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t2_t2_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t2_t2_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t2_t2_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t2_t2_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t2_t2_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t2_t2_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t2_t2_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t2_t2_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t2_t2_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t2_t2_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t2_t2_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t2_t2_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t2_t2_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t2_t2_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t2_t2_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t2_t2_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t2_t2_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t2_t2_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t2_t2_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t2_t2_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t2_t2_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t2_t2_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t2_t2_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t2_t2_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t2_t2_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t2_t2_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t2_t2_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t2_t2_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t2_t2_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t2_t2_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t2_t2_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t2_t2_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t2_t2_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t2_t2_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t2_t2_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t2_t2_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t2_t2_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t2_t2_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t2_t2_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t2_t2_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t2_t2_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t2_t2_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t2_t2_out = { AES_r1_t2_t2_k0, AES_r1_t2_t2_k0, ( AES_r1_t2_t2_k0 ^ AES_r1_t2_t2_k1 ), AES_r1_t2_t2_k1 };
    assign AES_r1_t2_t3_clk = AES_r1_t2_clk;
    assign AES_r1_t2_t3_in = AES_r1_t2_b3;
    assign AES_r1_t2_p3 = AES_r1_t2_t3_out;
    assign AES_r1_t2_t3_s0_clk = AES_r1_t2_t3_clk;
    assign AES_r1_t2_t3_s0_in = AES_r1_t2_t3_in;
    assign AES_r1_t2_t3_k0 = AES_r1_t2_t3_s0_out;
    always @ (  posedge AES_r1_t2_t3_s0_clk)
    begin
        case ( AES_r1_t2_t3_s0_in ) 
        8'h00:
        begin
            AES_r1_t2_t3_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t2_t3_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t2_t3_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t2_t3_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t2_t3_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t2_t3_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t2_t3_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t2_t3_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t2_t3_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t2_t3_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t2_t3_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t2_t3_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t2_t3_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t2_t3_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t2_t3_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t2_t3_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t2_t3_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t2_t3_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t2_t3_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t2_t3_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t2_t3_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t2_t3_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t2_t3_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t2_t3_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t2_t3_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t2_t3_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t2_t3_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t2_t3_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t2_t3_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t2_t3_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t2_t3_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t2_t3_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t2_t3_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t2_t3_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t2_t3_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t2_t3_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t2_t3_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t2_t3_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t2_t3_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t2_t3_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t2_t3_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t2_t3_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t3_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t2_t3_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t2_t3_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t2_t3_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t2_t3_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t2_t3_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t2_t3_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t2_t3_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t2_t3_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t2_t3_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t2_t3_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t2_t3_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t2_t3_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t2_t3_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t2_t3_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t2_t3_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t2_t3_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t2_t3_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t2_t3_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t2_t3_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t2_t3_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t2_t3_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t2_t3_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t2_t3_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t2_t3_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t2_t3_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t2_t3_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t2_t3_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t2_t3_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t2_t3_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t2_t3_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t2_t3_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t2_t3_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t2_t3_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t2_t3_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t2_t3_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t2_t3_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t2_t3_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t2_t3_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t2_t3_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t2_t3_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t2_t3_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t2_t3_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t2_t3_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t2_t3_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t2_t3_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t2_t3_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t2_t3_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t2_t3_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t2_t3_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t2_t3_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t2_t3_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t2_t3_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t2_t3_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t2_t3_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t2_t3_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t2_t3_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t2_t3_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t2_t3_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t2_t3_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t2_t3_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t2_t3_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t2_t3_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t2_t3_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t2_t3_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t2_t3_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t2_t3_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t2_t3_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t2_t3_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t2_t3_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t2_t3_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t2_t3_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t2_t3_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t2_t3_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t2_t3_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t2_t3_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t2_t3_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t2_t3_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t2_t3_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t2_t3_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t2_t3_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t2_t3_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t2_t3_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t2_t3_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t2_t3_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t2_t3_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t2_t3_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t2_t3_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t2_t3_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t2_t3_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t2_t3_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t2_t3_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t2_t3_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t2_t3_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t2_t3_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t2_t3_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t2_t3_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t2_t3_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t2_t3_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t2_t3_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t2_t3_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t2_t3_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t2_t3_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t2_t3_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t2_t3_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t2_t3_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t2_t3_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t2_t3_s4_clk = AES_r1_t2_t3_clk;
    assign AES_r1_t2_t3_s4_in = AES_r1_t2_t3_in;
    assign AES_r1_t2_t3_k1 = AES_r1_t2_t3_s4_out;
    always @ (  posedge AES_r1_t2_t3_s4_clk)
    begin
        case ( AES_r1_t2_t3_s4_in ) 
        8'h00:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t2_t3_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t2_t3_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t2_t3_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t2_t3_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t2_t3_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t2_t3_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t2_t3_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t2_t3_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t2_t3_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t2_t3_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t2_t3_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t2_t3_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t2_t3_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t2_t3_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t2_t3_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t2_t3_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t2_t3_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t2_t3_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t2_t3_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t2_t3_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t2_t3_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t2_t3_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t2_t3_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t2_t3_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t2_t3_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t2_t3_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t2_t3_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t2_t3_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t2_t3_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t2_t3_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t2_t3_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t2_t3_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t2_t3_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t2_t3_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t2_t3_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t2_t3_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t2_t3_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t2_t3_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t2_t3_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t2_t3_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t2_t3_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t2_t3_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t2_t3_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t2_t3_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t2_t3_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t2_t3_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t2_t3_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t2_t3_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t2_t3_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t2_t3_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t2_t3_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t2_t3_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t2_t3_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t2_t3_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t2_t3_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t2_t3_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t2_t3_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t2_t3_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t2_t3_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t2_t3_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t2_t3_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t2_t3_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t2_t3_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t2_t3_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t2_t3_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t2_t3_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t2_t3_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t2_t3_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t2_t3_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t2_t3_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t2_t3_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t2_t3_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t2_t3_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t2_t3_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t2_t3_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t2_t3_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t2_t3_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t2_t3_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t2_t3_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t2_t3_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t2_t3_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t2_t3_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t2_t3_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t2_t3_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t2_t3_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t2_t3_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t2_t3_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t2_t3_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t2_t3_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t2_t3_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t2_t3_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t2_t3_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t2_t3_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t2_t3_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t2_t3_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t2_t3_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t2_t3_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t2_t3_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t2_t3_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t2_t3_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t2_t3_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t2_t3_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t2_t3_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t2_t3_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t2_t3_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t2_t3_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t2_t3_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t2_t3_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t2_t3_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t2_t3_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t2_t3_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t2_t3_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t2_t3_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t2_t3_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t2_t3_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t2_t3_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t2_t3_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t2_t3_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t2_t3_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t2_t3_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t2_t3_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t2_t3_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t2_t3_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t2_t3_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t2_t3_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t2_t3_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t2_t3_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t2_t3_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t2_t3_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t2_t3_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t2_t3_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t2_t3_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t2_t3_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t2_t3_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t2_t3_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t2_t3_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t2_t3_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t2_t3_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t2_t3_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t2_t3_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t2_t3_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t2_t3_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t2_t3_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t2_t3_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t2_t3_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t2_t3_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t2_t3_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t2_t3_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t2_t3_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t2_t3_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t2_t3_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t2_t3_out = { AES_r1_t2_t3_k0, AES_r1_t2_t3_k0, ( AES_r1_t2_t3_k0 ^ AES_r1_t2_t3_k1 ), AES_r1_t2_t3_k1 };
    assign AES_r1_t3_clk = AES_r1_clk;
    assign AES_r1_t3_state = AES_r1_s3;
    assign AES_r1_p30 = AES_r1_t3_p0;
    assign AES_r1_p31 = AES_r1_t3_p1;
    assign AES_r1_p32 = AES_r1_t3_p2;
    assign AES_r1_p33 = AES_r1_t3_p3;
    assign AES_r1_t3_p0 = { AES_r1_t3_k0[7:0], AES_r1_t3_k0[31:8] };
    assign AES_r1_t3_p1 = { AES_r1_t3_k1[15:0], AES_r1_t3_k1[31:16] };
    assign AES_r1_t3_p2 = { AES_r1_t3_k2[23:0], AES_r1_t3_k2[31:24] };
    assign AES_r1_t3_b0 = AES_r1_t3_state[31:24];
    assign AES_r1_t3_b1 = AES_r1_t3_state[23:16];
    assign AES_r1_t3_b2 = AES_r1_t3_state[15:8];
    assign AES_r1_t3_b3 = AES_r1_t3_state[7:0];
    assign AES_r1_t3_t0_clk = AES_r1_t3_clk;
    assign AES_r1_t3_t0_in = AES_r1_t3_b0;
    assign AES_r1_t3_k0 = AES_r1_t3_t0_out;
    assign AES_r1_t3_t0_s0_clk = AES_r1_t3_t0_clk;
    assign AES_r1_t3_t0_s0_in = AES_r1_t3_t0_in;
    assign AES_r1_t3_t0_k0 = AES_r1_t3_t0_s0_out;
    always @ (  posedge AES_r1_t3_t0_s0_clk)
    begin
        case ( AES_r1_t3_t0_s0_in ) 
        8'h00:
        begin
            AES_r1_t3_t0_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t3_t0_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t3_t0_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t3_t0_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t3_t0_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t3_t0_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t3_t0_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t3_t0_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t3_t0_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t3_t0_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t3_t0_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t3_t0_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t3_t0_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t3_t0_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t3_t0_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t3_t0_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t3_t0_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t3_t0_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t3_t0_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t3_t0_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t3_t0_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t3_t0_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t3_t0_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t3_t0_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t3_t0_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t3_t0_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t3_t0_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t3_t0_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t3_t0_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t3_t0_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t3_t0_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t3_t0_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t3_t0_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t3_t0_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t3_t0_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t3_t0_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t3_t0_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t3_t0_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t3_t0_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t3_t0_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t3_t0_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t3_t0_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t0_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t3_t0_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t3_t0_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t3_t0_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t3_t0_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t3_t0_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t3_t0_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t3_t0_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t3_t0_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t3_t0_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t3_t0_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t3_t0_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t3_t0_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t3_t0_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t3_t0_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t3_t0_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t3_t0_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t3_t0_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t3_t0_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t3_t0_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t3_t0_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t3_t0_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t3_t0_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t3_t0_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t3_t0_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t3_t0_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t3_t0_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t3_t0_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t3_t0_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t3_t0_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t3_t0_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t3_t0_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t3_t0_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t3_t0_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t3_t0_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t3_t0_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t3_t0_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t3_t0_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t3_t0_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t3_t0_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t3_t0_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t3_t0_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t3_t0_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t3_t0_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t3_t0_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t3_t0_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t3_t0_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t3_t0_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t3_t0_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t3_t0_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t3_t0_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t3_t0_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t3_t0_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t3_t0_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t3_t0_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t3_t0_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t3_t0_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t3_t0_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t3_t0_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t3_t0_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t3_t0_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t3_t0_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t3_t0_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t3_t0_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t3_t0_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t3_t0_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t3_t0_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t3_t0_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t3_t0_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t3_t0_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t3_t0_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t3_t0_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t3_t0_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t3_t0_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t3_t0_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t3_t0_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t3_t0_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t3_t0_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t3_t0_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t3_t0_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t3_t0_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t3_t0_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t3_t0_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t3_t0_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t3_t0_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t3_t0_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t3_t0_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t3_t0_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t3_t0_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t3_t0_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t3_t0_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t3_t0_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t3_t0_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t3_t0_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t3_t0_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t3_t0_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t3_t0_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t3_t0_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t3_t0_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t3_t0_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t3_t0_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t3_t0_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t3_t0_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t3_t0_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t3_t0_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t3_t0_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t3_t0_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t3_t0_s4_clk = AES_r1_t3_t0_clk;
    assign AES_r1_t3_t0_s4_in = AES_r1_t3_t0_in;
    assign AES_r1_t3_t0_k1 = AES_r1_t3_t0_s4_out;
    always @ (  posedge AES_r1_t3_t0_s4_clk)
    begin
        case ( AES_r1_t3_t0_s4_in ) 
        8'h00:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t3_t0_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t3_t0_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t3_t0_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t3_t0_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t3_t0_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t3_t0_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t3_t0_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t3_t0_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t3_t0_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t3_t0_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t3_t0_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t3_t0_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t3_t0_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t3_t0_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t3_t0_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t3_t0_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t3_t0_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t3_t0_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t3_t0_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t3_t0_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t3_t0_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t3_t0_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t3_t0_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t3_t0_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t3_t0_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t3_t0_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t3_t0_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t3_t0_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t3_t0_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t3_t0_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t3_t0_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t3_t0_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t3_t0_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t3_t0_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t3_t0_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t3_t0_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t3_t0_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t3_t0_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t3_t0_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t3_t0_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t3_t0_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t3_t0_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t3_t0_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t3_t0_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t3_t0_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t3_t0_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t3_t0_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t3_t0_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t3_t0_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t3_t0_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t3_t0_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t3_t0_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t3_t0_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t3_t0_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t3_t0_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t3_t0_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t3_t0_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t3_t0_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t3_t0_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t3_t0_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t3_t0_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t3_t0_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t3_t0_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t3_t0_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t3_t0_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t3_t0_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t3_t0_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t3_t0_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t3_t0_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t3_t0_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t3_t0_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t3_t0_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t3_t0_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t3_t0_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t3_t0_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t3_t0_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t3_t0_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t3_t0_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t3_t0_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t3_t0_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t3_t0_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t3_t0_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t3_t0_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t3_t0_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t3_t0_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t3_t0_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t3_t0_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t3_t0_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t3_t0_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t3_t0_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t3_t0_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t3_t0_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t3_t0_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t3_t0_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t3_t0_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t3_t0_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t3_t0_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t3_t0_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t3_t0_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t3_t0_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t3_t0_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t3_t0_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t3_t0_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t3_t0_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t3_t0_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t3_t0_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t3_t0_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t3_t0_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t3_t0_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t3_t0_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t3_t0_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t3_t0_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t3_t0_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t3_t0_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t3_t0_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t3_t0_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t3_t0_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t3_t0_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t3_t0_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t3_t0_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t3_t0_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t3_t0_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t3_t0_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t3_t0_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t3_t0_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t3_t0_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t3_t0_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t3_t0_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t3_t0_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t3_t0_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t3_t0_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t3_t0_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t3_t0_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t3_t0_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t3_t0_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t3_t0_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t3_t0_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t3_t0_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t3_t0_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t3_t0_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t3_t0_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t3_t0_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t3_t0_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t3_t0_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t3_t0_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t3_t0_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t3_t0_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t3_t0_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t3_t0_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t3_t0_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t3_t0_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t3_t0_out = { AES_r1_t3_t0_k0, AES_r1_t3_t0_k0, ( AES_r1_t3_t0_k0 ^ AES_r1_t3_t0_k1 ), AES_r1_t3_t0_k1 };
    assign AES_r1_t3_t1_clk = AES_r1_t3_clk;
    assign AES_r1_t3_t1_in = AES_r1_t3_b1;
    assign AES_r1_t3_k1 = AES_r1_t3_t1_out;
    assign AES_r1_t3_t1_s0_clk = AES_r1_t3_t1_clk;
    assign AES_r1_t3_t1_s0_in = AES_r1_t3_t1_in;
    assign AES_r1_t3_t1_k0 = AES_r1_t3_t1_s0_out;
    always @ (  posedge AES_r1_t3_t1_s0_clk)
    begin
        case ( AES_r1_t3_t1_s0_in ) 
        8'h00:
        begin
            AES_r1_t3_t1_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t3_t1_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t3_t1_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t3_t1_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t3_t1_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t3_t1_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t3_t1_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t3_t1_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t3_t1_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t3_t1_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t3_t1_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t3_t1_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t3_t1_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t3_t1_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t3_t1_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t3_t1_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t3_t1_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t3_t1_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t3_t1_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t3_t1_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t3_t1_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t3_t1_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t3_t1_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t3_t1_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t3_t1_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t3_t1_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t3_t1_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t3_t1_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t3_t1_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t3_t1_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t3_t1_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t3_t1_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t3_t1_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t3_t1_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t3_t1_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t3_t1_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t3_t1_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t3_t1_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t3_t1_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t3_t1_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t3_t1_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t3_t1_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t1_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t3_t1_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t3_t1_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t3_t1_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t3_t1_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t3_t1_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t3_t1_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t3_t1_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t3_t1_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t3_t1_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t3_t1_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t3_t1_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t3_t1_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t3_t1_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t3_t1_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t3_t1_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t3_t1_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t3_t1_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t3_t1_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t3_t1_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t3_t1_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t3_t1_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t3_t1_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t3_t1_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t3_t1_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t3_t1_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t3_t1_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t3_t1_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t3_t1_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t3_t1_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t3_t1_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t3_t1_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t3_t1_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t3_t1_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t3_t1_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t3_t1_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t3_t1_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t3_t1_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t3_t1_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t3_t1_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t3_t1_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t3_t1_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t3_t1_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t3_t1_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t3_t1_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t3_t1_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t3_t1_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t3_t1_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t3_t1_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t3_t1_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t3_t1_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t3_t1_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t3_t1_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t3_t1_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t3_t1_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t3_t1_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t3_t1_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t3_t1_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t3_t1_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t3_t1_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t3_t1_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t3_t1_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t3_t1_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t3_t1_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t3_t1_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t3_t1_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t3_t1_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t3_t1_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t3_t1_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t3_t1_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t3_t1_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t3_t1_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t3_t1_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t3_t1_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t3_t1_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t3_t1_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t3_t1_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t3_t1_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t3_t1_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t3_t1_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t3_t1_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t3_t1_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t3_t1_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t3_t1_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t3_t1_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t3_t1_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t3_t1_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t3_t1_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t3_t1_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t3_t1_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t3_t1_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t3_t1_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t3_t1_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t3_t1_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t3_t1_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t3_t1_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t3_t1_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t3_t1_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t3_t1_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t3_t1_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t3_t1_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t3_t1_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t3_t1_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t3_t1_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t3_t1_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t3_t1_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t3_t1_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t3_t1_s4_clk = AES_r1_t3_t1_clk;
    assign AES_r1_t3_t1_s4_in = AES_r1_t3_t1_in;
    assign AES_r1_t3_t1_k1 = AES_r1_t3_t1_s4_out;
    always @ (  posedge AES_r1_t3_t1_s4_clk)
    begin
        case ( AES_r1_t3_t1_s4_in ) 
        8'h00:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t3_t1_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t3_t1_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t3_t1_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t3_t1_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t3_t1_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t3_t1_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t3_t1_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t3_t1_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t3_t1_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t3_t1_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t3_t1_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t3_t1_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t3_t1_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t3_t1_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t3_t1_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t3_t1_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t3_t1_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t3_t1_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t3_t1_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t3_t1_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t3_t1_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t3_t1_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t3_t1_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t3_t1_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t3_t1_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t3_t1_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t3_t1_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t3_t1_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t3_t1_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t3_t1_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t3_t1_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t3_t1_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t3_t1_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t3_t1_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t3_t1_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t3_t1_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t3_t1_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t3_t1_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t3_t1_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t3_t1_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t3_t1_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t3_t1_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t3_t1_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t3_t1_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t3_t1_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t3_t1_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t3_t1_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t3_t1_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t3_t1_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t3_t1_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t3_t1_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t3_t1_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t3_t1_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t3_t1_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t3_t1_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t3_t1_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t3_t1_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t3_t1_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t3_t1_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t3_t1_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t3_t1_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t3_t1_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t3_t1_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t3_t1_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t3_t1_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t3_t1_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t3_t1_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t3_t1_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t3_t1_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t3_t1_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t3_t1_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t3_t1_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t3_t1_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t3_t1_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t3_t1_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t3_t1_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t3_t1_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t3_t1_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t3_t1_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t3_t1_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t3_t1_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t3_t1_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t3_t1_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t3_t1_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t3_t1_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t3_t1_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t3_t1_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t3_t1_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t3_t1_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t3_t1_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t3_t1_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t3_t1_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t3_t1_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t3_t1_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t3_t1_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t3_t1_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t3_t1_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t3_t1_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t3_t1_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t3_t1_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t3_t1_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t3_t1_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t3_t1_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t3_t1_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t3_t1_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t3_t1_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t3_t1_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t3_t1_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t3_t1_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t3_t1_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t3_t1_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t3_t1_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t3_t1_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t3_t1_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t3_t1_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t3_t1_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t3_t1_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t3_t1_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t3_t1_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t3_t1_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t3_t1_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t3_t1_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t3_t1_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t3_t1_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t3_t1_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t3_t1_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t3_t1_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t3_t1_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t3_t1_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t3_t1_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t3_t1_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t3_t1_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t3_t1_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t3_t1_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t3_t1_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t3_t1_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t3_t1_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t3_t1_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t3_t1_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t3_t1_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t3_t1_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t3_t1_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t3_t1_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t3_t1_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t3_t1_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t3_t1_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t3_t1_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t3_t1_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t3_t1_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t3_t1_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t3_t1_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t3_t1_out = { AES_r1_t3_t1_k0, AES_r1_t3_t1_k0, ( AES_r1_t3_t1_k0 ^ AES_r1_t3_t1_k1 ), AES_r1_t3_t1_k1 };
    assign AES_r1_t3_t2_clk = AES_r1_t3_clk;
    assign AES_r1_t3_t2_in = AES_r1_t3_b2;
    assign AES_r1_t3_k2 = AES_r1_t3_t2_out;
    assign AES_r1_t3_t2_s0_clk = AES_r1_t3_t2_clk;
    assign AES_r1_t3_t2_s0_in = AES_r1_t3_t2_in;
    assign AES_r1_t3_t2_k0 = AES_r1_t3_t2_s0_out;
    always @ (  posedge AES_r1_t3_t2_s0_clk)
    begin
        case ( AES_r1_t3_t2_s0_in ) 
        8'h00:
        begin
            AES_r1_t3_t2_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t3_t2_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t3_t2_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t3_t2_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t3_t2_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t3_t2_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t3_t2_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t3_t2_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t3_t2_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t3_t2_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t3_t2_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t3_t2_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t3_t2_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t3_t2_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t3_t2_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t3_t2_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t3_t2_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t3_t2_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t3_t2_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t3_t2_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t3_t2_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t3_t2_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t3_t2_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t3_t2_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t3_t2_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t3_t2_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t3_t2_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t3_t2_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t3_t2_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t3_t2_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t3_t2_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t3_t2_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t3_t2_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t3_t2_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t3_t2_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t3_t2_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t3_t2_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t3_t2_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t3_t2_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t3_t2_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t3_t2_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t3_t2_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t2_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t3_t2_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t3_t2_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t3_t2_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t3_t2_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t3_t2_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t3_t2_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t3_t2_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t3_t2_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t3_t2_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t3_t2_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t3_t2_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t3_t2_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t3_t2_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t3_t2_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t3_t2_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t3_t2_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t3_t2_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t3_t2_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t3_t2_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t3_t2_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t3_t2_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t3_t2_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t3_t2_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t3_t2_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t3_t2_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t3_t2_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t3_t2_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t3_t2_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t3_t2_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t3_t2_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t3_t2_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t3_t2_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t3_t2_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t3_t2_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t3_t2_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t3_t2_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t3_t2_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t3_t2_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t3_t2_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t3_t2_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t3_t2_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t3_t2_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t3_t2_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t3_t2_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t3_t2_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t3_t2_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t3_t2_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t3_t2_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t3_t2_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t3_t2_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t3_t2_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t3_t2_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t3_t2_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t3_t2_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t3_t2_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t3_t2_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t3_t2_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t3_t2_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t3_t2_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t3_t2_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t3_t2_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t3_t2_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t3_t2_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t3_t2_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t3_t2_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t3_t2_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t3_t2_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t3_t2_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t3_t2_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t3_t2_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t3_t2_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t3_t2_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t3_t2_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t3_t2_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t3_t2_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t3_t2_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t3_t2_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t3_t2_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t3_t2_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t3_t2_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t3_t2_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t3_t2_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t3_t2_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t3_t2_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t3_t2_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t3_t2_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t3_t2_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t3_t2_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t3_t2_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t3_t2_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t3_t2_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t3_t2_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t3_t2_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t3_t2_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t3_t2_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t3_t2_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t3_t2_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t3_t2_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t3_t2_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t3_t2_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t3_t2_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t3_t2_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t3_t2_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t3_t2_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t3_t2_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t3_t2_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t3_t2_s4_clk = AES_r1_t3_t2_clk;
    assign AES_r1_t3_t2_s4_in = AES_r1_t3_t2_in;
    assign AES_r1_t3_t2_k1 = AES_r1_t3_t2_s4_out;
    always @ (  posedge AES_r1_t3_t2_s4_clk)
    begin
        case ( AES_r1_t3_t2_s4_in ) 
        8'h00:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t3_t2_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t3_t2_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t3_t2_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t3_t2_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t3_t2_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t3_t2_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t3_t2_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t3_t2_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t3_t2_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t3_t2_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t3_t2_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t3_t2_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t3_t2_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t3_t2_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t3_t2_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t3_t2_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t3_t2_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t3_t2_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t3_t2_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t3_t2_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t3_t2_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t3_t2_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t3_t2_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t3_t2_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t3_t2_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t3_t2_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t3_t2_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t3_t2_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t3_t2_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t3_t2_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t3_t2_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t3_t2_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t3_t2_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t3_t2_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t3_t2_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t3_t2_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t3_t2_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t3_t2_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t3_t2_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t3_t2_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t3_t2_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t3_t2_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t3_t2_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t3_t2_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t3_t2_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t3_t2_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t3_t2_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t3_t2_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t3_t2_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t3_t2_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t3_t2_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t3_t2_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t3_t2_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t3_t2_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t3_t2_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t3_t2_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t3_t2_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t3_t2_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t3_t2_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t3_t2_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t3_t2_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t3_t2_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t3_t2_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t3_t2_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t3_t2_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t3_t2_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t3_t2_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t3_t2_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t3_t2_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t3_t2_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t3_t2_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t3_t2_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t3_t2_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t3_t2_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t3_t2_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t3_t2_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t3_t2_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t3_t2_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t3_t2_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t3_t2_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t3_t2_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t3_t2_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t3_t2_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t3_t2_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t3_t2_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t3_t2_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t3_t2_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t3_t2_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t3_t2_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t3_t2_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t3_t2_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t3_t2_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t3_t2_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t3_t2_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t3_t2_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t3_t2_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t3_t2_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t3_t2_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t3_t2_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t3_t2_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t3_t2_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t3_t2_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t3_t2_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t3_t2_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t3_t2_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t3_t2_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t3_t2_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t3_t2_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t3_t2_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t3_t2_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t3_t2_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t3_t2_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t3_t2_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t3_t2_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t3_t2_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t3_t2_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t3_t2_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t3_t2_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t3_t2_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t3_t2_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t3_t2_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t3_t2_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t3_t2_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t3_t2_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t3_t2_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t3_t2_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t3_t2_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t3_t2_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t3_t2_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t3_t2_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t3_t2_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t3_t2_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t3_t2_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t3_t2_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t3_t2_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t3_t2_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t3_t2_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t3_t2_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t3_t2_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t3_t2_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t3_t2_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t3_t2_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t3_t2_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t3_t2_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t3_t2_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t3_t2_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t3_t2_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t3_t2_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t3_t2_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t3_t2_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t3_t2_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t3_t2_out = { AES_r1_t3_t2_k0, AES_r1_t3_t2_k0, ( AES_r1_t3_t2_k0 ^ AES_r1_t3_t2_k1 ), AES_r1_t3_t2_k1 };
    assign AES_r1_t3_t3_clk = AES_r1_t3_clk;
    assign AES_r1_t3_t3_in = AES_r1_t3_b3;
    assign AES_r1_t3_p3 = AES_r1_t3_t3_out;
    assign AES_r1_t3_t3_s0_clk = AES_r1_t3_t3_clk;
    assign AES_r1_t3_t3_s0_in = AES_r1_t3_t3_in;
    assign AES_r1_t3_t3_k0 = AES_r1_t3_t3_s0_out;
    always @ (  posedge AES_r1_t3_t3_s0_clk)
    begin
        case ( AES_r1_t3_t3_s0_in ) 
        8'h00:
        begin
            AES_r1_t3_t3_s0_out <= 8'h63;
        end
        8'h01:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7c;
        end
        8'h02:
        begin
            AES_r1_t3_t3_s0_out <= 8'h77;
        end
        8'h03:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7b;
        end
        8'h04:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf2;
        end
        8'h05:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6b;
        end
        8'h06:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6f;
        end
        8'h07:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc5;
        end
        8'h08:
        begin
            AES_r1_t3_t3_s0_out <= 8'h30;
        end
        8'h09:
        begin
            AES_r1_t3_t3_s0_out <= 8'h01;
        end
        8'h0a:
        begin
            AES_r1_t3_t3_s0_out <= 8'h67;
        end
        8'h0b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2b;
        end
        8'h0c:
        begin
            AES_r1_t3_t3_s0_out <= 8'hfe;
        end
        8'h0d:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd7;
        end
        8'h0e:
        begin
            AES_r1_t3_t3_s0_out <= 8'hab;
        end
        8'h0f:
        begin
            AES_r1_t3_t3_s0_out <= 8'h76;
        end
        8'h10:
        begin
            AES_r1_t3_t3_s0_out <= 8'hca;
        end
        8'h11:
        begin
            AES_r1_t3_t3_s0_out <= 8'h82;
        end
        8'h12:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc9;
        end
        8'h13:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7d;
        end
        8'h14:
        begin
            AES_r1_t3_t3_s0_out <= 8'hfa;
        end
        8'h15:
        begin
            AES_r1_t3_t3_s0_out <= 8'h59;
        end
        8'h16:
        begin
            AES_r1_t3_t3_s0_out <= 8'h47;
        end
        8'h17:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf0;
        end
        8'h18:
        begin
            AES_r1_t3_t3_s0_out <= 8'had;
        end
        8'h19:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd4;
        end
        8'h1a:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha2;
        end
        8'h1b:
        begin
            AES_r1_t3_t3_s0_out <= 8'haf;
        end
        8'h1c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9c;
        end
        8'h1d:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha4;
        end
        8'h1e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h72;
        end
        8'h1f:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc0;
        end
        8'h20:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb7;
        end
        8'h21:
        begin
            AES_r1_t3_t3_s0_out <= 8'hfd;
        end
        8'h22:
        begin
            AES_r1_t3_t3_s0_out <= 8'h93;
        end
        8'h23:
        begin
            AES_r1_t3_t3_s0_out <= 8'h26;
        end
        8'h24:
        begin
            AES_r1_t3_t3_s0_out <= 8'h36;
        end
        8'h25:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3f;
        end
        8'h26:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf7;
        end
        8'h27:
        begin
            AES_r1_t3_t3_s0_out <= 8'hcc;
        end
        8'h28:
        begin
            AES_r1_t3_t3_s0_out <= 8'h34;
        end
        8'h29:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha5;
        end
        8'h2a:
        begin
            AES_r1_t3_t3_s0_out <= 8'he5;
        end
        8'h2b:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf1;
        end
        8'h2c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h71;
        end
        8'h2d:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd8;
        end
        8'h2e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h31;
        end
        8'h2f:
        begin
            AES_r1_t3_t3_s0_out <= 8'h15;
        end
        8'h30:
        begin
            AES_r1_t3_t3_s0_out <= 8'h04;
        end
        8'h31:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc7;
        end
        8'h32:
        begin
            AES_r1_t3_t3_s0_out <= 8'h23;
        end
        8'h33:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc3;
        end
        8'h34:
        begin
            AES_r1_t3_t3_s0_out <= 8'h18;
        end
        8'h35:
        begin
            AES_r1_t3_t3_s0_out <= 8'h96;
        end
        8'h36:
        begin
            AES_r1_t3_t3_s0_out <= 8'h05;
        end
        8'h37:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9a;
        end
        8'h38:
        begin
            AES_r1_t3_t3_s0_out <= 8'h07;
        end
        8'h39:
        begin
            AES_r1_t3_t3_s0_out <= 8'h12;
        end
        8'h3a:
        begin
            AES_r1_t3_t3_s0_out <= 8'h80;
        end
        8'h3b:
        begin
            AES_r1_t3_t3_s0_out <= 8'he2;
        end
        8'h3c:
        begin
            AES_r1_t3_t3_s0_out <= 8'heb;
        end
        8'h3d:
        begin
            AES_r1_t3_t3_s0_out <= 8'h27;
        end
        8'h3e:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb2;
        end
        8'h3f:
        begin
            AES_r1_t3_t3_s0_out <= 8'h75;
        end
        8'h40:
        begin
            AES_r1_t3_t3_s0_out <= 8'h09;
        end
        8'h41:
        begin
            AES_r1_t3_t3_s0_out <= 8'h83;
        end
        8'h42:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2c;
        end
        8'h43:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1a;
        end
        8'h44:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1b;
        end
        8'h45:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6e;
        end
        8'h46:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5a;
        end
        8'h47:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha0;
        end
        8'h48:
        begin
            AES_r1_t3_t3_s0_out <= 8'h52;
        end
        8'h49:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3b;
        end
        8'h4a:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd6;
        end
        8'h4b:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb3;
        end
        8'h4c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h29;
        end
        8'h4d:
        begin
            AES_r1_t3_t3_s0_out <= 8'he3;
        end
        8'h4e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2f;
        end
        8'h4f:
        begin
            AES_r1_t3_t3_s0_out <= 8'h84;
        end
        8'h50:
        begin
            AES_r1_t3_t3_s0_out <= 8'h53;
        end
        8'h51:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd1;
        end
        8'h52:
        begin
            AES_r1_t3_t3_s0_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t3_s0_out <= 8'hed;
        end
        8'h54:
        begin
            AES_r1_t3_t3_s0_out <= 8'h20;
        end
        8'h55:
        begin
            AES_r1_t3_t3_s0_out <= 8'hfc;
        end
        8'h56:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb1;
        end
        8'h57:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5b;
        end
        8'h58:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6a;
        end
        8'h59:
        begin
            AES_r1_t3_t3_s0_out <= 8'hcb;
        end
        8'h5a:
        begin
            AES_r1_t3_t3_s0_out <= 8'hbe;
        end
        8'h5b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h39;
        end
        8'h5c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4a;
        end
        8'h5d:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4c;
        end
        8'h5e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h58;
        end
        8'h5f:
        begin
            AES_r1_t3_t3_s0_out <= 8'hcf;
        end
        8'h60:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd0;
        end
        8'h61:
        begin
            AES_r1_t3_t3_s0_out <= 8'hef;
        end
        8'h62:
        begin
            AES_r1_t3_t3_s0_out <= 8'haa;
        end
        8'h63:
        begin
            AES_r1_t3_t3_s0_out <= 8'hfb;
        end
        8'h64:
        begin
            AES_r1_t3_t3_s0_out <= 8'h43;
        end
        8'h65:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4d;
        end
        8'h66:
        begin
            AES_r1_t3_t3_s0_out <= 8'h33;
        end
        8'h67:
        begin
            AES_r1_t3_t3_s0_out <= 8'h85;
        end
        8'h68:
        begin
            AES_r1_t3_t3_s0_out <= 8'h45;
        end
        8'h69:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf9;
        end
        8'h6a:
        begin
            AES_r1_t3_t3_s0_out <= 8'h02;
        end
        8'h6b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7f;
        end
        8'h6c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h50;
        end
        8'h6d:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3c;
        end
        8'h6e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9f;
        end
        8'h6f:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha8;
        end
        8'h70:
        begin
            AES_r1_t3_t3_s0_out <= 8'h51;
        end
        8'h71:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha3;
        end
        8'h72:
        begin
            AES_r1_t3_t3_s0_out <= 8'h40;
        end
        8'h73:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8f;
        end
        8'h74:
        begin
            AES_r1_t3_t3_s0_out <= 8'h92;
        end
        8'h75:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9d;
        end
        8'h76:
        begin
            AES_r1_t3_t3_s0_out <= 8'h38;
        end
        8'h77:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf5;
        end
        8'h78:
        begin
            AES_r1_t3_t3_s0_out <= 8'hbc;
        end
        8'h79:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb6;
        end
        8'h7a:
        begin
            AES_r1_t3_t3_s0_out <= 8'hda;
        end
        8'h7b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h21;
        end
        8'h7c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h10;
        end
        8'h7d:
        begin
            AES_r1_t3_t3_s0_out <= 8'hff;
        end
        8'h7e:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf3;
        end
        8'h7f:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd2;
        end
        8'h80:
        begin
            AES_r1_t3_t3_s0_out <= 8'hcd;
        end
        8'h81:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0c;
        end
        8'h82:
        begin
            AES_r1_t3_t3_s0_out <= 8'h13;
        end
        8'h83:
        begin
            AES_r1_t3_t3_s0_out <= 8'hec;
        end
        8'h84:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5f;
        end
        8'h85:
        begin
            AES_r1_t3_t3_s0_out <= 8'h97;
        end
        8'h86:
        begin
            AES_r1_t3_t3_s0_out <= 8'h44;
        end
        8'h87:
        begin
            AES_r1_t3_t3_s0_out <= 8'h17;
        end
        8'h88:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc4;
        end
        8'h89:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha7;
        end
        8'h8a:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7e;
        end
        8'h8b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3d;
        end
        8'h8c:
        begin
            AES_r1_t3_t3_s0_out <= 8'h64;
        end
        8'h8d:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5d;
        end
        8'h8e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h19;
        end
        8'h8f:
        begin
            AES_r1_t3_t3_s0_out <= 8'h73;
        end
        8'h90:
        begin
            AES_r1_t3_t3_s0_out <= 8'h60;
        end
        8'h91:
        begin
            AES_r1_t3_t3_s0_out <= 8'h81;
        end
        8'h92:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4f;
        end
        8'h93:
        begin
            AES_r1_t3_t3_s0_out <= 8'hdc;
        end
        8'h94:
        begin
            AES_r1_t3_t3_s0_out <= 8'h22;
        end
        8'h95:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2a;
        end
        8'h96:
        begin
            AES_r1_t3_t3_s0_out <= 8'h90;
        end
        8'h97:
        begin
            AES_r1_t3_t3_s0_out <= 8'h88;
        end
        8'h98:
        begin
            AES_r1_t3_t3_s0_out <= 8'h46;
        end
        8'h99:
        begin
            AES_r1_t3_t3_s0_out <= 8'hee;
        end
        8'h9a:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb8;
        end
        8'h9b:
        begin
            AES_r1_t3_t3_s0_out <= 8'h14;
        end
        8'h9c:
        begin
            AES_r1_t3_t3_s0_out <= 8'hde;
        end
        8'h9d:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5e;
        end
        8'h9e:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0b;
        end
        8'h9f:
        begin
            AES_r1_t3_t3_s0_out <= 8'hdb;
        end
        8'ha0:
        begin
            AES_r1_t3_t3_s0_out <= 8'he0;
        end
        8'ha1:
        begin
            AES_r1_t3_t3_s0_out <= 8'h32;
        end
        8'ha2:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3a;
        end
        8'ha3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0a;
        end
        8'ha4:
        begin
            AES_r1_t3_t3_s0_out <= 8'h49;
        end
        8'ha5:
        begin
            AES_r1_t3_t3_s0_out <= 8'h06;
        end
        8'ha6:
        begin
            AES_r1_t3_t3_s0_out <= 8'h24;
        end
        8'ha7:
        begin
            AES_r1_t3_t3_s0_out <= 8'h5c;
        end
        8'ha8:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc2;
        end
        8'ha9:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd3;
        end
        8'haa:
        begin
            AES_r1_t3_t3_s0_out <= 8'hac;
        end
        8'hab:
        begin
            AES_r1_t3_t3_s0_out <= 8'h62;
        end
        8'hac:
        begin
            AES_r1_t3_t3_s0_out <= 8'h91;
        end
        8'had:
        begin
            AES_r1_t3_t3_s0_out <= 8'h95;
        end
        8'hae:
        begin
            AES_r1_t3_t3_s0_out <= 8'he4;
        end
        8'haf:
        begin
            AES_r1_t3_t3_s0_out <= 8'h79;
        end
        8'hb0:
        begin
            AES_r1_t3_t3_s0_out <= 8'he7;
        end
        8'hb1:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc8;
        end
        8'hb2:
        begin
            AES_r1_t3_t3_s0_out <= 8'h37;
        end
        8'hb3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6d;
        end
        8'hb4:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8d;
        end
        8'hb5:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd5;
        end
        8'hb6:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4e;
        end
        8'hb7:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha9;
        end
        8'hb8:
        begin
            AES_r1_t3_t3_s0_out <= 8'h6c;
        end
        8'hb9:
        begin
            AES_r1_t3_t3_s0_out <= 8'h56;
        end
        8'hba:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf4;
        end
        8'hbb:
        begin
            AES_r1_t3_t3_s0_out <= 8'hea;
        end
        8'hbc:
        begin
            AES_r1_t3_t3_s0_out <= 8'h65;
        end
        8'hbd:
        begin
            AES_r1_t3_t3_s0_out <= 8'h7a;
        end
        8'hbe:
        begin
            AES_r1_t3_t3_s0_out <= 8'hae;
        end
        8'hbf:
        begin
            AES_r1_t3_t3_s0_out <= 8'h08;
        end
        8'hc0:
        begin
            AES_r1_t3_t3_s0_out <= 8'hba;
        end
        8'hc1:
        begin
            AES_r1_t3_t3_s0_out <= 8'h78;
        end
        8'hc2:
        begin
            AES_r1_t3_t3_s0_out <= 8'h25;
        end
        8'hc3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2e;
        end
        8'hc4:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1c;
        end
        8'hc5:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha6;
        end
        8'hc6:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb4;
        end
        8'hc7:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc6;
        end
        8'hc8:
        begin
            AES_r1_t3_t3_s0_out <= 8'he8;
        end
        8'hc9:
        begin
            AES_r1_t3_t3_s0_out <= 8'hdd;
        end
        8'hca:
        begin
            AES_r1_t3_t3_s0_out <= 8'h74;
        end
        8'hcb:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1f;
        end
        8'hcc:
        begin
            AES_r1_t3_t3_s0_out <= 8'h4b;
        end
        8'hcd:
        begin
            AES_r1_t3_t3_s0_out <= 8'hbd;
        end
        8'hce:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8b;
        end
        8'hcf:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8a;
        end
        8'hd0:
        begin
            AES_r1_t3_t3_s0_out <= 8'h70;
        end
        8'hd1:
        begin
            AES_r1_t3_t3_s0_out <= 8'h3e;
        end
        8'hd2:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb5;
        end
        8'hd3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h66;
        end
        8'hd4:
        begin
            AES_r1_t3_t3_s0_out <= 8'h48;
        end
        8'hd5:
        begin
            AES_r1_t3_t3_s0_out <= 8'h03;
        end
        8'hd6:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf6;
        end
        8'hd7:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0e;
        end
        8'hd8:
        begin
            AES_r1_t3_t3_s0_out <= 8'h61;
        end
        8'hd9:
        begin
            AES_r1_t3_t3_s0_out <= 8'h35;
        end
        8'hda:
        begin
            AES_r1_t3_t3_s0_out <= 8'h57;
        end
        8'hdb:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb9;
        end
        8'hdc:
        begin
            AES_r1_t3_t3_s0_out <= 8'h86;
        end
        8'hdd:
        begin
            AES_r1_t3_t3_s0_out <= 8'hc1;
        end
        8'hde:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1d;
        end
        8'hdf:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9e;
        end
        8'he0:
        begin
            AES_r1_t3_t3_s0_out <= 8'he1;
        end
        8'he1:
        begin
            AES_r1_t3_t3_s0_out <= 8'hf8;
        end
        8'he2:
        begin
            AES_r1_t3_t3_s0_out <= 8'h98;
        end
        8'he3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h11;
        end
        8'he4:
        begin
            AES_r1_t3_t3_s0_out <= 8'h69;
        end
        8'he5:
        begin
            AES_r1_t3_t3_s0_out <= 8'hd9;
        end
        8'he6:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8e;
        end
        8'he7:
        begin
            AES_r1_t3_t3_s0_out <= 8'h94;
        end
        8'he8:
        begin
            AES_r1_t3_t3_s0_out <= 8'h9b;
        end
        8'he9:
        begin
            AES_r1_t3_t3_s0_out <= 8'h1e;
        end
        8'hea:
        begin
            AES_r1_t3_t3_s0_out <= 8'h87;
        end
        8'heb:
        begin
            AES_r1_t3_t3_s0_out <= 8'he9;
        end
        8'hec:
        begin
            AES_r1_t3_t3_s0_out <= 8'hce;
        end
        8'hed:
        begin
            AES_r1_t3_t3_s0_out <= 8'h55;
        end
        8'hee:
        begin
            AES_r1_t3_t3_s0_out <= 8'h28;
        end
        8'hef:
        begin
            AES_r1_t3_t3_s0_out <= 8'hdf;
        end
        8'hf0:
        begin
            AES_r1_t3_t3_s0_out <= 8'h8c;
        end
        8'hf1:
        begin
            AES_r1_t3_t3_s0_out <= 8'ha1;
        end
        8'hf2:
        begin
            AES_r1_t3_t3_s0_out <= 8'h89;
        end
        8'hf3:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0d;
        end
        8'hf4:
        begin
            AES_r1_t3_t3_s0_out <= 8'hbf;
        end
        8'hf5:
        begin
            AES_r1_t3_t3_s0_out <= 8'he6;
        end
        8'hf6:
        begin
            AES_r1_t3_t3_s0_out <= 8'h42;
        end
        8'hf7:
        begin
            AES_r1_t3_t3_s0_out <= 8'h68;
        end
        8'hf8:
        begin
            AES_r1_t3_t3_s0_out <= 8'h41;
        end
        8'hf9:
        begin
            AES_r1_t3_t3_s0_out <= 8'h99;
        end
        8'hfa:
        begin
            AES_r1_t3_t3_s0_out <= 8'h2d;
        end
        8'hfb:
        begin
            AES_r1_t3_t3_s0_out <= 8'h0f;
        end
        8'hfc:
        begin
            AES_r1_t3_t3_s0_out <= 8'hb0;
        end
        8'hfd:
        begin
            AES_r1_t3_t3_s0_out <= 8'h54;
        end
        8'hfe:
        begin
            AES_r1_t3_t3_s0_out <= 8'hbb;
        end
        8'hff:
        begin
            AES_r1_t3_t3_s0_out <= 8'h16;
        end
        endcase
    end
    assign AES_r1_t3_t3_s4_clk = AES_r1_t3_t3_clk;
    assign AES_r1_t3_t3_s4_in = AES_r1_t3_t3_in;
    assign AES_r1_t3_t3_k1 = AES_r1_t3_t3_s4_out;
    always @ (  posedge AES_r1_t3_t3_s4_clk)
    begin
        case ( AES_r1_t3_t3_s4_in ) 
        8'h00:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc6;
        end
        8'h01:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf8;
        end
        8'h02:
        begin
            AES_r1_t3_t3_s4_out <= 8'hee;
        end
        8'h03:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf6;
        end
        8'h04:
        begin
            AES_r1_t3_t3_s4_out <= 8'hff;
        end
        8'h05:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd6;
        end
        8'h06:
        begin
            AES_r1_t3_t3_s4_out <= 8'hde;
        end
        8'h07:
        begin
            AES_r1_t3_t3_s4_out <= 8'h91;
        end
        8'h08:
        begin
            AES_r1_t3_t3_s4_out <= 8'h60;
        end
        8'h09:
        begin
            AES_r1_t3_t3_s4_out <= 8'h02;
        end
        8'h0a:
        begin
            AES_r1_t3_t3_s4_out <= 8'hce;
        end
        8'h0b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h56;
        end
        8'h0c:
        begin
            AES_r1_t3_t3_s4_out <= 8'he7;
        end
        8'h0d:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb5;
        end
        8'h0e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4d;
        end
        8'h0f:
        begin
            AES_r1_t3_t3_s4_out <= 8'hec;
        end
        8'h10:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8f;
        end
        8'h11:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1f;
        end
        8'h12:
        begin
            AES_r1_t3_t3_s4_out <= 8'h89;
        end
        8'h13:
        begin
            AES_r1_t3_t3_s4_out <= 8'hfa;
        end
        8'h14:
        begin
            AES_r1_t3_t3_s4_out <= 8'hef;
        end
        8'h15:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb2;
        end
        8'h16:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8e;
        end
        8'h17:
        begin
            AES_r1_t3_t3_s4_out <= 8'hfb;
        end
        8'h18:
        begin
            AES_r1_t3_t3_s4_out <= 8'h41;
        end
        8'h19:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb3;
        end
        8'h1a:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5f;
        end
        8'h1b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h45;
        end
        8'h1c:
        begin
            AES_r1_t3_t3_s4_out <= 8'h23;
        end
        8'h1d:
        begin
            AES_r1_t3_t3_s4_out <= 8'h53;
        end
        8'h1e:
        begin
            AES_r1_t3_t3_s4_out <= 8'he4;
        end
        8'h1f:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9b;
        end
        8'h20:
        begin
            AES_r1_t3_t3_s4_out <= 8'h75;
        end
        8'h21:
        begin
            AES_r1_t3_t3_s4_out <= 8'he1;
        end
        8'h22:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3d;
        end
        8'h23:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4c;
        end
        8'h24:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6c;
        end
        8'h25:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7e;
        end
        8'h26:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf5;
        end
        8'h27:
        begin
            AES_r1_t3_t3_s4_out <= 8'h83;
        end
        8'h28:
        begin
            AES_r1_t3_t3_s4_out <= 8'h68;
        end
        8'h29:
        begin
            AES_r1_t3_t3_s4_out <= 8'h51;
        end
        8'h2a:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd1;
        end
        8'h2b:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf9;
        end
        8'h2c:
        begin
            AES_r1_t3_t3_s4_out <= 8'he2;
        end
        8'h2d:
        begin
            AES_r1_t3_t3_s4_out <= 8'hab;
        end
        8'h2e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h62;
        end
        8'h2f:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2a;
        end
        8'h30:
        begin
            AES_r1_t3_t3_s4_out <= 8'h08;
        end
        8'h31:
        begin
            AES_r1_t3_t3_s4_out <= 8'h95;
        end
        8'h32:
        begin
            AES_r1_t3_t3_s4_out <= 8'h46;
        end
        8'h33:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9d;
        end
        8'h34:
        begin
            AES_r1_t3_t3_s4_out <= 8'h30;
        end
        8'h35:
        begin
            AES_r1_t3_t3_s4_out <= 8'h37;
        end
        8'h36:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0a;
        end
        8'h37:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2f;
        end
        8'h38:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0e;
        end
        8'h39:
        begin
            AES_r1_t3_t3_s4_out <= 8'h24;
        end
        8'h3a:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1b;
        end
        8'h3b:
        begin
            AES_r1_t3_t3_s4_out <= 8'hdf;
        end
        8'h3c:
        begin
            AES_r1_t3_t3_s4_out <= 8'hcd;
        end
        8'h3d:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4e;
        end
        8'h3e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7f;
        end
        8'h3f:
        begin
            AES_r1_t3_t3_s4_out <= 8'hea;
        end
        8'h40:
        begin
            AES_r1_t3_t3_s4_out <= 8'h12;
        end
        8'h41:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1d;
        end
        8'h42:
        begin
            AES_r1_t3_t3_s4_out <= 8'h58;
        end
        8'h43:
        begin
            AES_r1_t3_t3_s4_out <= 8'h34;
        end
        8'h44:
        begin
            AES_r1_t3_t3_s4_out <= 8'h36;
        end
        8'h45:
        begin
            AES_r1_t3_t3_s4_out <= 8'hdc;
        end
        8'h46:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb4;
        end
        8'h47:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5b;
        end
        8'h48:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha4;
        end
        8'h49:
        begin
            AES_r1_t3_t3_s4_out <= 8'h76;
        end
        8'h4a:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb7;
        end
        8'h4b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7d;
        end
        8'h4c:
        begin
            AES_r1_t3_t3_s4_out <= 8'h52;
        end
        8'h4d:
        begin
            AES_r1_t3_t3_s4_out <= 8'hdd;
        end
        8'h4e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5e;
        end
        8'h4f:
        begin
            AES_r1_t3_t3_s4_out <= 8'h13;
        end
        8'h50:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha6;
        end
        8'h51:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb9;
        end
        8'h52:
        begin
            AES_r1_t3_t3_s4_out <= 8'h00;
        end
        8'h53:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc1;
        end
        8'h54:
        begin
            AES_r1_t3_t3_s4_out <= 8'h40;
        end
        8'h55:
        begin
            AES_r1_t3_t3_s4_out <= 8'he3;
        end
        8'h56:
        begin
            AES_r1_t3_t3_s4_out <= 8'h79;
        end
        8'h57:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb6;
        end
        8'h58:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd4;
        end
        8'h59:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8d;
        end
        8'h5a:
        begin
            AES_r1_t3_t3_s4_out <= 8'h67;
        end
        8'h5b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h72;
        end
        8'h5c:
        begin
            AES_r1_t3_t3_s4_out <= 8'h94;
        end
        8'h5d:
        begin
            AES_r1_t3_t3_s4_out <= 8'h98;
        end
        8'h5e:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb0;
        end
        8'h5f:
        begin
            AES_r1_t3_t3_s4_out <= 8'h85;
        end
        8'h60:
        begin
            AES_r1_t3_t3_s4_out <= 8'hbb;
        end
        8'h61:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc5;
        end
        8'h62:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4f;
        end
        8'h63:
        begin
            AES_r1_t3_t3_s4_out <= 8'hed;
        end
        8'h64:
        begin
            AES_r1_t3_t3_s4_out <= 8'h86;
        end
        8'h65:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9a;
        end
        8'h66:
        begin
            AES_r1_t3_t3_s4_out <= 8'h66;
        end
        8'h67:
        begin
            AES_r1_t3_t3_s4_out <= 8'h11;
        end
        8'h68:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8a;
        end
        8'h69:
        begin
            AES_r1_t3_t3_s4_out <= 8'he9;
        end
        8'h6a:
        begin
            AES_r1_t3_t3_s4_out <= 8'h04;
        end
        8'h6b:
        begin
            AES_r1_t3_t3_s4_out <= 8'hfe;
        end
        8'h6c:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha0;
        end
        8'h6d:
        begin
            AES_r1_t3_t3_s4_out <= 8'h78;
        end
        8'h6e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h25;
        end
        8'h6f:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4b;
        end
        8'h70:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha2;
        end
        8'h71:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5d;
        end
        8'h72:
        begin
            AES_r1_t3_t3_s4_out <= 8'h80;
        end
        8'h73:
        begin
            AES_r1_t3_t3_s4_out <= 8'h05;
        end
        8'h74:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3f;
        end
        8'h75:
        begin
            AES_r1_t3_t3_s4_out <= 8'h21;
        end
        8'h76:
        begin
            AES_r1_t3_t3_s4_out <= 8'h70;
        end
        8'h77:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf1;
        end
        8'h78:
        begin
            AES_r1_t3_t3_s4_out <= 8'h63;
        end
        8'h79:
        begin
            AES_r1_t3_t3_s4_out <= 8'h77;
        end
        8'h7a:
        begin
            AES_r1_t3_t3_s4_out <= 8'haf;
        end
        8'h7b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h42;
        end
        8'h7c:
        begin
            AES_r1_t3_t3_s4_out <= 8'h20;
        end
        8'h7d:
        begin
            AES_r1_t3_t3_s4_out <= 8'he5;
        end
        8'h7e:
        begin
            AES_r1_t3_t3_s4_out <= 8'hfd;
        end
        8'h7f:
        begin
            AES_r1_t3_t3_s4_out <= 8'hbf;
        end
        8'h80:
        begin
            AES_r1_t3_t3_s4_out <= 8'h81;
        end
        8'h81:
        begin
            AES_r1_t3_t3_s4_out <= 8'h18;
        end
        8'h82:
        begin
            AES_r1_t3_t3_s4_out <= 8'h26;
        end
        8'h83:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc3;
        end
        8'h84:
        begin
            AES_r1_t3_t3_s4_out <= 8'hbe;
        end
        8'h85:
        begin
            AES_r1_t3_t3_s4_out <= 8'h35;
        end
        8'h86:
        begin
            AES_r1_t3_t3_s4_out <= 8'h88;
        end
        8'h87:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2e;
        end
        8'h88:
        begin
            AES_r1_t3_t3_s4_out <= 8'h93;
        end
        8'h89:
        begin
            AES_r1_t3_t3_s4_out <= 8'h55;
        end
        8'h8a:
        begin
            AES_r1_t3_t3_s4_out <= 8'hfc;
        end
        8'h8b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7a;
        end
        8'h8c:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc8;
        end
        8'h8d:
        begin
            AES_r1_t3_t3_s4_out <= 8'hba;
        end
        8'h8e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h32;
        end
        8'h8f:
        begin
            AES_r1_t3_t3_s4_out <= 8'he6;
        end
        8'h90:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc0;
        end
        8'h91:
        begin
            AES_r1_t3_t3_s4_out <= 8'h19;
        end
        8'h92:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9e;
        end
        8'h93:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha3;
        end
        8'h94:
        begin
            AES_r1_t3_t3_s4_out <= 8'h44;
        end
        8'h95:
        begin
            AES_r1_t3_t3_s4_out <= 8'h54;
        end
        8'h96:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3b;
        end
        8'h97:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0b;
        end
        8'h98:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8c;
        end
        8'h99:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc7;
        end
        8'h9a:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6b;
        end
        8'h9b:
        begin
            AES_r1_t3_t3_s4_out <= 8'h28;
        end
        8'h9c:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha7;
        end
        8'h9d:
        begin
            AES_r1_t3_t3_s4_out <= 8'hbc;
        end
        8'h9e:
        begin
            AES_r1_t3_t3_s4_out <= 8'h16;
        end
        8'h9f:
        begin
            AES_r1_t3_t3_s4_out <= 8'had;
        end
        8'ha0:
        begin
            AES_r1_t3_t3_s4_out <= 8'hdb;
        end
        8'ha1:
        begin
            AES_r1_t3_t3_s4_out <= 8'h64;
        end
        8'ha2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h74;
        end
        8'ha3:
        begin
            AES_r1_t3_t3_s4_out <= 8'h14;
        end
        8'ha4:
        begin
            AES_r1_t3_t3_s4_out <= 8'h92;
        end
        8'ha5:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0c;
        end
        8'ha6:
        begin
            AES_r1_t3_t3_s4_out <= 8'h48;
        end
        8'ha7:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb8;
        end
        8'ha8:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9f;
        end
        8'ha9:
        begin
            AES_r1_t3_t3_s4_out <= 8'hbd;
        end
        8'haa:
        begin
            AES_r1_t3_t3_s4_out <= 8'h43;
        end
        8'hab:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc4;
        end
        8'hac:
        begin
            AES_r1_t3_t3_s4_out <= 8'h39;
        end
        8'had:
        begin
            AES_r1_t3_t3_s4_out <= 8'h31;
        end
        8'hae:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd3;
        end
        8'haf:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf2;
        end
        8'hb0:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd5;
        end
        8'hb1:
        begin
            AES_r1_t3_t3_s4_out <= 8'h8b;
        end
        8'hb2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6e;
        end
        8'hb3:
        begin
            AES_r1_t3_t3_s4_out <= 8'hda;
        end
        8'hb4:
        begin
            AES_r1_t3_t3_s4_out <= 8'h01;
        end
        8'hb5:
        begin
            AES_r1_t3_t3_s4_out <= 8'hb1;
        end
        8'hb6:
        begin
            AES_r1_t3_t3_s4_out <= 8'h9c;
        end
        8'hb7:
        begin
            AES_r1_t3_t3_s4_out <= 8'h49;
        end
        8'hb8:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd8;
        end
        8'hb9:
        begin
            AES_r1_t3_t3_s4_out <= 8'hac;
        end
        8'hba:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf3;
        end
        8'hbb:
        begin
            AES_r1_t3_t3_s4_out <= 8'hcf;
        end
        8'hbc:
        begin
            AES_r1_t3_t3_s4_out <= 8'hca;
        end
        8'hbd:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf4;
        end
        8'hbe:
        begin
            AES_r1_t3_t3_s4_out <= 8'h47;
        end
        8'hbf:
        begin
            AES_r1_t3_t3_s4_out <= 8'h10;
        end
        8'hc0:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6f;
        end
        8'hc1:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf0;
        end
        8'hc2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h4a;
        end
        8'hc3:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5c;
        end
        8'hc4:
        begin
            AES_r1_t3_t3_s4_out <= 8'h38;
        end
        8'hc5:
        begin
            AES_r1_t3_t3_s4_out <= 8'h57;
        end
        8'hc6:
        begin
            AES_r1_t3_t3_s4_out <= 8'h73;
        end
        8'hc7:
        begin
            AES_r1_t3_t3_s4_out <= 8'h97;
        end
        8'hc8:
        begin
            AES_r1_t3_t3_s4_out <= 8'hcb;
        end
        8'hc9:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha1;
        end
        8'hca:
        begin
            AES_r1_t3_t3_s4_out <= 8'he8;
        end
        8'hcb:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3e;
        end
        8'hcc:
        begin
            AES_r1_t3_t3_s4_out <= 8'h96;
        end
        8'hcd:
        begin
            AES_r1_t3_t3_s4_out <= 8'h61;
        end
        8'hce:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0d;
        end
        8'hcf:
        begin
            AES_r1_t3_t3_s4_out <= 8'h0f;
        end
        8'hd0:
        begin
            AES_r1_t3_t3_s4_out <= 8'he0;
        end
        8'hd1:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7c;
        end
        8'hd2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h71;
        end
        8'hd3:
        begin
            AES_r1_t3_t3_s4_out <= 8'hcc;
        end
        8'hd4:
        begin
            AES_r1_t3_t3_s4_out <= 8'h90;
        end
        8'hd5:
        begin
            AES_r1_t3_t3_s4_out <= 8'h06;
        end
        8'hd6:
        begin
            AES_r1_t3_t3_s4_out <= 8'hf7;
        end
        8'hd7:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1c;
        end
        8'hd8:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc2;
        end
        8'hd9:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6a;
        end
        8'hda:
        begin
            AES_r1_t3_t3_s4_out <= 8'hae;
        end
        8'hdb:
        begin
            AES_r1_t3_t3_s4_out <= 8'h69;
        end
        8'hdc:
        begin
            AES_r1_t3_t3_s4_out <= 8'h17;
        end
        8'hdd:
        begin
            AES_r1_t3_t3_s4_out <= 8'h99;
        end
        8'hde:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3a;
        end
        8'hdf:
        begin
            AES_r1_t3_t3_s4_out <= 8'h27;
        end
        8'he0:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd9;
        end
        8'he1:
        begin
            AES_r1_t3_t3_s4_out <= 8'heb;
        end
        8'he2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2b;
        end
        8'he3:
        begin
            AES_r1_t3_t3_s4_out <= 8'h22;
        end
        8'he4:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd2;
        end
        8'he5:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha9;
        end
        8'he6:
        begin
            AES_r1_t3_t3_s4_out <= 8'h07;
        end
        8'he7:
        begin
            AES_r1_t3_t3_s4_out <= 8'h33;
        end
        8'he8:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2d;
        end
        8'he9:
        begin
            AES_r1_t3_t3_s4_out <= 8'h3c;
        end
        8'hea:
        begin
            AES_r1_t3_t3_s4_out <= 8'h15;
        end
        8'heb:
        begin
            AES_r1_t3_t3_s4_out <= 8'hc9;
        end
        8'hec:
        begin
            AES_r1_t3_t3_s4_out <= 8'h87;
        end
        8'hed:
        begin
            AES_r1_t3_t3_s4_out <= 8'haa;
        end
        8'hee:
        begin
            AES_r1_t3_t3_s4_out <= 8'h50;
        end
        8'hef:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha5;
        end
        8'hf0:
        begin
            AES_r1_t3_t3_s4_out <= 8'h03;
        end
        8'hf1:
        begin
            AES_r1_t3_t3_s4_out <= 8'h59;
        end
        8'hf2:
        begin
            AES_r1_t3_t3_s4_out <= 8'h09;
        end
        8'hf3:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1a;
        end
        8'hf4:
        begin
            AES_r1_t3_t3_s4_out <= 8'h65;
        end
        8'hf5:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd7;
        end
        8'hf6:
        begin
            AES_r1_t3_t3_s4_out <= 8'h84;
        end
        8'hf7:
        begin
            AES_r1_t3_t3_s4_out <= 8'hd0;
        end
        8'hf8:
        begin
            AES_r1_t3_t3_s4_out <= 8'h82;
        end
        8'hf9:
        begin
            AES_r1_t3_t3_s4_out <= 8'h29;
        end
        8'hfa:
        begin
            AES_r1_t3_t3_s4_out <= 8'h5a;
        end
        8'hfb:
        begin
            AES_r1_t3_t3_s4_out <= 8'h1e;
        end
        8'hfc:
        begin
            AES_r1_t3_t3_s4_out <= 8'h7b;
        end
        8'hfd:
        begin
            AES_r1_t3_t3_s4_out <= 8'ha8;
        end
        8'hfe:
        begin
            AES_r1_t3_t3_s4_out <= 8'h6d;
        end
        8'hff:
        begin
            AES_r1_t3_t3_s4_out <= 8'h2c;
        end
        endcase
    end
    assign AES_r1_t3_t3_out = { AES_r1_t3_t3_k0, AES_r1_t3_t3_k0, ( AES_r1_t3_t3_k0 ^ AES_r1_t3_t3_k1 ), AES_r1_t3_t3_k1 };
    assign AES_r1_z0 = ( ( ( ( AES_r1_p00 ^ AES_r1_p11 ) ^ AES_r1_p22 ) ^ AES_r1_p33 ) ^ AES_r1_k0 );
    assign AES_r1_z1 = ( ( ( ( AES_r1_p03 ^ AES_r1_p10 ) ^ AES_r1_p21 ) ^ AES_r1_p32 ) ^ AES_r1_k1 );
    assign AES_r1_z2 = ( ( ( ( AES_r1_p02 ^ AES_r1_p13 ) ^ AES_r1_p20 ) ^ AES_r1_p31 ) ^ AES_r1_k2 );
    assign AES_r1_z3 = ( ( ( ( AES_r1_p01 ^ AES_r1_p12 ) ^ AES_r1_p23 ) ^ AES_r1_p30 ) ^ AES_r1_k3 );
    always @ (  posedge AES_r1_clk)
    begin
        AES_r1_state_out <= { AES_r1_z0, AES_r1_z1, AES_r1_z2, AES_r1_z3 };
    end
endmodule 


