module ram_2x3 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [2:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [2:0] W0_data;
	reg [2:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 3'bxxx);
endmodule
module ram_2x8 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [7:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [7:0] W0_data;
	reg [7:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 8'bxxxxxxxx);
endmodule
module ram_data_2x64 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [63:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [63:0] W0_data;
	reg [63:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [63:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module ram_2x1 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input W0_data;
	reg Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 1'bx);
endmodule
module ram_param_2x2 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [1:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [1:0] W0_data;
	reg [1:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 2'bxx);
endmodule
module ram_size_2x4 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [3:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [3:0] W0_data;
	reg [3:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 4'bxxxx);
endmodule
module ram_address_2x32 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [31:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [31:0] W0_data;
	reg [31:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module Queue_37 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_data,
	io_enq_bits_strb,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_data,
	io_deq_bits_strb,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [63:0] io_enq_bits_data;
	input [7:0] io_enq_bits_strb;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [63:0] io_deq_bits_data;
	output wire [7:0] io_deq_bits_strb;
	output wire io_deq_bits_last;
	reg ram_last;
	reg [7:0] ram_strb;
	reg [63:0] ram_data;
	reg full;
	wire _io_deq_valid_output = io_enq_valid | full;
	wire do_enq = (~(~full & io_deq_ready) & ~full) & io_enq_valid;
	always @(posedge clock) begin
		if (do_enq) begin
			ram_last <= io_enq_bits_last;
			ram_strb <= io_enq_bits_strb;
			ram_data <= io_enq_bits_data;
		end
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == ((full & io_deq_ready) & _io_deq_valid_output)))
			full <= do_enq;
	end
	wire [31:0] _RANDOM [0:2];
	assign io_enq_ready = ~full;
	assign io_deq_valid = _io_deq_valid_output;
	assign io_deq_bits_data = (full ? ram_data : io_enq_bits_data);
	assign io_deq_bits_strb = (full ? ram_strb : io_enq_bits_strb);
	assign io_deq_bits_last = (full ? ram_last : io_enq_bits_last);
endmodule
module IntXbar_1 (
	auto_int_in_3_0,
	auto_int_in_2_0,
	auto_int_in_1_0,
	auto_int_in_1_1,
	auto_int_in_0_0,
	auto_int_out_0,
	auto_int_out_1,
	auto_int_out_2,
	auto_int_out_3,
	auto_int_out_4
);
	input auto_int_in_3_0;
	input auto_int_in_2_0;
	input auto_int_in_1_0;
	input auto_int_in_1_1;
	input auto_int_in_0_0;
	output wire auto_int_out_0;
	output wire auto_int_out_1;
	output wire auto_int_out_2;
	output wire auto_int_out_3;
	output wire auto_int_out_4;
	assign auto_int_out_0 = auto_int_in_0_0;
	assign auto_int_out_1 = auto_int_in_1_0;
	assign auto_int_out_2 = auto_int_in_1_1;
	assign auto_int_out_3 = auto_int_in_2_0;
	assign auto_int_out_4 = auto_int_in_3_0;
endmodule
module TLMonitor_40 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [3:0] io_in_a_bits_size;
	input [5:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [7:0] io_in_a_bits_mask;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [5:0] io_in_d_bits_source;
	input [2:0] io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] _plusarg_reader_1_out;
	wire [31:0] _plusarg_reader_out;
	wire [26:0] _GEN = {23'h000000, io_in_a_bits_size};
	wire _a_first_T_1 = io_in_a_ready & io_in_a_valid;
	reg [8:0] a_first_counter;
	reg [2:0] opcode;
	reg [3:0] size;
	reg [5:0] source;
	reg [31:0] address;
	reg [8:0] d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [5:0] source_1;
	reg [2:0] sink;
	reg denied;
	reg [63:0] inflight;
	reg [255:0] inflight_opcodes;
	reg [511:0] inflight_sizes;
	reg [8:0] a_first_counter_1;
	wire a_first_1 = a_first_counter_1 == 9'h000;
	reg [8:0] d_first_counter_1;
	wire d_first_1 = d_first_counter_1 == 9'h000;
	wire [63:0] _GEN_0 = {58'h000000000000000, io_in_a_bits_source};
	wire _GEN_1 = _a_first_T_1 & a_first_1;
	wire d_release_ack = io_in_d_bits_opcode == 3'h6;
	wire [63:0] _GEN_2 = {58'h000000000000000, io_in_d_bits_source};
	reg [31:0] watchdog;
	reg [63:0] inflight_1;
	reg [511:0] inflight_sizes_1;
	reg [8:0] d_first_counter_2;
	wire d_first_2 = d_first_counter_2 == 9'h000;
	reg [31:0] watchdog_1;
	wire [23:0] _GEN_3 = 24'h951240;
	wire [23:0] _GEN_4 = 24'h911240;
	wire source_ok = ((((((((((((((~(|io_in_a_bits_source[5:2]) | (io_in_a_bits_source[5:2] == 4'h1)) | (io_in_a_bits_source[5:2] == 4'h2)) | (io_in_a_bits_source[5:2] == 4'h3)) | (io_in_a_bits_source[5:2] == 4'h4)) | (io_in_a_bits_source[5:2] == 4'h5)) | (io_in_a_bits_source[5:2] == 4'h6)) | (io_in_a_bits_source[5:2] == 4'h7)) | (io_in_a_bits_source[5:2] == 4'h8)) | (io_in_a_bits_source[5:2] == 4'h9)) | (io_in_a_bits_source[5:2] == 4'ha)) | (io_in_a_bits_source[5:2] == 4'hb)) | (io_in_a_bits_source[5:2] == 4'hc)) | (io_in_a_bits_source[5:2] == 4'hd)) | (io_in_a_bits_source[5:2] == 4'he)) | &io_in_a_bits_source[5:2];
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << _GEN;
	wire [11:0] _GEN_5 = io_in_a_bits_address[11:0] & ~_is_aligned_mask_T_1[11:0];
	wire _mask_T = io_in_a_bits_size > 4'h2;
	wire mask_size = io_in_a_bits_size[1:0] == 2'h2;
	wire mask_acc = _mask_T | (mask_size & ~io_in_a_bits_address[2]);
	wire mask_acc_1 = _mask_T | (mask_size & io_in_a_bits_address[2]);
	wire mask_size_1 = io_in_a_bits_size[1:0] == 2'h1;
	wire mask_eq_2 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1];
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1];
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1];
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = io_in_a_bits_address[2] & io_in_a_bits_address[1];
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [7:0] mask = {mask_acc_5 | (mask_eq_5 & io_in_a_bits_address[0]), mask_acc_5 | (mask_eq_5 & ~io_in_a_bits_address[0]), mask_acc_4 | (mask_eq_4 & io_in_a_bits_address[0]), mask_acc_4 | (mask_eq_4 & ~io_in_a_bits_address[0]), mask_acc_3 | (mask_eq_3 & io_in_a_bits_address[0]), mask_acc_3 | (mask_eq_3 & ~io_in_a_bits_address[0]), mask_acc_2 | (mask_eq_2 & io_in_a_bits_address[0]), mask_acc_2 | (mask_eq_2 & ~io_in_a_bits_address[0])};
	wire _GEN_6 = io_in_a_bits_size < 4'hd;
	wire _GEN_7 = _GEN_6 & (((((((((((((((~(|io_in_a_bits_source[5:2]) | (io_in_a_bits_source[5:2] == 4'h1)) | (io_in_a_bits_source[5:2] == 4'h2)) | (io_in_a_bits_source[5:2] == 4'h3)) | (io_in_a_bits_source[5:2] == 4'h4)) | (io_in_a_bits_source[5:2] == 4'h5)) | (io_in_a_bits_source[5:2] == 4'h6)) | (io_in_a_bits_source[5:2] == 4'h7)) | (io_in_a_bits_source[5:2] == 4'h8)) | (io_in_a_bits_source[5:2] == 4'h9)) | (io_in_a_bits_source[5:2] == 4'ha)) | (io_in_a_bits_source[5:2] == 4'hb)) | (io_in_a_bits_source[5:2] == 4'hc)) | (io_in_a_bits_source[5:2] == 4'hd)) | (io_in_a_bits_source[5:2] == 4'he)) | &io_in_a_bits_source[5:2]);
	wire _GEN_8 = {io_in_a_bits_address[31:28], io_in_a_bits_address[27:16] ^ 12'h800} == 16'h0000;
	wire _GEN_9 = io_in_a_bits_address[31:28] == 4'h8;
	wire _GEN_10 = _GEN_8 | _GEN_9;
	wire _GEN_11 = (_GEN_7 & (io_in_a_bits_size == 4'h6)) & _GEN_10;
	wire _GEN_12 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h6)) & ~reset;
	wire _GEN_13 = io_in_a_bits_mask != 8'hff;
	wire _GEN_14 = (io_in_a_valid & &io_in_a_bits_opcode) & ~reset;
	wire _GEN_15 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h4)) & ~reset;
	wire _GEN_16 = {io_in_a_bits_address[31:14], ~io_in_a_bits_address[13:12]} == 20'h00000;
	wire _GEN_17 = _GEN_6 & _GEN_16;
	wire _GEN_18 = io_in_a_bits_size < 4'h7;
	wire _GEN_19 = io_in_a_bits_address[31:13] == 19'h00000;
	wire _GEN_20 = {io_in_a_bits_address[31:21], io_in_a_bits_address[20:17] ^ 4'h8, io_in_a_bits_address[15:12]} == 19'h00000;
	wire _GEN_21 = {io_in_a_bits_address[31:26], io_in_a_bits_address[25:16] ^ 10'h200} == 16'h0000;
	wire _GEN_22 = {io_in_a_bits_address[31:26], io_in_a_bits_address[25:12] ^ 14'h2010} == 20'h00000;
	wire _GEN_23 = {io_in_a_bits_address[31:28], ~io_in_a_bits_address[27:26]} == 6'h00;
	wire _GEN_24 = {io_in_a_bits_address[31:29], io_in_a_bits_address[28:12] ^ 17'h10020} == 20'h00000;
	wire _GEN_25 = io_in_a_bits_mask != mask;
	wire _GEN_26 = _GEN_7 & (_GEN_17 | (_GEN_18 & (((((((_GEN_19 | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9)));
	wire _GEN_27 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h0)) & ~reset;
	wire _GEN_28 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h1)) & ~reset;
	wire _GEN_29 = (_GEN_7 & (io_in_a_bits_size < 4'h4)) & ((((((((_GEN_19 | _GEN_16) | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9);
	wire _GEN_30 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h2)) & ~reset;
	wire _GEN_31 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h3)) & ~reset;
	wire _GEN_32 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h5)) & ~reset;
	wire source_ok_1 = (((((((((((((((io_in_d_bits_source[5:2] == 4'h0) | (io_in_d_bits_source[5:2] == 4'h1)) | (io_in_d_bits_source[5:2] == 4'h2)) | (io_in_d_bits_source[5:2] == 4'h3)) | (io_in_d_bits_source[5:2] == 4'h4)) | (io_in_d_bits_source[5:2] == 4'h5)) | (io_in_d_bits_source[5:2] == 4'h6)) | (io_in_d_bits_source[5:2] == 4'h7)) | (io_in_d_bits_source[5:2] == 4'h8)) | (io_in_d_bits_source[5:2] == 4'h9)) | (io_in_d_bits_source[5:2] == 4'ha)) | (io_in_d_bits_source[5:2] == 4'hb)) | (io_in_d_bits_source[5:2] == 4'hc)) | (io_in_d_bits_source[5:2] == 4'hd)) | (io_in_d_bits_source[5:2] == 4'he)) | &io_in_d_bits_source[5:2];
	wire _GEN_33 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h6)) & ~reset;
	wire _GEN_34 = io_in_d_bits_size < 4'h3;
	wire _GEN_35 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h4)) & ~reset;
	wire _GEN_36 = io_in_d_bits_param == 2'h2;
	wire _GEN_37 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h5)) & ~reset;
	wire _GEN_38 = ~io_in_d_bits_denied | io_in_d_bits_corrupt;
	wire _GEN_39 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h0)) & ~reset;
	wire _GEN_40 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h1)) & ~reset;
	wire _GEN_41 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h2)) & ~reset;
	wire _GEN_42 = (io_in_a_valid & |a_first_counter) & ~reset;
	wire _GEN_43 = (io_in_d_valid & |d_first_counter) & ~reset;
	wire [255:0] _a_opcode_lookup_T_1 = inflight_opcodes >> {248'h00000000000000000000000000000000000000000000000000000000000000, io_in_d_bits_source, 2'h0};
	wire [511:0] _GEN_44 = {503'h0, io_in_d_bits_source, 3'h0};
	wire _same_cycle_resp_T_1 = io_in_a_valid & a_first_1;
	wire [63:0] a_set_wo_ready = (_same_cycle_resp_T_1 ? 64'h0000000000000001 << _GEN_0 : 64'h0000000000000000);
	wire _GEN_45 = io_in_d_valid & d_first_1;
	wire _GEN_46 = _GEN_45 & ~d_release_ack;
	wire same_cycle_resp = _same_cycle_resp_T_1 & (io_in_a_bits_source == io_in_d_bits_source);
	wire _GEN_47 = (_GEN_46 & same_cycle_resp) & ~reset;
	wire _GEN_48 = (_GEN_46 & ~same_cycle_resp) & ~reset;
	wire [7:0] _GEN_49 = {4'h0, io_in_d_bits_size};
	wire _GEN_50 = ((io_in_d_valid & d_first_2) & d_release_ack) & ~reset;
	wire [63:0] _GEN_51 = inflight >> _GEN_0;
	wire [63:0] _GEN_52 = inflight >> _GEN_2;
	wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _GEN_44;
	wire [63:0] _GEN_53 = inflight_1 >> _GEN_2;
	wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _GEN_44;
	always @(posedge clock) begin
		if (_GEN_12 & ~_GEN_11) begin
			$error("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12) begin
			$error("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & ~source_ok) begin
			$error("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & ~_mask_T) begin
			$error("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & _GEN_13) begin
			$error("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~_GEN_11) begin
			$error("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14) begin
			$error("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~source_ok) begin
			$error("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~_mask_T) begin
			$error("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14) begin
			$error("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & _GEN_13) begin
			$error("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~_GEN_7) begin
			$error("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~(_GEN_17 | (_GEN_18 & ((((((((_GEN_19 | ({io_in_a_bits_address[31:17], ~io_in_a_bits_address[16]} == 16'h0000)) | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9)))) begin
			$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Get carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Get address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Get contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & ~_GEN_26) begin
			$error("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & ~source_ok) begin
			$error("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel PutFull address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & _GEN_25) begin
			$error("Assertion failed: 'A' channel PutFull contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & ~_GEN_26) begin
			$error("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & ~source_ok) begin
			$error("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & |(io_in_a_bits_mask & ~mask)) begin
			$error("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & ~_GEN_29) begin
			$error("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & ~_GEN_29) begin
			$error("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Logical carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Logical address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Logical contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & ~(_GEN_7 & (_GEN_17 | (_GEN_18 & _GEN_10)))) begin
			$error("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Hint carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Hint address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Hint contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if ((io_in_d_valid & ~reset) & &io_in_d_bits_opcode) begin
			$error("Assertion failed: 'D' channel has invalid opcode (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & _GEN_34) begin
			$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & io_in_d_bits_denied) begin
			$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel Grant carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & _GEN_34) begin
			$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & &io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & _GEN_36) begin
			$error("Assertion failed: 'D' channel Grant carries toN param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel Grant is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & _GEN_34) begin
			$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & &io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & _GEN_36) begin
			$error("Assertion failed: 'D' channel GrantData carries toN param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & ~_GEN_38) begin
			$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & ~_GEN_38) begin
			$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel HintAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_opcode != opcode)) begin
			$error("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_size != size)) begin
			$error("Assertion failed: 'A' channel size changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_source != source)) begin
			$error("Assertion failed: 'A' channel source changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_address != address)) begin
			$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_opcode != opcode_1)) begin
			$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_param != param_1)) begin
			$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_size != size_1)) begin
			$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_source != source_1)) begin
			$error("Assertion failed: 'D' channel source changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_sink != sink)) begin
			$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_denied != denied)) begin
			$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if ((_GEN_1 & ~reset) & _GEN_51[0]) begin
			$error("Assertion failed: 'A' channel re-used a source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if ((_GEN_46 & ~reset) & ~(_GEN_52[0] | same_cycle_resp)) begin
			$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_47 & ~((io_in_d_bits_opcode == _GEN_4[io_in_a_bits_opcode * 3+:3]) | (io_in_d_bits_opcode == _GEN_3[io_in_a_bits_opcode * 3+:3]))) begin
			$error("Assertion failed: 'D' channel contains improper opcode response (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_47 & (io_in_a_bits_size != io_in_d_bits_size)) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_48 & ~((io_in_d_bits_opcode == _GEN_4[_a_opcode_lookup_T_1[3:1] * 3+:3]) | (io_in_d_bits_opcode == _GEN_3[_a_opcode_lookup_T_1[3:1] * 3+:3]))) begin
			$error("Assertion failed: 'D' channel contains improper opcode response (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_48 & (_GEN_49 != {1'h0, _a_size_lookup_T_1[7:1]})) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if ((((((_GEN_45 & a_first_1) & io_in_a_valid) & (io_in_a_bits_source == io_in_d_bits_source)) & ~d_release_ack) & ~reset) & ~(~io_in_d_ready | io_in_a_ready)) begin
			$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~((a_set_wo_ready != (_GEN_46 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000)) | (a_set_wo_ready == 64'h0000000000000000))) begin
			$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency > 0 (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~(((inflight == 64'h0000000000000000) | (_plusarg_reader_out == 32'h00000000)) | (watchdog < _plusarg_reader_out))) begin
			$error("Assertion failed: TileLink timeout expired (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_50 & ~_GEN_53[0]) begin
			$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_50 & (_GEN_49 != {1'h0, _c_size_lookup_T_1[7:1]})) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~(((inflight_1 == 64'h0000000000000000) | (_plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < _plusarg_reader_1_out))) begin
			$error("Assertion failed: TileLink timeout expired (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:191:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
	end
	wire [26:0] _a_first_beats1_decode_T_1 = 27'h0000fff << _GEN;
	wire [26:0] _a_first_beats1_decode_T_5 = 27'h0000fff << _GEN;
	wire [26:0] _GEN_54 = {23'h000000, io_in_d_bits_size};
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << _GEN_54;
	wire [26:0] _d_first_beats1_decode_T_5 = 27'h0000fff << _GEN_54;
	wire [26:0] _d_first_beats1_decode_T_9 = 27'h0000fff << _GEN_54;
	wire [526:0] _GEN_55 = {518'h0, io_in_d_bits_source, 3'h0};
	wire [526:0] _d_opcodes_clr_T_5 = 527'hf << {519'h0, io_in_d_bits_source, 2'h0};
	wire [514:0] _a_opcodes_set_T_1 = {511'h0, (_GEN_1 ? {io_in_a_bits_opcode, 1'h1} : 4'h0)} << {507'h0, io_in_a_bits_source, 2'h0};
	wire [526:0] _d_sizes_clr_T_5 = 527'hff << _GEN_55;
	wire [515:0] _a_sizes_set_T_1 = {511'h0, (_GEN_1 ? {io_in_a_bits_size, 1'h1} : 5'h00)} << {507'h0, io_in_a_bits_source, 3'h0};
	wire [526:0] _d_sizes_clr_T_11 = 527'hff << _GEN_55;
	wire _d_first_T_2 = io_in_d_ready & io_in_d_valid;
	wire _GEN_56 = (_d_first_T_2 & d_first_1) & ~d_release_ack;
	wire _GEN_57 = (_d_first_T_2 & d_first_2) & d_release_ack;
	always @(posedge clock) begin
		if (reset) begin
			a_first_counter <= 9'h000;
			d_first_counter <= 9'h000;
			inflight <= 64'h0000000000000000;
			inflight_opcodes <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			inflight_sizes <= 512'h0;
			a_first_counter_1 <= 9'h000;
			d_first_counter_1 <= 9'h000;
			watchdog <= 32'h00000000;
			inflight_1 <= 64'h0000000000000000;
			inflight_sizes_1 <= 512'h0;
			d_first_counter_2 <= 9'h000;
			watchdog_1 <= 32'h00000000;
		end
		else begin
			if (_a_first_T_1) begin
				if (|a_first_counter)
					a_first_counter <= a_first_counter - 9'h001;
				else
					a_first_counter <= (io_in_a_bits_opcode[2] ? 9'h000 : ~_a_first_beats1_decode_T_1[11:3]);
				if (a_first_1)
					a_first_counter_1 <= (io_in_a_bits_opcode[2] ? 9'h000 : ~_a_first_beats1_decode_T_5[11:3]);
				else
					a_first_counter_1 <= a_first_counter_1 - 9'h001;
			end
			if (_d_first_T_2) begin
				if (|d_first_counter)
					d_first_counter <= d_first_counter - 9'h001;
				else
					d_first_counter <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_1[11:3] : 9'h000);
				if (d_first_1)
					d_first_counter_1 <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_5[11:3] : 9'h000);
				else
					d_first_counter_1 <= d_first_counter_1 - 9'h001;
				if (d_first_2)
					d_first_counter_2 <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_9[11:3] : 9'h000);
				else
					d_first_counter_2 <= d_first_counter_2 - 9'h001;
				watchdog_1 <= 32'h00000000;
			end
			else
				watchdog_1 <= watchdog_1 + 32'h00000001;
			inflight <= (inflight | (_GEN_1 ? 64'h0000000000000001 << _GEN_0 : 64'h0000000000000000)) & ~(_GEN_56 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000);
			inflight_opcodes <= (inflight_opcodes | (_GEN_1 ? _a_opcodes_set_T_1[255:0] : 256'h0000000000000000000000000000000000000000000000000000000000000000)) & ~(_GEN_56 ? _d_opcodes_clr_T_5[255:0] : 256'h0000000000000000000000000000000000000000000000000000000000000000);
			inflight_sizes <= (inflight_sizes | (_GEN_1 ? _a_sizes_set_T_1[511:0] : 512'h0)) & ~(_GEN_56 ? _d_sizes_clr_T_5[511:0] : 512'h0);
			if (_a_first_T_1 | _d_first_T_2)
				watchdog <= 32'h00000000;
			else
				watchdog <= watchdog + 32'h00000001;
			inflight_1 <= inflight_1 & ~(_GEN_57 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000);
			inflight_sizes_1 <= inflight_sizes_1 & ~(_GEN_57 ? _d_sizes_clr_T_11[511:0] : 512'h0);
		end
		if (_a_first_T_1 & ~(|a_first_counter)) begin
			opcode <= io_in_a_bits_opcode;
			size <= io_in_a_bits_size;
			source <= io_in_a_bits_source;
			address <= io_in_a_bits_address;
		end
		if (_d_first_T_2 & ~(|d_first_counter)) begin
			opcode_1 <= io_in_d_bits_opcode;
			param_1 <= io_in_d_bits_param;
			size_1 <= io_in_d_bits_size;
			source_1 <= io_in_d_bits_source;
			sink <= io_in_d_bits_sink;
			denied <= io_in_d_bits_denied;
		end
	end
	wire [31:0] _RANDOM [0:57];
	plusarg_reader #(
		.DEFAULT(0),
		.FORMAT("tilelink_timeout=%d"),
		.WIDTH(32)
	) plusarg_reader(.out(_plusarg_reader_out));
	plusarg_reader #(
		.DEFAULT(0),
		.FORMAT("tilelink_timeout=%d"),
		.WIDTH(32)
	) plusarg_reader_1(.out(_plusarg_reader_1_out));
endmodule
module ram_source_2x6 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input R0_addr;
	input R0_en;
	input R0_clk;
	output wire [5:0] R0_data;
	input W0_addr;
	input W0_en;
	input W0_clk;
	input [5:0] W0_data;
	reg [5:0] Memory [0:1];
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	reg [31:0] _RANDOM_MEM;
	assign R0_data = (R0_en ? Memory[R0_addr] : 6'bxxxxxx);
endmodule
module Queue_52 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_address,
	io_enq_bits_mask,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_address,
	io_deq_bits_mask,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [2:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input [5:0] io_enq_bits_source;
	input [31:0] io_enq_bits_address;
	input [7:0] io_enq_bits_mask;
	input [63:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [2:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire [5:0] io_deq_bits_source;
	output wire [31:0] io_deq_bits_address;
	output wire [7:0] io_deq_bits_mask;
	output wire [63:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	wire do_deq = io_deq_ready & ~empty;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	wire [31:0] _RANDOM [0:0];
	ram_2x3 ram_opcode_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_opcode),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_opcode)
	);
	ram_2x3 ram_param_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_param),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_param)
	);
	ram_size_2x4 ram_size_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_size),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_size)
	);
	ram_source_2x6 ram_source_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_source),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_source)
	);
	ram_address_2x32 ram_address_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_address),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_address)
	);
	ram_2x8 ram_mask_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_mask),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_mask)
	);
	ram_data_2x64 ram_data_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_data)
	);
	ram_2x1 ram_corrupt_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_corrupt),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_corrupt)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module Queue_53 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_opcode,
	io_enq_bits_param,
	io_enq_bits_size,
	io_enq_bits_source,
	io_enq_bits_sink,
	io_enq_bits_denied,
	io_enq_bits_data,
	io_enq_bits_corrupt,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_opcode,
	io_deq_bits_param,
	io_deq_bits_size,
	io_deq_bits_source,
	io_deq_bits_sink,
	io_deq_bits_denied,
	io_deq_bits_data,
	io_deq_bits_corrupt
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [2:0] io_enq_bits_opcode;
	input [1:0] io_enq_bits_param;
	input [3:0] io_enq_bits_size;
	input [5:0] io_enq_bits_source;
	input [2:0] io_enq_bits_sink;
	input io_enq_bits_denied;
	input [63:0] io_enq_bits_data;
	input io_enq_bits_corrupt;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [2:0] io_deq_bits_opcode;
	output wire [1:0] io_deq_bits_param;
	output wire [3:0] io_deq_bits_size;
	output wire [5:0] io_deq_bits_source;
	output wire [2:0] io_deq_bits_sink;
	output wire io_deq_bits_denied;
	output wire [63:0] io_deq_bits_data;
	output wire io_deq_bits_corrupt;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	wire do_deq = io_deq_ready & ~empty;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	wire [31:0] _RANDOM [0:0];
	ram_2x3 ram_opcode_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_opcode),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_opcode)
	);
	ram_param_2x2 ram_param_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_param),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_param)
	);
	ram_size_2x4 ram_size_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_size),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_size)
	);
	ram_source_2x6 ram_source_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_source),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_source)
	);
	ram_2x3 ram_sink_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_sink),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_sink)
	);
	ram_2x1 ram_denied_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_denied),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_denied)
	);
	ram_data_2x64 ram_data_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_data),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_data)
	);
	ram_2x1 ram_corrupt_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_corrupt),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_corrupt)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module TLBuffer_14 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_param,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_sink,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_param,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_a_bits_corrupt,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [3:0] auto_in_a_bits_size;
	input [5:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [7:0] auto_in_a_bits_mask;
	input [63:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [1:0] auto_in_d_bits_param;
	output wire [3:0] auto_in_d_bits_size;
	output wire [5:0] auto_in_d_bits_source;
	output wire [2:0] auto_in_d_bits_sink;
	output wire auto_in_d_bits_denied;
	output wire [63:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [2:0] auto_out_a_bits_param;
	output wire [3:0] auto_out_a_bits_size;
	output wire [5:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_a_bits_corrupt;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [5:0] auto_out_d_bits_source;
	input [2:0] auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire _nodeIn_d_q_io_deq_valid;
	wire [2:0] _nodeIn_d_q_io_deq_bits_opcode;
	wire [1:0] _nodeIn_d_q_io_deq_bits_param;
	wire [3:0] _nodeIn_d_q_io_deq_bits_size;
	wire [5:0] _nodeIn_d_q_io_deq_bits_source;
	wire [2:0] _nodeIn_d_q_io_deq_bits_sink;
	wire _nodeIn_d_q_io_deq_bits_denied;
	wire _nodeIn_d_q_io_deq_bits_corrupt;
	wire _nodeOut_a_q_io_enq_ready;
	TLMonitor_40 monitor(
		.clock(clock),
		.reset(reset),
		.io_in_a_ready(_nodeOut_a_q_io_enq_ready),
		.io_in_a_valid(auto_in_a_valid),
		.io_in_a_bits_opcode(auto_in_a_bits_opcode),
		.io_in_a_bits_size(auto_in_a_bits_size),
		.io_in_a_bits_source(auto_in_a_bits_source),
		.io_in_a_bits_address(auto_in_a_bits_address),
		.io_in_a_bits_mask(auto_in_a_bits_mask),
		.io_in_d_ready(auto_in_d_ready),
		.io_in_d_valid(_nodeIn_d_q_io_deq_valid),
		.io_in_d_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),
		.io_in_d_bits_param(_nodeIn_d_q_io_deq_bits_param),
		.io_in_d_bits_size(_nodeIn_d_q_io_deq_bits_size),
		.io_in_d_bits_source(_nodeIn_d_q_io_deq_bits_source),
		.io_in_d_bits_sink(_nodeIn_d_q_io_deq_bits_sink),
		.io_in_d_bits_denied(_nodeIn_d_q_io_deq_bits_denied),
		.io_in_d_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)
	);
	Queue_52 nodeOut_a_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_nodeOut_a_q_io_enq_ready),
		.io_enq_valid(auto_in_a_valid),
		.io_enq_bits_opcode(auto_in_a_bits_opcode),
		.io_enq_bits_param(3'h0),
		.io_enq_bits_size(auto_in_a_bits_size),
		.io_enq_bits_source(auto_in_a_bits_source),
		.io_enq_bits_address(auto_in_a_bits_address),
		.io_enq_bits_mask(auto_in_a_bits_mask),
		.io_enq_bits_data(auto_in_a_bits_data),
		.io_enq_bits_corrupt(1'h0),
		.io_deq_ready(auto_out_a_ready),
		.io_deq_valid(auto_out_a_valid),
		.io_deq_bits_opcode(auto_out_a_bits_opcode),
		.io_deq_bits_param(auto_out_a_bits_param),
		.io_deq_bits_size(auto_out_a_bits_size),
		.io_deq_bits_source(auto_out_a_bits_source),
		.io_deq_bits_address(auto_out_a_bits_address),
		.io_deq_bits_mask(auto_out_a_bits_mask),
		.io_deq_bits_data(auto_out_a_bits_data),
		.io_deq_bits_corrupt(auto_out_a_bits_corrupt)
	);
	Queue_53 nodeIn_d_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(auto_out_d_ready),
		.io_enq_valid(auto_out_d_valid),
		.io_enq_bits_opcode(auto_out_d_bits_opcode),
		.io_enq_bits_param(auto_out_d_bits_param),
		.io_enq_bits_size(auto_out_d_bits_size),
		.io_enq_bits_source(auto_out_d_bits_source),
		.io_enq_bits_sink(auto_out_d_bits_sink),
		.io_enq_bits_denied(auto_out_d_bits_denied),
		.io_enq_bits_data(auto_out_d_bits_data),
		.io_enq_bits_corrupt(auto_out_d_bits_corrupt),
		.io_deq_ready(auto_in_d_ready),
		.io_deq_valid(_nodeIn_d_q_io_deq_valid),
		.io_deq_bits_opcode(_nodeIn_d_q_io_deq_bits_opcode),
		.io_deq_bits_param(_nodeIn_d_q_io_deq_bits_param),
		.io_deq_bits_size(_nodeIn_d_q_io_deq_bits_size),
		.io_deq_bits_source(_nodeIn_d_q_io_deq_bits_source),
		.io_deq_bits_sink(_nodeIn_d_q_io_deq_bits_sink),
		.io_deq_bits_denied(_nodeIn_d_q_io_deq_bits_denied),
		.io_deq_bits_data(auto_in_d_bits_data),
		.io_deq_bits_corrupt(_nodeIn_d_q_io_deq_bits_corrupt)
	);
	assign auto_in_a_ready = _nodeOut_a_q_io_enq_ready;
	assign auto_in_d_valid = _nodeIn_d_q_io_deq_valid;
	assign auto_in_d_bits_opcode = _nodeIn_d_q_io_deq_bits_opcode;
	assign auto_in_d_bits_param = _nodeIn_d_q_io_deq_bits_param;
	assign auto_in_d_bits_size = _nodeIn_d_q_io_deq_bits_size;
	assign auto_in_d_bits_source = _nodeIn_d_q_io_deq_bits_source;
	assign auto_in_d_bits_sink = _nodeIn_d_q_io_deq_bits_sink;
	assign auto_in_d_bits_denied = _nodeIn_d_q_io_deq_bits_denied;
	assign auto_in_d_bits_corrupt = _nodeIn_d_q_io_deq_bits_corrupt;
endmodule
module TLMonitor_41 (
	clock,
	reset,
	io_in_a_ready,
	io_in_a_valid,
	io_in_a_bits_opcode,
	io_in_a_bits_size,
	io_in_a_bits_source,
	io_in_a_bits_address,
	io_in_a_bits_mask,
	io_in_d_ready,
	io_in_d_valid,
	io_in_d_bits_opcode,
	io_in_d_bits_param,
	io_in_d_bits_size,
	io_in_d_bits_source,
	io_in_d_bits_sink,
	io_in_d_bits_denied,
	io_in_d_bits_corrupt
);
	input clock;
	input reset;
	input io_in_a_ready;
	input io_in_a_valid;
	input [2:0] io_in_a_bits_opcode;
	input [3:0] io_in_a_bits_size;
	input [5:0] io_in_a_bits_source;
	input [31:0] io_in_a_bits_address;
	input [7:0] io_in_a_bits_mask;
	input io_in_d_ready;
	input io_in_d_valid;
	input [2:0] io_in_d_bits_opcode;
	input [1:0] io_in_d_bits_param;
	input [3:0] io_in_d_bits_size;
	input [5:0] io_in_d_bits_source;
	input [2:0] io_in_d_bits_sink;
	input io_in_d_bits_denied;
	input io_in_d_bits_corrupt;
	wire [31:0] _plusarg_reader_1_out;
	wire [31:0] _plusarg_reader_out;
	wire [26:0] _GEN = {23'h000000, io_in_a_bits_size};
	wire _a_first_T_1 = io_in_a_ready & io_in_a_valid;
	reg [8:0] a_first_counter;
	reg [2:0] opcode;
	reg [3:0] size;
	reg [5:0] source;
	reg [31:0] address;
	reg [8:0] d_first_counter;
	reg [2:0] opcode_1;
	reg [1:0] param_1;
	reg [3:0] size_1;
	reg [5:0] source_1;
	reg [2:0] sink;
	reg denied;
	reg [63:0] inflight;
	reg [255:0] inflight_opcodes;
	reg [511:0] inflight_sizes;
	reg [8:0] a_first_counter_1;
	wire a_first_1 = a_first_counter_1 == 9'h000;
	reg [8:0] d_first_counter_1;
	wire d_first_1 = d_first_counter_1 == 9'h000;
	wire [63:0] _GEN_0 = {58'h000000000000000, io_in_a_bits_source};
	wire _GEN_1 = _a_first_T_1 & a_first_1;
	wire d_release_ack = io_in_d_bits_opcode == 3'h6;
	wire [63:0] _GEN_2 = {58'h000000000000000, io_in_d_bits_source};
	reg [31:0] watchdog;
	reg [63:0] inflight_1;
	reg [511:0] inflight_sizes_1;
	reg [8:0] d_first_counter_2;
	wire d_first_2 = d_first_counter_2 == 9'h000;
	reg [31:0] watchdog_1;
	wire [23:0] _GEN_3 = 24'h951240;
	wire [23:0] _GEN_4 = 24'h911240;
	wire source_ok = ((((((((((((((~(|io_in_a_bits_source[5:2]) | (io_in_a_bits_source[5:2] == 4'h1)) | (io_in_a_bits_source[5:2] == 4'h2)) | (io_in_a_bits_source[5:2] == 4'h3)) | (io_in_a_bits_source[5:2] == 4'h4)) | (io_in_a_bits_source[5:2] == 4'h5)) | (io_in_a_bits_source[5:2] == 4'h6)) | (io_in_a_bits_source[5:2] == 4'h7)) | (io_in_a_bits_source[5:2] == 4'h8)) | (io_in_a_bits_source[5:2] == 4'h9)) | (io_in_a_bits_source[5:2] == 4'ha)) | (io_in_a_bits_source[5:2] == 4'hb)) | (io_in_a_bits_source[5:2] == 4'hc)) | (io_in_a_bits_source[5:2] == 4'hd)) | (io_in_a_bits_source[5:2] == 4'he)) | &io_in_a_bits_source[5:2];
	wire [26:0] _is_aligned_mask_T_1 = 27'h0000fff << _GEN;
	wire [11:0] _GEN_5 = io_in_a_bits_address[11:0] & ~_is_aligned_mask_T_1[11:0];
	wire _mask_T = io_in_a_bits_size > 4'h2;
	wire mask_size = io_in_a_bits_size[1:0] == 2'h2;
	wire mask_acc = _mask_T | (mask_size & ~io_in_a_bits_address[2]);
	wire mask_acc_1 = _mask_T | (mask_size & io_in_a_bits_address[2]);
	wire mask_size_1 = io_in_a_bits_size[1:0] == 2'h1;
	wire mask_eq_2 = ~io_in_a_bits_address[2] & ~io_in_a_bits_address[1];
	wire mask_acc_2 = mask_acc | (mask_size_1 & mask_eq_2);
	wire mask_eq_3 = ~io_in_a_bits_address[2] & io_in_a_bits_address[1];
	wire mask_acc_3 = mask_acc | (mask_size_1 & mask_eq_3);
	wire mask_eq_4 = io_in_a_bits_address[2] & ~io_in_a_bits_address[1];
	wire mask_acc_4 = mask_acc_1 | (mask_size_1 & mask_eq_4);
	wire mask_eq_5 = io_in_a_bits_address[2] & io_in_a_bits_address[1];
	wire mask_acc_5 = mask_acc_1 | (mask_size_1 & mask_eq_5);
	wire [7:0] mask = {mask_acc_5 | (mask_eq_5 & io_in_a_bits_address[0]), mask_acc_5 | (mask_eq_5 & ~io_in_a_bits_address[0]), mask_acc_4 | (mask_eq_4 & io_in_a_bits_address[0]), mask_acc_4 | (mask_eq_4 & ~io_in_a_bits_address[0]), mask_acc_3 | (mask_eq_3 & io_in_a_bits_address[0]), mask_acc_3 | (mask_eq_3 & ~io_in_a_bits_address[0]), mask_acc_2 | (mask_eq_2 & io_in_a_bits_address[0]), mask_acc_2 | (mask_eq_2 & ~io_in_a_bits_address[0])};
	wire _GEN_6 = io_in_a_bits_size < 4'hd;
	wire _GEN_7 = _GEN_6 & (((((((((((((((~(|io_in_a_bits_source[5:2]) | (io_in_a_bits_source[5:2] == 4'h1)) | (io_in_a_bits_source[5:2] == 4'h2)) | (io_in_a_bits_source[5:2] == 4'h3)) | (io_in_a_bits_source[5:2] == 4'h4)) | (io_in_a_bits_source[5:2] == 4'h5)) | (io_in_a_bits_source[5:2] == 4'h6)) | (io_in_a_bits_source[5:2] == 4'h7)) | (io_in_a_bits_source[5:2] == 4'h8)) | (io_in_a_bits_source[5:2] == 4'h9)) | (io_in_a_bits_source[5:2] == 4'ha)) | (io_in_a_bits_source[5:2] == 4'hb)) | (io_in_a_bits_source[5:2] == 4'hc)) | (io_in_a_bits_source[5:2] == 4'hd)) | (io_in_a_bits_source[5:2] == 4'he)) | &io_in_a_bits_source[5:2]);
	wire _GEN_8 = {io_in_a_bits_address[31:28], io_in_a_bits_address[27:16] ^ 12'h800} == 16'h0000;
	wire _GEN_9 = io_in_a_bits_address[31:28] == 4'h8;
	wire _GEN_10 = _GEN_8 | _GEN_9;
	wire _GEN_11 = (_GEN_7 & (io_in_a_bits_size == 4'h6)) & _GEN_10;
	wire _GEN_12 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h6)) & ~reset;
	wire _GEN_13 = io_in_a_bits_mask != 8'hff;
	wire _GEN_14 = (io_in_a_valid & &io_in_a_bits_opcode) & ~reset;
	wire _GEN_15 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h4)) & ~reset;
	wire _GEN_16 = {io_in_a_bits_address[31:14], ~io_in_a_bits_address[13:12]} == 20'h00000;
	wire _GEN_17 = _GEN_6 & _GEN_16;
	wire _GEN_18 = io_in_a_bits_size < 4'h7;
	wire _GEN_19 = io_in_a_bits_address[31:13] == 19'h00000;
	wire _GEN_20 = {io_in_a_bits_address[31:21], io_in_a_bits_address[20:17] ^ 4'h8, io_in_a_bits_address[15:12]} == 19'h00000;
	wire _GEN_21 = {io_in_a_bits_address[31:26], io_in_a_bits_address[25:16] ^ 10'h200} == 16'h0000;
	wire _GEN_22 = {io_in_a_bits_address[31:26], io_in_a_bits_address[25:12] ^ 14'h2010} == 20'h00000;
	wire _GEN_23 = {io_in_a_bits_address[31:28], ~io_in_a_bits_address[27:26]} == 6'h00;
	wire _GEN_24 = {io_in_a_bits_address[31:29], io_in_a_bits_address[28:12] ^ 17'h10020} == 20'h00000;
	wire _GEN_25 = io_in_a_bits_mask != mask;
	wire _GEN_26 = _GEN_7 & (_GEN_17 | (_GEN_18 & (((((((_GEN_19 | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9)));
	wire _GEN_27 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h0)) & ~reset;
	wire _GEN_28 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h1)) & ~reset;
	wire _GEN_29 = (_GEN_7 & (io_in_a_bits_size < 4'h4)) & ((((((((_GEN_19 | _GEN_16) | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9);
	wire _GEN_30 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h2)) & ~reset;
	wire _GEN_31 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h3)) & ~reset;
	wire _GEN_32 = (io_in_a_valid & (io_in_a_bits_opcode == 3'h5)) & ~reset;
	wire source_ok_1 = (((((((((((((((io_in_d_bits_source[5:2] == 4'h0) | (io_in_d_bits_source[5:2] == 4'h1)) | (io_in_d_bits_source[5:2] == 4'h2)) | (io_in_d_bits_source[5:2] == 4'h3)) | (io_in_d_bits_source[5:2] == 4'h4)) | (io_in_d_bits_source[5:2] == 4'h5)) | (io_in_d_bits_source[5:2] == 4'h6)) | (io_in_d_bits_source[5:2] == 4'h7)) | (io_in_d_bits_source[5:2] == 4'h8)) | (io_in_d_bits_source[5:2] == 4'h9)) | (io_in_d_bits_source[5:2] == 4'ha)) | (io_in_d_bits_source[5:2] == 4'hb)) | (io_in_d_bits_source[5:2] == 4'hc)) | (io_in_d_bits_source[5:2] == 4'hd)) | (io_in_d_bits_source[5:2] == 4'he)) | &io_in_d_bits_source[5:2];
	wire _GEN_33 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h6)) & ~reset;
	wire _GEN_34 = io_in_d_bits_size < 4'h3;
	wire _GEN_35 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h4)) & ~reset;
	wire _GEN_36 = io_in_d_bits_param == 2'h2;
	wire _GEN_37 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h5)) & ~reset;
	wire _GEN_38 = ~io_in_d_bits_denied | io_in_d_bits_corrupt;
	wire _GEN_39 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h0)) & ~reset;
	wire _GEN_40 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h1)) & ~reset;
	wire _GEN_41 = (io_in_d_valid & (io_in_d_bits_opcode == 3'h2)) & ~reset;
	wire _GEN_42 = (io_in_a_valid & |a_first_counter) & ~reset;
	wire _GEN_43 = (io_in_d_valid & |d_first_counter) & ~reset;
	wire [255:0] _a_opcode_lookup_T_1 = inflight_opcodes >> {248'h00000000000000000000000000000000000000000000000000000000000000, io_in_d_bits_source, 2'h0};
	wire [511:0] _GEN_44 = {503'h0, io_in_d_bits_source, 3'h0};
	wire _same_cycle_resp_T_1 = io_in_a_valid & a_first_1;
	wire [63:0] a_set_wo_ready = (_same_cycle_resp_T_1 ? 64'h0000000000000001 << _GEN_0 : 64'h0000000000000000);
	wire _GEN_45 = io_in_d_valid & d_first_1;
	wire _GEN_46 = _GEN_45 & ~d_release_ack;
	wire same_cycle_resp = _same_cycle_resp_T_1 & (io_in_a_bits_source == io_in_d_bits_source);
	wire _GEN_47 = (_GEN_46 & same_cycle_resp) & ~reset;
	wire _GEN_48 = (_GEN_46 & ~same_cycle_resp) & ~reset;
	wire [7:0] _GEN_49 = {4'h0, io_in_d_bits_size};
	wire _GEN_50 = ((io_in_d_valid & d_first_2) & d_release_ack) & ~reset;
	wire [63:0] _GEN_51 = inflight >> _GEN_0;
	wire [63:0] _GEN_52 = inflight >> _GEN_2;
	wire [511:0] _a_size_lookup_T_1 = inflight_sizes >> _GEN_44;
	wire [63:0] _GEN_53 = inflight_1 >> _GEN_2;
	wire [511:0] _c_size_lookup_T_1 = inflight_sizes_1 >> _GEN_44;
	always @(posedge clock) begin
		if (_GEN_12 & ~_GEN_11) begin
			$error("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12) begin
			$error("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & ~source_ok) begin
			$error("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & ~_mask_T) begin
			$error("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_12 & _GEN_13) begin
			$error("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~_GEN_11) begin
			$error("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14) begin
			$error("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~source_ok) begin
			$error("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & ~_mask_T) begin
			$error("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14) begin
			$error("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_14 & _GEN_13) begin
			$error("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~_GEN_7) begin
			$error("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~(_GEN_17 | (_GEN_18 & ((((((((_GEN_19 | ({io_in_a_bits_address[31:17], ~io_in_a_bits_address[16]} == 16'h0000)) | _GEN_20) | _GEN_21) | _GEN_22) | _GEN_8) | _GEN_23) | _GEN_24) | _GEN_9)))) begin
			$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Get carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Get address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_15 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Get contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & ~_GEN_26) begin
			$error("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & ~source_ok) begin
			$error("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel PutFull address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_27 & _GEN_25) begin
			$error("Assertion failed: 'A' channel PutFull contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & ~_GEN_26) begin
			$error("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & ~source_ok) begin
			$error("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_28 & |(io_in_a_bits_mask & ~mask)) begin
			$error("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & ~_GEN_29) begin
			$error("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_30 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & ~_GEN_29) begin
			$error("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Logical carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Logical address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_31 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Logical contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & ~(_GEN_7 & (_GEN_17 | (_GEN_18 & _GEN_10)))) begin
			$error("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & ~source_ok) begin
			$error("Assertion failed: 'A' channel Hint carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & |_GEN_5) begin
			$error("Assertion failed: 'A' channel Hint address not aligned to size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_32 & _GEN_25) begin
			$error("Assertion failed: 'A' channel Hint contains invalid mask (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if ((io_in_d_valid & ~reset) & &io_in_d_bits_opcode) begin
			$error("Assertion failed: 'D' channel has invalid opcode (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & _GEN_34) begin
			$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_33 & io_in_d_bits_denied) begin
			$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel Grant carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & _GEN_34) begin
			$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & &io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & _GEN_36) begin
			$error("Assertion failed: 'D' channel Grant carries toN param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_35 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel Grant is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & _GEN_34) begin
			$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & &io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & _GEN_36) begin
			$error("Assertion failed: 'D' channel GrantData carries toN param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_37 & ~_GEN_38) begin
			$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_39 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_40 & ~_GEN_38) begin
			$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & ~source_ok_1) begin
			$error("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & |io_in_d_bits_param) begin
			$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_41 & io_in_d_bits_corrupt) begin
			$error("Assertion failed: 'D' channel HintAck is corrupt (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_opcode != opcode)) begin
			$error("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_size != size)) begin
			$error("Assertion failed: 'A' channel size changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_source != source)) begin
			$error("Assertion failed: 'A' channel source changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_42 & (io_in_a_bits_address != address)) begin
			$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_opcode != opcode_1)) begin
			$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_param != param_1)) begin
			$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_size != size_1)) begin
			$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_source != source_1)) begin
			$error("Assertion failed: 'D' channel source changed within multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_sink != sink)) begin
			$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_43 & (io_in_d_bits_denied != denied)) begin
			$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if ((_GEN_1 & ~reset) & _GEN_51[0]) begin
			$error("Assertion failed: 'A' channel re-used a source ID (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if ((_GEN_46 & ~reset) & ~(_GEN_52[0] | same_cycle_resp)) begin
			$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_47 & ~((io_in_d_bits_opcode == _GEN_4[io_in_a_bits_opcode * 3+:3]) | (io_in_d_bits_opcode == _GEN_3[io_in_a_bits_opcode * 3+:3]))) begin
			$error("Assertion failed: 'D' channel contains improper opcode response (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_47 & (io_in_a_bits_size != io_in_d_bits_size)) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_48 & ~((io_in_d_bits_opcode == _GEN_4[_a_opcode_lookup_T_1[3:1] * 3+:3]) | (io_in_d_bits_opcode == _GEN_3[_a_opcode_lookup_T_1[3:1] * 3+:3]))) begin
			$error("Assertion failed: 'D' channel contains improper opcode response (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_48 & (_GEN_49 != {1'h0, _a_size_lookup_T_1[7:1]})) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if ((((((_GEN_45 & a_first_1) & io_in_a_valid) & (io_in_a_bits_source == io_in_d_bits_source)) & ~d_release_ack) & ~reset) & ~(~io_in_d_ready | io_in_a_ready)) begin
			$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~((a_set_wo_ready != (_GEN_46 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000)) | (a_set_wo_ready == 64'h0000000000000000))) begin
			$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency > 0 (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~(((inflight == 64'h0000000000000000) | (_plusarg_reader_out == 32'h00000000)) | (watchdog < _plusarg_reader_out))) begin
			$error("Assertion failed: TileLink timeout expired (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_50 & ~_GEN_53[0]) begin
			$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (_GEN_50 & (_GEN_49 != {1'h0, _c_size_lookup_T_1[7:1]})) begin
			$error("Assertion failed: 'D' channel contains improper response size (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:49 assert(cond, message)\n");
			$fatal;
		end
		if (~reset & ~(((inflight_1 == 64'h0000000000000000) | (_plusarg_reader_1_out == 32'h00000000)) | (watchdog_1 < _plusarg_reader_1_out))) begin
			$error("Assertion failed: TileLink timeout expired (connected at generators/cva6/src/main/scala/cva6/CVA6Tile.scala:192:5)\n    at Monitor.scala:42 assert(cond, message)\n");
			$fatal;
		end
	end
	wire [26:0] _a_first_beats1_decode_T_1 = 27'h0000fff << _GEN;
	wire [26:0] _a_first_beats1_decode_T_5 = 27'h0000fff << _GEN;
	wire [26:0] _GEN_54 = {23'h000000, io_in_d_bits_size};
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << _GEN_54;
	wire [26:0] _d_first_beats1_decode_T_5 = 27'h0000fff << _GEN_54;
	wire [26:0] _d_first_beats1_decode_T_9 = 27'h0000fff << _GEN_54;
	wire [526:0] _GEN_55 = {518'h0, io_in_d_bits_source, 3'h0};
	wire [526:0] _d_opcodes_clr_T_5 = 527'hf << {519'h0, io_in_d_bits_source, 2'h0};
	wire [514:0] _a_opcodes_set_T_1 = {511'h0, (_GEN_1 ? {io_in_a_bits_opcode, 1'h1} : 4'h0)} << {507'h0, io_in_a_bits_source, 2'h0};
	wire [526:0] _d_sizes_clr_T_5 = 527'hff << _GEN_55;
	wire [515:0] _a_sizes_set_T_1 = {511'h0, (_GEN_1 ? {io_in_a_bits_size, 1'h1} : 5'h00)} << {507'h0, io_in_a_bits_source, 3'h0};
	wire [526:0] _d_sizes_clr_T_11 = 527'hff << _GEN_55;
	wire _d_first_T_2 = io_in_d_ready & io_in_d_valid;
	wire _GEN_56 = (_d_first_T_2 & d_first_1) & ~d_release_ack;
	wire _GEN_57 = (_d_first_T_2 & d_first_2) & d_release_ack;
	always @(posedge clock) begin
		if (reset) begin
			a_first_counter <= 9'h000;
			d_first_counter <= 9'h000;
			inflight <= 64'h0000000000000000;
			inflight_opcodes <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
			inflight_sizes <= 512'h0;
			a_first_counter_1 <= 9'h000;
			d_first_counter_1 <= 9'h000;
			watchdog <= 32'h00000000;
			inflight_1 <= 64'h0000000000000000;
			inflight_sizes_1 <= 512'h0;
			d_first_counter_2 <= 9'h000;
			watchdog_1 <= 32'h00000000;
		end
		else begin
			if (_a_first_T_1) begin
				if (|a_first_counter)
					a_first_counter <= a_first_counter - 9'h001;
				else
					a_first_counter <= (io_in_a_bits_opcode[2] ? 9'h000 : ~_a_first_beats1_decode_T_1[11:3]);
				if (a_first_1)
					a_first_counter_1 <= (io_in_a_bits_opcode[2] ? 9'h000 : ~_a_first_beats1_decode_T_5[11:3]);
				else
					a_first_counter_1 <= a_first_counter_1 - 9'h001;
			end
			if (_d_first_T_2) begin
				if (|d_first_counter)
					d_first_counter <= d_first_counter - 9'h001;
				else
					d_first_counter <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_1[11:3] : 9'h000);
				if (d_first_1)
					d_first_counter_1 <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_5[11:3] : 9'h000);
				else
					d_first_counter_1 <= d_first_counter_1 - 9'h001;
				if (d_first_2)
					d_first_counter_2 <= (io_in_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_9[11:3] : 9'h000);
				else
					d_first_counter_2 <= d_first_counter_2 - 9'h001;
				watchdog_1 <= 32'h00000000;
			end
			else
				watchdog_1 <= watchdog_1 + 32'h00000001;
			inflight <= (inflight | (_GEN_1 ? 64'h0000000000000001 << _GEN_0 : 64'h0000000000000000)) & ~(_GEN_56 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000);
			inflight_opcodes <= (inflight_opcodes | (_GEN_1 ? _a_opcodes_set_T_1[255:0] : 256'h0000000000000000000000000000000000000000000000000000000000000000)) & ~(_GEN_56 ? _d_opcodes_clr_T_5[255:0] : 256'h0000000000000000000000000000000000000000000000000000000000000000);
			inflight_sizes <= (inflight_sizes | (_GEN_1 ? _a_sizes_set_T_1[511:0] : 512'h0)) & ~(_GEN_56 ? _d_sizes_clr_T_5[511:0] : 512'h0);
			if (_a_first_T_1 | _d_first_T_2)
				watchdog <= 32'h00000000;
			else
				watchdog <= watchdog + 32'h00000001;
			inflight_1 <= inflight_1 & ~(_GEN_57 ? 64'h0000000000000001 << _GEN_2 : 64'h0000000000000000);
			inflight_sizes_1 <= inflight_sizes_1 & ~(_GEN_57 ? _d_sizes_clr_T_11[511:0] : 512'h0);
		end
		if (_a_first_T_1 & ~(|a_first_counter)) begin
			opcode <= io_in_a_bits_opcode;
			size <= io_in_a_bits_size;
			source <= io_in_a_bits_source;
			address <= io_in_a_bits_address;
		end
		if (_d_first_T_2 & ~(|d_first_counter)) begin
			opcode_1 <= io_in_d_bits_opcode;
			param_1 <= io_in_d_bits_param;
			size_1 <= io_in_d_bits_size;
			source_1 <= io_in_d_bits_source;
			sink <= io_in_d_bits_sink;
			denied <= io_in_d_bits_denied;
		end
	end
	wire [31:0] _RANDOM [0:57];
	plusarg_reader #(
		.DEFAULT(0),
		.FORMAT("tilelink_timeout=%d"),
		.WIDTH(32)
	) plusarg_reader(.out(_plusarg_reader_out));
	plusarg_reader #(
		.DEFAULT(0),
		.FORMAT("tilelink_timeout=%d"),
		.WIDTH(32)
	) plusarg_reader_1(.out(_plusarg_reader_1_out));
endmodule
module TLFIFOFixer_5 (
	clock,
	reset,
	auto_in_a_ready,
	auto_in_a_valid,
	auto_in_a_bits_opcode,
	auto_in_a_bits_size,
	auto_in_a_bits_source,
	auto_in_a_bits_address,
	auto_in_a_bits_mask,
	auto_in_a_bits_data,
	auto_in_d_ready,
	auto_in_d_valid,
	auto_in_d_bits_opcode,
	auto_in_d_bits_size,
	auto_in_d_bits_source,
	auto_in_d_bits_denied,
	auto_in_d_bits_data,
	auto_in_d_bits_corrupt,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_param,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_sink,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_a_ready;
	input auto_in_a_valid;
	input [2:0] auto_in_a_bits_opcode;
	input [3:0] auto_in_a_bits_size;
	input [5:0] auto_in_a_bits_source;
	input [31:0] auto_in_a_bits_address;
	input [7:0] auto_in_a_bits_mask;
	input [63:0] auto_in_a_bits_data;
	input auto_in_d_ready;
	output wire auto_in_d_valid;
	output wire [2:0] auto_in_d_bits_opcode;
	output wire [3:0] auto_in_d_bits_size;
	output wire [5:0] auto_in_d_bits_source;
	output wire auto_in_d_bits_denied;
	output wire [63:0] auto_in_d_bits_data;
	output wire auto_in_d_bits_corrupt;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [3:0] auto_out_a_bits_size;
	output wire [5:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [1:0] auto_out_d_bits_param;
	input [3:0] auto_out_d_bits_size;
	input [5:0] auto_out_d_bits_source;
	input [2:0] auto_out_d_bits_sink;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire a_id = (({auto_in_a_bits_address[31], auto_in_a_bits_address[27:26]} == 3'h0) | ({auto_in_a_bits_address[31], auto_in_a_bits_address[27:26], ~auto_in_a_bits_address[16], auto_in_a_bits_address[12]} == 5'h00)) | ({auto_in_a_bits_address[31], ~auto_in_a_bits_address[27:26]} == 3'h0);
	reg [8:0] a_first_counter;
	wire a_first = a_first_counter == 9'h000;
	reg [8:0] d_first_counter;
	reg flight_0;
	reg flight_1;
	reg flight_2;
	reg flight_3;
	reg flight_4;
	reg flight_5;
	reg flight_6;
	reg flight_7;
	reg flight_8;
	reg flight_9;
	reg flight_10;
	reg flight_11;
	reg flight_12;
	reg flight_13;
	reg flight_14;
	reg flight_15;
	reg flight_16;
	reg flight_17;
	reg flight_18;
	reg flight_19;
	reg flight_20;
	reg flight_21;
	reg flight_22;
	reg flight_23;
	reg flight_24;
	reg flight_25;
	reg flight_26;
	reg flight_27;
	reg flight_28;
	reg flight_29;
	reg flight_30;
	reg flight_31;
	reg flight_32;
	reg flight_33;
	reg flight_34;
	reg flight_35;
	reg flight_36;
	reg flight_37;
	reg flight_38;
	reg flight_39;
	reg flight_40;
	reg flight_41;
	reg flight_42;
	reg flight_43;
	reg flight_44;
	reg flight_45;
	reg flight_46;
	reg flight_47;
	reg flight_48;
	reg flight_49;
	reg flight_50;
	reg flight_51;
	reg flight_52;
	reg flight_53;
	reg flight_54;
	reg flight_55;
	reg flight_56;
	reg flight_57;
	reg flight_58;
	reg flight_59;
	reg flight_60;
	reg flight_61;
	reg flight_62;
	reg flight_63;
	wire stalls_a_sel = auto_in_a_bits_source[5:2] == 4'h0;
	reg stalls_id;
	wire stalls_a_sel_1 = auto_in_a_bits_source[5:2] == 4'h1;
	reg stalls_id_1;
	wire stalls_a_sel_2 = auto_in_a_bits_source[5:2] == 4'h2;
	reg stalls_id_2;
	wire stalls_a_sel_3 = auto_in_a_bits_source[5:2] == 4'h3;
	reg stalls_id_3;
	wire stalls_a_sel_4 = auto_in_a_bits_source[5:2] == 4'h4;
	reg stalls_id_4;
	wire stalls_a_sel_5 = auto_in_a_bits_source[5:2] == 4'h5;
	reg stalls_id_5;
	wire stalls_a_sel_6 = auto_in_a_bits_source[5:2] == 4'h6;
	reg stalls_id_6;
	wire stalls_a_sel_7 = auto_in_a_bits_source[5:2] == 4'h7;
	reg stalls_id_7;
	wire stalls_a_sel_8 = auto_in_a_bits_source[5:2] == 4'h8;
	reg stalls_id_8;
	wire stalls_a_sel_9 = auto_in_a_bits_source[5:2] == 4'h9;
	reg stalls_id_9;
	wire stalls_a_sel_10 = auto_in_a_bits_source[5:2] == 4'ha;
	reg stalls_id_10;
	wire stalls_a_sel_11 = auto_in_a_bits_source[5:2] == 4'hb;
	reg stalls_id_11;
	wire stalls_a_sel_12 = auto_in_a_bits_source[5:2] == 4'hc;
	reg stalls_id_12;
	wire stalls_a_sel_13 = auto_in_a_bits_source[5:2] == 4'hd;
	reg stalls_id_13;
	wire stalls_a_sel_14 = auto_in_a_bits_source[5:2] == 4'he;
	reg stalls_id_14;
	reg stalls_id_15;
	wire stall = (((((((((((((((((stalls_a_sel & a_first) & (((flight_0 | flight_1) | flight_2) | flight_3)) & (~a_id | (stalls_id != a_id))) | (((stalls_a_sel_1 & a_first) & (((flight_4 | flight_5) | flight_6) | flight_7)) & (~a_id | (stalls_id_1 != a_id)))) | (((stalls_a_sel_2 & a_first) & (((flight_8 | flight_9) | flight_10) | flight_11)) & (~a_id | (stalls_id_2 != a_id)))) | (((stalls_a_sel_3 & a_first) & (((flight_12 | flight_13) | flight_14) | flight_15)) & (~a_id | (stalls_id_3 != a_id)))) | (((stalls_a_sel_4 & a_first) & (((flight_16 | flight_17) | flight_18) | flight_19)) & (~a_id | (stalls_id_4 != a_id)))) | (((stalls_a_sel_5 & a_first) & (((flight_20 | flight_21) | flight_22) | flight_23)) & (~a_id | (stalls_id_5 != a_id)))) | (((stalls_a_sel_6 & a_first) & (((flight_24 | flight_25) | flight_26) | flight_27)) & (~a_id | (stalls_id_6 != a_id)))) | (((stalls_a_sel_7 & a_first) & (((flight_28 | flight_29) | flight_30) | flight_31)) & (~a_id | (stalls_id_7 != a_id)))) | (((stalls_a_sel_8 & a_first) & (((flight_32 | flight_33) | flight_34) | flight_35)) & (~a_id | (stalls_id_8 != a_id)))) | (((stalls_a_sel_9 & a_first) & (((flight_36 | flight_37) | flight_38) | flight_39)) & (~a_id | (stalls_id_9 != a_id)))) | (((stalls_a_sel_10 & a_first) & (((flight_40 | flight_41) | flight_42) | flight_43)) & (~a_id | (stalls_id_10 != a_id)))) | (((stalls_a_sel_11 & a_first) & (((flight_44 | flight_45) | flight_46) | flight_47)) & (~a_id | (stalls_id_11 != a_id)))) | (((stalls_a_sel_12 & a_first) & (((flight_48 | flight_49) | flight_50) | flight_51)) & (~a_id | (stalls_id_12 != a_id)))) | (((stalls_a_sel_13 & a_first) & (((flight_52 | flight_53) | flight_54) | flight_55)) & (~a_id | (stalls_id_13 != a_id)))) | (((stalls_a_sel_14 & a_first) & (((flight_56 | flight_57) | flight_58) | flight_59)) & (~a_id | (stalls_id_14 != a_id)))) | (((&auto_in_a_bits_source[5:2] & a_first) & (((flight_60 | flight_61) | flight_62) | flight_63)) & (~a_id | (stalls_id_15 != a_id)));
	wire nodeIn_a_ready = auto_out_a_ready & ~stall;
	wire [26:0] _a_first_beats1_decode_T_1 = 27'h0000fff << auto_in_a_bits_size;
	wire [26:0] _d_first_beats1_decode_T_1 = 27'h0000fff << auto_out_d_bits_size;
	wire d_first_first = d_first_counter == 9'h000;
	wire _GEN = ((d_first_first & (auto_out_d_bits_opcode != 3'h6)) & auto_in_d_ready) & auto_out_d_valid;
	wire _stalls_id_T_60 = nodeIn_a_ready & auto_in_a_valid;
	wire _GEN_0 = a_first & _stalls_id_T_60;
	always @(posedge clock) begin
		if (reset) begin
			a_first_counter <= 9'h000;
			d_first_counter <= 9'h000;
			flight_0 <= 1'h0;
			flight_1 <= 1'h0;
			flight_2 <= 1'h0;
			flight_3 <= 1'h0;
			flight_4 <= 1'h0;
			flight_5 <= 1'h0;
			flight_6 <= 1'h0;
			flight_7 <= 1'h0;
			flight_8 <= 1'h0;
			flight_9 <= 1'h0;
			flight_10 <= 1'h0;
			flight_11 <= 1'h0;
			flight_12 <= 1'h0;
			flight_13 <= 1'h0;
			flight_14 <= 1'h0;
			flight_15 <= 1'h0;
			flight_16 <= 1'h0;
			flight_17 <= 1'h0;
			flight_18 <= 1'h0;
			flight_19 <= 1'h0;
			flight_20 <= 1'h0;
			flight_21 <= 1'h0;
			flight_22 <= 1'h0;
			flight_23 <= 1'h0;
			flight_24 <= 1'h0;
			flight_25 <= 1'h0;
			flight_26 <= 1'h0;
			flight_27 <= 1'h0;
			flight_28 <= 1'h0;
			flight_29 <= 1'h0;
			flight_30 <= 1'h0;
			flight_31 <= 1'h0;
			flight_32 <= 1'h0;
			flight_33 <= 1'h0;
			flight_34 <= 1'h0;
			flight_35 <= 1'h0;
			flight_36 <= 1'h0;
			flight_37 <= 1'h0;
			flight_38 <= 1'h0;
			flight_39 <= 1'h0;
			flight_40 <= 1'h0;
			flight_41 <= 1'h0;
			flight_42 <= 1'h0;
			flight_43 <= 1'h0;
			flight_44 <= 1'h0;
			flight_45 <= 1'h0;
			flight_46 <= 1'h0;
			flight_47 <= 1'h0;
			flight_48 <= 1'h0;
			flight_49 <= 1'h0;
			flight_50 <= 1'h0;
			flight_51 <= 1'h0;
			flight_52 <= 1'h0;
			flight_53 <= 1'h0;
			flight_54 <= 1'h0;
			flight_55 <= 1'h0;
			flight_56 <= 1'h0;
			flight_57 <= 1'h0;
			flight_58 <= 1'h0;
			flight_59 <= 1'h0;
			flight_60 <= 1'h0;
			flight_61 <= 1'h0;
			flight_62 <= 1'h0;
			flight_63 <= 1'h0;
		end
		else begin
			if (_stalls_id_T_60) begin
				if (a_first)
					a_first_counter <= (auto_in_a_bits_opcode[2] ? 9'h000 : ~_a_first_beats1_decode_T_1[11:3]);
				else
					a_first_counter <= a_first_counter - 9'h001;
			end
			if (auto_in_d_ready & auto_out_d_valid) begin
				if (d_first_first)
					d_first_counter <= (auto_out_d_bits_opcode[0] ? ~_d_first_beats1_decode_T_1[11:3] : 9'h000);
				else
					d_first_counter <= d_first_counter - 9'h001;
			end
			flight_0 <= ~(_GEN & (auto_out_d_bits_source == 6'h00)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h00)) | flight_0);
			flight_1 <= ~(_GEN & (auto_out_d_bits_source == 6'h01)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h01)) | flight_1);
			flight_2 <= ~(_GEN & (auto_out_d_bits_source == 6'h02)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h02)) | flight_2);
			flight_3 <= ~(_GEN & (auto_out_d_bits_source == 6'h03)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h03)) | flight_3);
			flight_4 <= ~(_GEN & (auto_out_d_bits_source == 6'h04)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h04)) | flight_4);
			flight_5 <= ~(_GEN & (auto_out_d_bits_source == 6'h05)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h05)) | flight_5);
			flight_6 <= ~(_GEN & (auto_out_d_bits_source == 6'h06)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h06)) | flight_6);
			flight_7 <= ~(_GEN & (auto_out_d_bits_source == 6'h07)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h07)) | flight_7);
			flight_8 <= ~(_GEN & (auto_out_d_bits_source == 6'h08)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h08)) | flight_8);
			flight_9 <= ~(_GEN & (auto_out_d_bits_source == 6'h09)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h09)) | flight_9);
			flight_10 <= ~(_GEN & (auto_out_d_bits_source == 6'h0a)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0a)) | flight_10);
			flight_11 <= ~(_GEN & (auto_out_d_bits_source == 6'h0b)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0b)) | flight_11);
			flight_12 <= ~(_GEN & (auto_out_d_bits_source == 6'h0c)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0c)) | flight_12);
			flight_13 <= ~(_GEN & (auto_out_d_bits_source == 6'h0d)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0d)) | flight_13);
			flight_14 <= ~(_GEN & (auto_out_d_bits_source == 6'h0e)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0e)) | flight_14);
			flight_15 <= ~(_GEN & (auto_out_d_bits_source == 6'h0f)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h0f)) | flight_15);
			flight_16 <= ~(_GEN & (auto_out_d_bits_source == 6'h10)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h10)) | flight_16);
			flight_17 <= ~(_GEN & (auto_out_d_bits_source == 6'h11)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h11)) | flight_17);
			flight_18 <= ~(_GEN & (auto_out_d_bits_source == 6'h12)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h12)) | flight_18);
			flight_19 <= ~(_GEN & (auto_out_d_bits_source == 6'h13)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h13)) | flight_19);
			flight_20 <= ~(_GEN & (auto_out_d_bits_source == 6'h14)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h14)) | flight_20);
			flight_21 <= ~(_GEN & (auto_out_d_bits_source == 6'h15)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h15)) | flight_21);
			flight_22 <= ~(_GEN & (auto_out_d_bits_source == 6'h16)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h16)) | flight_22);
			flight_23 <= ~(_GEN & (auto_out_d_bits_source == 6'h17)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h17)) | flight_23);
			flight_24 <= ~(_GEN & (auto_out_d_bits_source == 6'h18)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h18)) | flight_24);
			flight_25 <= ~(_GEN & (auto_out_d_bits_source == 6'h19)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h19)) | flight_25);
			flight_26 <= ~(_GEN & (auto_out_d_bits_source == 6'h1a)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1a)) | flight_26);
			flight_27 <= ~(_GEN & (auto_out_d_bits_source == 6'h1b)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1b)) | flight_27);
			flight_28 <= ~(_GEN & (auto_out_d_bits_source == 6'h1c)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1c)) | flight_28);
			flight_29 <= ~(_GEN & (auto_out_d_bits_source == 6'h1d)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1d)) | flight_29);
			flight_30 <= ~(_GEN & (auto_out_d_bits_source == 6'h1e)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1e)) | flight_30);
			flight_31 <= ~(_GEN & (auto_out_d_bits_source == 6'h1f)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h1f)) | flight_31);
			flight_32 <= ~(_GEN & (auto_out_d_bits_source == 6'h20)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h20)) | flight_32);
			flight_33 <= ~(_GEN & (auto_out_d_bits_source == 6'h21)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h21)) | flight_33);
			flight_34 <= ~(_GEN & (auto_out_d_bits_source == 6'h22)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h22)) | flight_34);
			flight_35 <= ~(_GEN & (auto_out_d_bits_source == 6'h23)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h23)) | flight_35);
			flight_36 <= ~(_GEN & (auto_out_d_bits_source == 6'h24)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h24)) | flight_36);
			flight_37 <= ~(_GEN & (auto_out_d_bits_source == 6'h25)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h25)) | flight_37);
			flight_38 <= ~(_GEN & (auto_out_d_bits_source == 6'h26)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h26)) | flight_38);
			flight_39 <= ~(_GEN & (auto_out_d_bits_source == 6'h27)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h27)) | flight_39);
			flight_40 <= ~(_GEN & (auto_out_d_bits_source == 6'h28)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h28)) | flight_40);
			flight_41 <= ~(_GEN & (auto_out_d_bits_source == 6'h29)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h29)) | flight_41);
			flight_42 <= ~(_GEN & (auto_out_d_bits_source == 6'h2a)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2a)) | flight_42);
			flight_43 <= ~(_GEN & (auto_out_d_bits_source == 6'h2b)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2b)) | flight_43);
			flight_44 <= ~(_GEN & (auto_out_d_bits_source == 6'h2c)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2c)) | flight_44);
			flight_45 <= ~(_GEN & (auto_out_d_bits_source == 6'h2d)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2d)) | flight_45);
			flight_46 <= ~(_GEN & (auto_out_d_bits_source == 6'h2e)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2e)) | flight_46);
			flight_47 <= ~(_GEN & (auto_out_d_bits_source == 6'h2f)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h2f)) | flight_47);
			flight_48 <= ~(_GEN & (auto_out_d_bits_source == 6'h30)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h30)) | flight_48);
			flight_49 <= ~(_GEN & (auto_out_d_bits_source == 6'h31)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h31)) | flight_49);
			flight_50 <= ~(_GEN & (auto_out_d_bits_source == 6'h32)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h32)) | flight_50);
			flight_51 <= ~(_GEN & (auto_out_d_bits_source == 6'h33)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h33)) | flight_51);
			flight_52 <= ~(_GEN & (auto_out_d_bits_source == 6'h34)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h34)) | flight_52);
			flight_53 <= ~(_GEN & (auto_out_d_bits_source == 6'h35)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h35)) | flight_53);
			flight_54 <= ~(_GEN & (auto_out_d_bits_source == 6'h36)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h36)) | flight_54);
			flight_55 <= ~(_GEN & (auto_out_d_bits_source == 6'h37)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h37)) | flight_55);
			flight_56 <= ~(_GEN & (auto_out_d_bits_source == 6'h38)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h38)) | flight_56);
			flight_57 <= ~(_GEN & (auto_out_d_bits_source == 6'h39)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h39)) | flight_57);
			flight_58 <= ~(_GEN & (auto_out_d_bits_source == 6'h3a)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h3a)) | flight_58);
			flight_59 <= ~(_GEN & (auto_out_d_bits_source == 6'h3b)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h3b)) | flight_59);
			flight_60 <= ~(_GEN & (auto_out_d_bits_source == 6'h3c)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h3c)) | flight_60);
			flight_61 <= ~(_GEN & (auto_out_d_bits_source == 6'h3d)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h3d)) | flight_61);
			flight_62 <= ~(_GEN & (auto_out_d_bits_source == 6'h3e)) & ((_GEN_0 & (auto_in_a_bits_source == 6'h3e)) | flight_62);
			flight_63 <= ~(_GEN & &auto_out_d_bits_source) & ((_GEN_0 & &auto_in_a_bits_source) | flight_63);
		end
		if (_stalls_id_T_60 & stalls_a_sel)
			stalls_id <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_1)
			stalls_id_1 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_2)
			stalls_id_2 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_3)
			stalls_id_3 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_4)
			stalls_id_4 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_5)
			stalls_id_5 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_6)
			stalls_id_6 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_7)
			stalls_id_7 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_8)
			stalls_id_8 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_9)
			stalls_id_9 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_10)
			stalls_id_10 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_11)
			stalls_id_11 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_12)
			stalls_id_12 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_13)
			stalls_id_13 <= a_id;
		if (_stalls_id_T_60 & stalls_a_sel_14)
			stalls_id_14 <= a_id;
		if (_stalls_id_T_60 & &auto_in_a_bits_source[5:2])
			stalls_id_15 <= a_id;
	end
	wire [31:0] _RANDOM [0:3];
	TLMonitor_41 monitor(
		.clock(clock),
		.reset(reset),
		.io_in_a_ready(nodeIn_a_ready),
		.io_in_a_valid(auto_in_a_valid),
		.io_in_a_bits_opcode(auto_in_a_bits_opcode),
		.io_in_a_bits_size(auto_in_a_bits_size),
		.io_in_a_bits_source(auto_in_a_bits_source),
		.io_in_a_bits_address(auto_in_a_bits_address),
		.io_in_a_bits_mask(auto_in_a_bits_mask),
		.io_in_d_ready(auto_in_d_ready),
		.io_in_d_valid(auto_out_d_valid),
		.io_in_d_bits_opcode(auto_out_d_bits_opcode),
		.io_in_d_bits_param(auto_out_d_bits_param),
		.io_in_d_bits_size(auto_out_d_bits_size),
		.io_in_d_bits_source(auto_out_d_bits_source),
		.io_in_d_bits_sink(auto_out_d_bits_sink),
		.io_in_d_bits_denied(auto_out_d_bits_denied),
		.io_in_d_bits_corrupt(auto_out_d_bits_corrupt)
	);
	assign auto_in_a_ready = nodeIn_a_ready;
	assign auto_in_d_valid = auto_out_d_valid;
	assign auto_in_d_bits_opcode = auto_out_d_bits_opcode;
	assign auto_in_d_bits_size = auto_out_d_bits_size;
	assign auto_in_d_bits_source = auto_out_d_bits_source;
	assign auto_in_d_bits_denied = auto_out_d_bits_denied;
	assign auto_in_d_bits_data = auto_out_d_bits_data;
	assign auto_in_d_bits_corrupt = auto_out_d_bits_corrupt;
	assign auto_out_a_valid = auto_in_a_valid & ~stall;
	assign auto_out_a_bits_opcode = auto_in_a_bits_opcode;
	assign auto_out_a_bits_size = auto_in_a_bits_size;
	assign auto_out_a_bits_source = auto_in_a_bits_source;
	assign auto_out_a_bits_address = auto_in_a_bits_address;
	assign auto_out_a_bits_mask = auto_in_a_bits_mask;
	assign auto_out_a_bits_data = auto_in_a_bits_data;
	assign auto_out_d_ready = auto_in_d_ready;
endmodule
module Queue_54 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_data,
	io_enq_bits_resp,
	io_enq_bits_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_data,
	io_deq_bits_resp,
	io_deq_bits_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [3:0] io_enq_bits_id;
	input [63:0] io_enq_bits_data;
	input [1:0] io_enq_bits_resp;
	input io_enq_bits_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [3:0] io_deq_bits_id;
	output wire [63:0] io_deq_bits_data;
	output wire [1:0] io_deq_bits_resp;
	output wire io_deq_bits_last;
	reg ram_last;
	reg [1:0] ram_resp;
	reg [63:0] ram_data;
	reg [3:0] ram_id;
	reg full;
	wire _io_deq_valid_output = io_enq_valid | full;
	wire do_enq = (~(~full & io_deq_ready) & ~full) & io_enq_valid;
	always @(posedge clock) begin
		if (do_enq) begin
			ram_last <= io_enq_bits_last;
			ram_resp <= io_enq_bits_resp;
			ram_data <= io_enq_bits_data;
			ram_id <= io_enq_bits_id;
		end
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == ((full & io_deq_ready) & _io_deq_valid_output)))
			full <= do_enq;
	end
	wire [31:0] _RANDOM [0:2];
	assign io_enq_ready = ~full;
	assign io_deq_valid = _io_deq_valid_output;
	assign io_deq_bits_id = (full ? ram_id : io_enq_bits_id);
	assign io_deq_bits_data = (full ? ram_data : io_enq_bits_data);
	assign io_deq_bits_resp = (full ? ram_resp : io_enq_bits_resp);
	assign io_deq_bits_last = (full ? ram_last : io_enq_bits_last);
endmodule
module Queue_55 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_resp,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_resp
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [3:0] io_enq_bits_id;
	input [1:0] io_enq_bits_resp;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [3:0] io_deq_bits_id;
	output wire [1:0] io_deq_bits_resp;
	reg [1:0] ram_resp;
	reg [3:0] ram_id;
	reg full;
	wire _io_deq_valid_output = io_enq_valid | full;
	wire do_enq = (~(~full & io_deq_ready) & ~full) & io_enq_valid;
	always @(posedge clock) begin
		if (do_enq) begin
			ram_resp <= io_enq_bits_resp;
			ram_id <= io_enq_bits_id;
		end
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == ((full & io_deq_ready) & _io_deq_valid_output)))
			full <= do_enq;
	end
	wire [31:0] _RANDOM [0:0];
	assign io_enq_ready = ~full;
	assign io_deq_valid = _io_deq_valid_output;
	assign io_deq_bits_id = (full ? ram_id : io_enq_bits_id);
	assign io_deq_bits_resp = (full ? ram_resp : io_enq_bits_resp);
endmodule
module AXI4ToTL (
	clock,
	reset,
	auto_in_aw_ready,
	auto_in_aw_valid,
	auto_in_aw_bits_id,
	auto_in_aw_bits_addr,
	auto_in_aw_bits_len,
	auto_in_aw_bits_size,
	auto_in_w_ready,
	auto_in_w_valid,
	auto_in_w_bits_data,
	auto_in_w_bits_strb,
	auto_in_w_bits_last,
	auto_in_b_ready,
	auto_in_b_valid,
	auto_in_b_bits_id,
	auto_in_b_bits_resp,
	auto_in_ar_ready,
	auto_in_ar_valid,
	auto_in_ar_bits_id,
	auto_in_ar_bits_addr,
	auto_in_ar_bits_len,
	auto_in_ar_bits_size,
	auto_in_r_ready,
	auto_in_r_valid,
	auto_in_r_bits_id,
	auto_in_r_bits_data,
	auto_in_r_bits_resp,
	auto_in_r_bits_last,
	auto_out_a_ready,
	auto_out_a_valid,
	auto_out_a_bits_opcode,
	auto_out_a_bits_size,
	auto_out_a_bits_source,
	auto_out_a_bits_address,
	auto_out_a_bits_mask,
	auto_out_a_bits_data,
	auto_out_d_ready,
	auto_out_d_valid,
	auto_out_d_bits_opcode,
	auto_out_d_bits_size,
	auto_out_d_bits_source,
	auto_out_d_bits_denied,
	auto_out_d_bits_data,
	auto_out_d_bits_corrupt
);
	input clock;
	input reset;
	output wire auto_in_aw_ready;
	input auto_in_aw_valid;
	input [3:0] auto_in_aw_bits_id;
	input [31:0] auto_in_aw_bits_addr;
	input [7:0] auto_in_aw_bits_len;
	input [2:0] auto_in_aw_bits_size;
	output wire auto_in_w_ready;
	input auto_in_w_valid;
	input [63:0] auto_in_w_bits_data;
	input [7:0] auto_in_w_bits_strb;
	input auto_in_w_bits_last;
	input auto_in_b_ready;
	output wire auto_in_b_valid;
	output wire [3:0] auto_in_b_bits_id;
	output wire [1:0] auto_in_b_bits_resp;
	output wire auto_in_ar_ready;
	input auto_in_ar_valid;
	input [3:0] auto_in_ar_bits_id;
	input [31:0] auto_in_ar_bits_addr;
	input [7:0] auto_in_ar_bits_len;
	input [2:0] auto_in_ar_bits_size;
	input auto_in_r_ready;
	output wire auto_in_r_valid;
	output wire [3:0] auto_in_r_bits_id;
	output wire [63:0] auto_in_r_bits_data;
	output wire [1:0] auto_in_r_bits_resp;
	output wire auto_in_r_bits_last;
	input auto_out_a_ready;
	output wire auto_out_a_valid;
	output wire [2:0] auto_out_a_bits_opcode;
	output wire [3:0] auto_out_a_bits_size;
	output wire [5:0] auto_out_a_bits_source;
	output wire [31:0] auto_out_a_bits_address;
	output wire [7:0] auto_out_a_bits_mask;
	output wire [63:0] auto_out_a_bits_data;
	output wire auto_out_d_ready;
	input auto_out_d_valid;
	input [2:0] auto_out_d_bits_opcode;
	input [3:0] auto_out_d_bits_size;
	input [5:0] auto_out_d_bits_source;
	input auto_out_d_bits_denied;
	input [63:0] auto_out_d_bits_data;
	input auto_out_d_bits_corrupt;
	wire w_out_ready;
	wire _q_b_deq_q_io_enq_ready;
	wire _q_b_deq_q_io_deq_valid;
	wire [3:0] _q_b_deq_q_io_deq_bits_id;
	wire _nodeIn_r_deq_q_io_enq_ready;
	wire [22:0] _r_size1_T_1 = {7'h00, auto_in_ar_bits_len, 8'hff} << auto_in_ar_bits_size;
	wire [13:0] _GEN = ~_r_size1_T_1[22:9];
	wire [7:0] r_size_hi = _r_size1_T_1[22:15] & {1'h1, _GEN[13:7]};
	wire [6:0] _r_size_T_6 = r_size_hi[7:1] | (_r_size1_T_1[14:8] & _GEN[6:0]);
	wire [2:0] _r_size_T_8 = _r_size_T_6[6:4] | _r_size_T_6[2:0];
	wire _r_size_T_10 = _r_size_T_8[2] | _r_size_T_8[0];
	wire [3:0] r_out_bits_a_size = {|r_size_hi, |_r_size_T_6[6:3], |_r_size_T_8[2:1], _r_size_T_10};
	wire [31:0] r_out_bits_a_address = (((r_out_bits_a_size < 4'hd) & ({auto_in_ar_bits_addr[31:14], ~auto_in_ar_bits_addr[13:12]} == 20'h00000)) | ((r_out_bits_a_size < 4'h7) & (((((((((auto_in_ar_bits_addr[31:13] == 19'h00000) | ({auto_in_ar_bits_addr[31:17], ~auto_in_ar_bits_addr[16]} == 16'h0000)) | ({auto_in_ar_bits_addr[31:21], auto_in_ar_bits_addr[20:17] ^ 4'h8, auto_in_ar_bits_addr[15:12]} == 19'h00000)) | ({auto_in_ar_bits_addr[31:26], auto_in_ar_bits_addr[25:16] ^ 10'h200} == 16'h0000)) | ({auto_in_ar_bits_addr[31:26], auto_in_ar_bits_addr[25:12] ^ 14'h2010} == 20'h00000)) | ({auto_in_ar_bits_addr[31:28], auto_in_ar_bits_addr[27:16] ^ 12'h800} == 16'h0000)) | ({auto_in_ar_bits_addr[31:28], ~auto_in_ar_bits_addr[27:26]} == 6'h00)) | ({auto_in_ar_bits_addr[31:29], auto_in_ar_bits_addr[28:12] ^ 17'h10020} == 20'h00000)) | (auto_in_ar_bits_addr[31:28] == 4'h8))) ? auto_in_ar_bits_addr : {29'h00000600, auto_in_ar_bits_addr[2:0]});
	reg [1:0] r_count_0;
	reg [1:0] r_count_1;
	reg [1:0] r_count_2;
	reg [1:0] r_count_3;
	reg [1:0] r_count_4;
	reg [1:0] r_count_5;
	reg [1:0] r_count_6;
	reg [1:0] r_count_7;
	reg [1:0] r_count_8;
	reg [1:0] r_count_9;
	reg [1:0] r_count_10;
	reg [1:0] r_count_11;
	reg [1:0] r_count_12;
	reg [1:0] r_count_13;
	reg [1:0] r_count_14;
	reg [1:0] r_count_15;
	wire [31:0] _GEN_0 = {r_count_15, r_count_14, r_count_13, r_count_12, r_count_11, r_count_10, r_count_9, r_count_8, r_count_7, r_count_6, r_count_5, r_count_4, r_count_3, r_count_2, r_count_1, r_count_0};
	wire _r_out_bits_a_mask_T = r_out_bits_a_size > 4'h2;
	wire [1:0] _GEN_1 = {|_r_size_T_8[2:1], _r_size_T_10};
	wire r_out_bits_a_mask_size = _GEN_1 == 2'h2;
	wire r_out_bits_a_mask_acc = _r_out_bits_a_mask_T | (r_out_bits_a_mask_size & ~r_out_bits_a_address[2]);
	wire r_out_bits_a_mask_acc_1 = _r_out_bits_a_mask_T | (r_out_bits_a_mask_size & r_out_bits_a_address[2]);
	wire r_out_bits_a_mask_size_1 = _GEN_1 == 2'h1;
	wire r_out_bits_a_mask_eq_2 = ~r_out_bits_a_address[2] & ~r_out_bits_a_address[1];
	wire r_out_bits_a_mask_acc_2 = r_out_bits_a_mask_acc | (r_out_bits_a_mask_size_1 & r_out_bits_a_mask_eq_2);
	wire r_out_bits_a_mask_eq_3 = ~r_out_bits_a_address[2] & r_out_bits_a_address[1];
	wire r_out_bits_a_mask_acc_3 = r_out_bits_a_mask_acc | (r_out_bits_a_mask_size_1 & r_out_bits_a_mask_eq_3);
	wire r_out_bits_a_mask_eq_4 = r_out_bits_a_address[2] & ~r_out_bits_a_address[1];
	wire r_out_bits_a_mask_acc_4 = r_out_bits_a_mask_acc_1 | (r_out_bits_a_mask_size_1 & r_out_bits_a_mask_eq_4);
	wire r_out_bits_a_mask_eq_5 = r_out_bits_a_address[2] & r_out_bits_a_address[1];
	wire r_out_bits_a_mask_acc_5 = r_out_bits_a_mask_acc_1 | (r_out_bits_a_mask_size_1 & r_out_bits_a_mask_eq_5);
	wire [22:0] _w_size1_T_1 = {7'h00, auto_in_aw_bits_len, 8'hff} << auto_in_aw_bits_size;
	wire [13:0] _GEN_2 = ~_w_size1_T_1[22:9];
	wire [7:0] w_size_hi = _w_size1_T_1[22:15] & {1'h1, _GEN_2[13:7]};
	wire [6:0] _w_size_T_6 = w_size_hi[7:1] | (_w_size1_T_1[14:8] & _GEN_2[6:0]);
	wire [2:0] _w_size_T_8 = _w_size_T_6[6:4] | _w_size_T_6[2:0];
	wire _w_size_T_10 = _w_size_T_8[2] | _w_size_T_8[0];
	wire [3:0] w_out_bits_a_size = {|w_size_hi, |_w_size_T_6[6:3], |_w_size_T_8[2:1], _w_size_T_10};
	reg [1:0] w_count_0;
	reg [1:0] w_count_1;
	reg [1:0] w_count_2;
	reg [1:0] w_count_3;
	reg [1:0] w_count_4;
	reg [1:0] w_count_5;
	reg [1:0] w_count_6;
	reg [1:0] w_count_7;
	reg [1:0] w_count_8;
	reg [1:0] w_count_9;
	reg [1:0] w_count_10;
	reg [1:0] w_count_11;
	reg [1:0] w_count_12;
	reg [1:0] w_count_13;
	reg [1:0] w_count_14;
	reg [1:0] w_count_15;
	wire [31:0] _GEN_3 = {w_count_15, w_count_14, w_count_13, w_count_12, w_count_11, w_count_10, w_count_9, w_count_8, w_count_7, w_count_6, w_count_5, w_count_4, w_count_3, w_count_2, w_count_1, w_count_0};
	wire nodeIn_aw_ready = (w_out_ready & auto_in_w_valid) & auto_in_w_bits_last;
	wire w_out_valid = auto_in_aw_valid & auto_in_w_valid;
	reg [7:0] beatsLeft;
	wire idle = beatsLeft == 8'h00;
	wire [1:0] readys_valid = {w_out_valid, auto_in_ar_valid};
	reg [1:0] readys_mask;
	wire [1:0] _readys_filter_T_1 = readys_valid & ~readys_mask;
	wire [1:0] readys_readys = ~({readys_mask[1], _readys_filter_T_1[1] | readys_mask[0]} & ({_readys_filter_T_1[0], w_out_valid} | _readys_filter_T_1));
	wire winner_0 = readys_readys[0] & auto_in_ar_valid;
	wire winner_1 = readys_readys[1] & w_out_valid;
	wire _nodeOut_a_valid_T = auto_in_ar_valid | w_out_valid;
	wire [29:0] _GEN_4 = 30'h00007fff << {26'h0000000, |r_size_hi, |_r_size_T_6[6:3], |_r_size_T_8[2:1], _r_size_T_10};
	wire [29:0] _GEN_5 = 30'h00007fff << {26'h0000000, |w_size_hi, |_w_size_T_6[6:3], |_w_size_T_8[2:1], _w_size_T_10};
	always @(posedge clock) begin
		if (~reset & ~(~auto_in_ar_valid | (_r_size1_T_1[22:8] == ~_GEN_4[14:0]))) begin
			$error("Assertion failed\n    at ToTL.scala:108 assert (!in.ar.valid || r_size1 === UIntToOH1(r_size, beatCountBits)) // because aligned\n");
			$fatal;
		end
		if (~reset & ~(~auto_in_aw_valid | (_w_size1_T_1[22:8] == ~_GEN_5[14:0]))) begin
			$error("Assertion failed\n    at ToTL.scala:144 assert (!in.aw.valid || w_size1 === UIntToOH1(w_size, beatCountBits)) // because aligned\n");
			$fatal;
		end
		if (~reset & ~((~auto_in_aw_valid | (auto_in_aw_bits_len == 8'h00)) | (auto_in_aw_bits_size == 3'h3))) begin
			$error("Assertion failed\n    at ToTL.scala:145 assert (!in.aw.valid || in.aw.bits.len === 0.U || in.aw.bits.size === log2Ceil(beatBytes).U) // because aligned\n");
			$fatal;
		end
		if (~reset & ~(~winner_0 | ~winner_1)) begin
			$error("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
			$fatal;
		end
		if (~reset & ~((~_nodeOut_a_valid_T | winner_0) | winner_1)) begin
			$error("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
			$fatal;
		end
	end
	reg state_0;
	reg state_1;
	wire muxState_0 = (idle ? winner_0 : state_0);
	wire muxState_1 = (idle ? winner_1 : state_1);
	wire r_out_ready = auto_out_a_ready & (idle ? readys_readys[0] : state_0);
	assign w_out_ready = auto_out_a_ready & (idle ? readys_readys[1] : state_1);
	wire nodeOut_a_valid = (idle ? _nodeOut_a_valid_T : (state_0 & auto_in_ar_valid) | (state_1 & w_out_valid));
	wire [1:0] ok_r_bits_resp = {auto_out_d_bits_denied | auto_out_d_bits_corrupt, 1'h0};
	wire [26:0] _d_last_beats1_decode_T_1 = 27'h0000fff << auto_out_d_bits_size;
	wire [8:0] d_last_beats1 = (auto_out_d_bits_opcode[0] ? ~_d_last_beats1_decode_T_1[11:3] : 9'h000);
	reg [8:0] d_last_counter;
	wire nodeOut_d_ready = (auto_out_d_bits_opcode[0] ? _nodeIn_r_deq_q_io_enq_ready : _q_b_deq_q_io_enq_ready);
	reg [1:0] b_count_0;
	reg [1:0] b_count_1;
	reg [1:0] b_count_2;
	reg [1:0] b_count_3;
	reg [1:0] b_count_4;
	reg [1:0] b_count_5;
	reg [1:0] b_count_6;
	reg [1:0] b_count_7;
	reg [1:0] b_count_8;
	reg [1:0] b_count_9;
	reg [1:0] b_count_10;
	reg [1:0] b_count_11;
	reg [1:0] b_count_12;
	reg [1:0] b_count_13;
	reg [1:0] b_count_14;
	reg [1:0] b_count_15;
	wire [31:0] _GEN_6 = {b_count_15, b_count_14, b_count_13, b_count_12, b_count_11, b_count_10, b_count_9, b_count_8, b_count_7, b_count_6, b_count_5, b_count_4, b_count_3, b_count_2, b_count_1, b_count_0};
	wire b_allow = _GEN_6[_q_b_deq_q_io_deq_bits_id * 2+:2] != _GEN_3[_q_b_deq_q_io_deq_bits_id * 2+:2];
	wire nodeIn_b_valid = _q_b_deq_q_io_deq_valid & b_allow;
	wire [1:0] _readys_mask_T = readys_readys & readys_valid;
	wire _GEN_7 = r_out_ready & auto_in_ar_valid;
	wire _GEN_8 = nodeIn_aw_ready & auto_in_aw_valid;
	wire latch = idle & auto_out_a_ready;
	wire _GEN_9 = auto_in_b_ready & nodeIn_b_valid;
	always @(posedge clock)
		if (reset) begin
			r_count_0 <= 2'h0;
			r_count_1 <= 2'h0;
			r_count_2 <= 2'h0;
			r_count_3 <= 2'h0;
			r_count_4 <= 2'h0;
			r_count_5 <= 2'h0;
			r_count_6 <= 2'h0;
			r_count_7 <= 2'h0;
			r_count_8 <= 2'h0;
			r_count_9 <= 2'h0;
			r_count_10 <= 2'h0;
			r_count_11 <= 2'h0;
			r_count_12 <= 2'h0;
			r_count_13 <= 2'h0;
			r_count_14 <= 2'h0;
			r_count_15 <= 2'h0;
			w_count_0 <= 2'h0;
			w_count_1 <= 2'h0;
			w_count_2 <= 2'h0;
			w_count_3 <= 2'h0;
			w_count_4 <= 2'h0;
			w_count_5 <= 2'h0;
			w_count_6 <= 2'h0;
			w_count_7 <= 2'h0;
			w_count_8 <= 2'h0;
			w_count_9 <= 2'h0;
			w_count_10 <= 2'h0;
			w_count_11 <= 2'h0;
			w_count_12 <= 2'h0;
			w_count_13 <= 2'h0;
			w_count_14 <= 2'h0;
			w_count_15 <= 2'h0;
			beatsLeft <= 8'h00;
			readys_mask <= 2'h3;
			state_0 <= 1'h0;
			state_1 <= 1'h0;
			d_last_counter <= 9'h000;
			b_count_0 <= 2'h0;
			b_count_1 <= 2'h0;
			b_count_2 <= 2'h0;
			b_count_3 <= 2'h0;
			b_count_4 <= 2'h0;
			b_count_5 <= 2'h0;
			b_count_6 <= 2'h0;
			b_count_7 <= 2'h0;
			b_count_8 <= 2'h0;
			b_count_9 <= 2'h0;
			b_count_10 <= 2'h0;
			b_count_11 <= 2'h0;
			b_count_12 <= 2'h0;
			b_count_13 <= 2'h0;
			b_count_14 <= 2'h0;
			b_count_15 <= 2'h0;
		end
		else begin
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h0))
				r_count_0 <= r_count_0 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h1))
				r_count_1 <= r_count_1 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h2))
				r_count_2 <= r_count_2 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h3))
				r_count_3 <= r_count_3 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h4))
				r_count_4 <= r_count_4 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h5))
				r_count_5 <= r_count_5 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h6))
				r_count_6 <= r_count_6 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h7))
				r_count_7 <= r_count_7 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h8))
				r_count_8 <= r_count_8 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'h9))
				r_count_9 <= r_count_9 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'ha))
				r_count_10 <= r_count_10 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'hb))
				r_count_11 <= r_count_11 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'hc))
				r_count_12 <= r_count_12 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'hd))
				r_count_13 <= r_count_13 + 2'h1;
			if (_GEN_7 & (auto_in_ar_bits_id == 4'he))
				r_count_14 <= r_count_14 + 2'h1;
			if (_GEN_7 & &auto_in_ar_bits_id)
				r_count_15 <= r_count_15 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h0))
				w_count_0 <= w_count_0 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h1))
				w_count_1 <= w_count_1 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h2))
				w_count_2 <= w_count_2 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h3))
				w_count_3 <= w_count_3 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h4))
				w_count_4 <= w_count_4 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h5))
				w_count_5 <= w_count_5 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h6))
				w_count_6 <= w_count_6 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h7))
				w_count_7 <= w_count_7 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h8))
				w_count_8 <= w_count_8 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'h9))
				w_count_9 <= w_count_9 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'ha))
				w_count_10 <= w_count_10 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'hb))
				w_count_11 <= w_count_11 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'hc))
				w_count_12 <= w_count_12 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'hd))
				w_count_13 <= w_count_13 + 2'h1;
			if (_GEN_8 & (auto_in_aw_bits_id == 4'he))
				w_count_14 <= w_count_14 + 2'h1;
			if (_GEN_8 & &auto_in_aw_bits_id)
				w_count_15 <= w_count_15 + 2'h1;
			if (latch)
				beatsLeft <= (winner_1 ? auto_in_aw_bits_len : 8'h00);
			else
				beatsLeft <= beatsLeft - {7'h00, auto_out_a_ready & nodeOut_a_valid};
			if (latch & |readys_valid)
				readys_mask <= _readys_mask_T | {_readys_mask_T[0], 1'h0};
			if (idle) begin
				state_0 <= winner_0;
				state_1 <= winner_1;
			end
			if (nodeOut_d_ready & auto_out_d_valid) begin
				if (d_last_counter == 9'h000)
					d_last_counter <= d_last_beats1;
				else
					d_last_counter <= d_last_counter - 9'h001;
			end
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h0))
				b_count_0 <= b_count_0 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h1))
				b_count_1 <= b_count_1 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h2))
				b_count_2 <= b_count_2 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h3))
				b_count_3 <= b_count_3 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h4))
				b_count_4 <= b_count_4 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h5))
				b_count_5 <= b_count_5 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h6))
				b_count_6 <= b_count_6 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h7))
				b_count_7 <= b_count_7 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h8))
				b_count_8 <= b_count_8 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'h9))
				b_count_9 <= b_count_9 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'ha))
				b_count_10 <= b_count_10 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'hb))
				b_count_11 <= b_count_11 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'hc))
				b_count_12 <= b_count_12 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'hd))
				b_count_13 <= b_count_13 + 2'h1;
			if (_GEN_9 & (_q_b_deq_q_io_deq_bits_id == 4'he))
				b_count_14 <= b_count_14 + 2'h1;
			if (_GEN_9 & &_q_b_deq_q_io_deq_bits_id)
				b_count_15 <= b_count_15 + 2'h1;
		end
	wire [31:0] _RANDOM [0:3];
	Queue_54 nodeIn_r_deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_nodeIn_r_deq_q_io_enq_ready),
		.io_enq_valid(auto_out_d_valid & auto_out_d_bits_opcode[0]),
		.io_enq_bits_id(auto_out_d_bits_source[5:2]),
		.io_enq_bits_data(auto_out_d_bits_data),
		.io_enq_bits_resp(ok_r_bits_resp),
		.io_enq_bits_last((d_last_counter == 9'h001) | (d_last_beats1 == 9'h000)),
		.io_deq_ready(auto_in_r_ready),
		.io_deq_valid(auto_in_r_valid),
		.io_deq_bits_id(auto_in_r_bits_id),
		.io_deq_bits_data(auto_in_r_bits_data),
		.io_deq_bits_resp(auto_in_r_bits_resp),
		.io_deq_bits_last(auto_in_r_bits_last)
	);
	Queue_55 q_b_deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_q_b_deq_q_io_enq_ready),
		.io_enq_valid(auto_out_d_valid & ~auto_out_d_bits_opcode[0]),
		.io_enq_bits_id(auto_out_d_bits_source[5:2]),
		.io_enq_bits_resp(ok_r_bits_resp),
		.io_deq_ready(auto_in_b_ready & b_allow),
		.io_deq_valid(_q_b_deq_q_io_deq_valid),
		.io_deq_bits_id(_q_b_deq_q_io_deq_bits_id),
		.io_deq_bits_resp(auto_in_b_bits_resp)
	);
	assign auto_in_aw_ready = nodeIn_aw_ready;
	assign auto_in_w_ready = w_out_ready & auto_in_aw_valid;
	assign auto_in_b_valid = nodeIn_b_valid;
	assign auto_in_b_bits_id = _q_b_deq_q_io_deq_bits_id;
	assign auto_in_ar_ready = r_out_ready;
	assign auto_out_a_valid = nodeOut_a_valid;
	assign auto_out_a_bits_opcode = {muxState_0, 1'h0, muxState_1};
	assign auto_out_a_bits_size = (muxState_0 ? r_out_bits_a_size : 4'h0) | (muxState_1 ? w_out_bits_a_size : 4'h0);
	assign auto_out_a_bits_source = (muxState_0 ? {auto_in_ar_bits_id, _GEN_0[auto_in_ar_bits_id * 2], 1'h0} : 6'h00) | (muxState_1 ? {auto_in_aw_bits_id, _GEN_3[auto_in_aw_bits_id * 2], 1'h1} : 6'h00);
	assign auto_out_a_bits_address = (muxState_0 ? r_out_bits_a_address : 32'h00000000) | (muxState_1 ? (((w_out_bits_a_size < 4'hd) & ({auto_in_aw_bits_addr[31:14], ~auto_in_aw_bits_addr[13:12]} == 20'h00000)) | ((w_out_bits_a_size < 4'h7) & ((((((((auto_in_aw_bits_addr[31:13] == 19'h00000) | ({auto_in_aw_bits_addr[31:21], auto_in_aw_bits_addr[20:17] ^ 4'h8, auto_in_aw_bits_addr[15:12]} == 19'h00000)) | ({auto_in_aw_bits_addr[31:26], auto_in_aw_bits_addr[25:16] ^ 10'h200} == 16'h0000)) | ({auto_in_aw_bits_addr[31:26], auto_in_aw_bits_addr[25:12] ^ 14'h2010} == 20'h00000)) | ({auto_in_aw_bits_addr[31:28], auto_in_aw_bits_addr[27:16] ^ 12'h800} == 16'h0000)) | ({auto_in_aw_bits_addr[31:28], ~auto_in_aw_bits_addr[27:26]} == 6'h00)) | ({auto_in_aw_bits_addr[31:29], auto_in_aw_bits_addr[28:12] ^ 17'h10020} == 20'h00000)) | (auto_in_aw_bits_addr[31:28] == 4'h8))) ? auto_in_aw_bits_addr : {29'h00000600, auto_in_aw_bits_addr[2:0]}) : 32'h00000000);
	assign auto_out_a_bits_mask = (muxState_0 ? {r_out_bits_a_mask_acc_5 | (r_out_bits_a_mask_eq_5 & r_out_bits_a_address[0]), r_out_bits_a_mask_acc_5 | (r_out_bits_a_mask_eq_5 & ~r_out_bits_a_address[0]), r_out_bits_a_mask_acc_4 | (r_out_bits_a_mask_eq_4 & r_out_bits_a_address[0]), r_out_bits_a_mask_acc_4 | (r_out_bits_a_mask_eq_4 & ~r_out_bits_a_address[0]), r_out_bits_a_mask_acc_3 | (r_out_bits_a_mask_eq_3 & r_out_bits_a_address[0]), r_out_bits_a_mask_acc_3 | (r_out_bits_a_mask_eq_3 & ~r_out_bits_a_address[0]), r_out_bits_a_mask_acc_2 | (r_out_bits_a_mask_eq_2 & r_out_bits_a_address[0]), r_out_bits_a_mask_acc_2 | (r_out_bits_a_mask_eq_2 & ~r_out_bits_a_address[0])} : 8'h00) | (muxState_1 ? auto_in_w_bits_strb : 8'h00);
	assign auto_out_a_bits_data = (muxState_1 ? auto_in_w_bits_data : 64'h0000000000000000);
	assign auto_out_d_ready = nodeOut_d_ready;
endmodule
module Queue_56 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_real_last,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_real_last
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input io_enq_bits_real_last;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire io_deq_bits_real_last;
	reg wrap;
	reg wrap_1;
	reg maybe_full;
	wire ptr_match = wrap == wrap_1;
	wire empty = ptr_match & ~maybe_full;
	wire full = ptr_match & maybe_full;
	wire do_enq = ~full & io_enq_valid;
	wire do_deq = io_deq_ready & ~empty;
	always @(posedge clock)
		if (reset) begin
			wrap <= 1'h0;
			wrap_1 <= 1'h0;
			maybe_full <= 1'h0;
		end
		else begin
			if (do_enq)
				wrap <= wrap - 1'h1;
			if (do_deq)
				wrap_1 <= wrap_1 - 1'h1;
			if (~(do_enq == do_deq))
				maybe_full <= do_enq;
		end
	wire [31:0] _RANDOM [0:0];
	ram_2x1 ram_real_last_ext(
		.R0_addr(wrap_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(io_deq_bits_real_last),
		.W0_addr(wrap),
		.W0_en(do_enq),
		.W0_clk(clock),
		.W0_data(io_enq_bits_real_last)
	);
	assign io_enq_ready = ~full;
	assign io_deq_valid = ~empty;
endmodule
module AXI4UserYanker_1 (
	clock,
	reset,
	auto_in_aw_ready,
	auto_in_aw_valid,
	auto_in_aw_bits_id,
	auto_in_aw_bits_addr,
	auto_in_aw_bits_len,
	auto_in_aw_bits_size,
	auto_in_aw_bits_echo_real_last,
	auto_in_w_ready,
	auto_in_w_valid,
	auto_in_w_bits_data,
	auto_in_w_bits_strb,
	auto_in_w_bits_last,
	auto_in_b_ready,
	auto_in_b_valid,
	auto_in_b_bits_id,
	auto_in_b_bits_resp,
	auto_in_b_bits_echo_real_last,
	auto_in_ar_ready,
	auto_in_ar_valid,
	auto_in_ar_bits_id,
	auto_in_ar_bits_addr,
	auto_in_ar_bits_len,
	auto_in_ar_bits_size,
	auto_in_ar_bits_echo_real_last,
	auto_in_r_ready,
	auto_in_r_valid,
	auto_in_r_bits_id,
	auto_in_r_bits_data,
	auto_in_r_bits_resp,
	auto_in_r_bits_echo_real_last,
	auto_in_r_bits_last,
	auto_out_aw_ready,
	auto_out_aw_valid,
	auto_out_aw_bits_id,
	auto_out_aw_bits_addr,
	auto_out_aw_bits_len,
	auto_out_aw_bits_size,
	auto_out_w_ready,
	auto_out_w_valid,
	auto_out_w_bits_data,
	auto_out_w_bits_strb,
	auto_out_w_bits_last,
	auto_out_b_ready,
	auto_out_b_valid,
	auto_out_b_bits_id,
	auto_out_b_bits_resp,
	auto_out_ar_ready,
	auto_out_ar_valid,
	auto_out_ar_bits_id,
	auto_out_ar_bits_addr,
	auto_out_ar_bits_len,
	auto_out_ar_bits_size,
	auto_out_r_ready,
	auto_out_r_valid,
	auto_out_r_bits_id,
	auto_out_r_bits_data,
	auto_out_r_bits_resp,
	auto_out_r_bits_last
);
	input clock;
	input reset;
	output wire auto_in_aw_ready;
	input auto_in_aw_valid;
	input [3:0] auto_in_aw_bits_id;
	input [31:0] auto_in_aw_bits_addr;
	input [7:0] auto_in_aw_bits_len;
	input [2:0] auto_in_aw_bits_size;
	input auto_in_aw_bits_echo_real_last;
	output wire auto_in_w_ready;
	input auto_in_w_valid;
	input [63:0] auto_in_w_bits_data;
	input [7:0] auto_in_w_bits_strb;
	input auto_in_w_bits_last;
	input auto_in_b_ready;
	output wire auto_in_b_valid;
	output wire [3:0] auto_in_b_bits_id;
	output wire [1:0] auto_in_b_bits_resp;
	output wire auto_in_b_bits_echo_real_last;
	output wire auto_in_ar_ready;
	input auto_in_ar_valid;
	input [3:0] auto_in_ar_bits_id;
	input [31:0] auto_in_ar_bits_addr;
	input [7:0] auto_in_ar_bits_len;
	input [2:0] auto_in_ar_bits_size;
	input auto_in_ar_bits_echo_real_last;
	input auto_in_r_ready;
	output wire auto_in_r_valid;
	output wire [3:0] auto_in_r_bits_id;
	output wire [63:0] auto_in_r_bits_data;
	output wire [1:0] auto_in_r_bits_resp;
	output wire auto_in_r_bits_echo_real_last;
	output wire auto_in_r_bits_last;
	input auto_out_aw_ready;
	output wire auto_out_aw_valid;
	output wire [3:0] auto_out_aw_bits_id;
	output wire [31:0] auto_out_aw_bits_addr;
	output wire [7:0] auto_out_aw_bits_len;
	output wire [2:0] auto_out_aw_bits_size;
	input auto_out_w_ready;
	output wire auto_out_w_valid;
	output wire [63:0] auto_out_w_bits_data;
	output wire [7:0] auto_out_w_bits_strb;
	output wire auto_out_w_bits_last;
	output wire auto_out_b_ready;
	input auto_out_b_valid;
	input [3:0] auto_out_b_bits_id;
	input [1:0] auto_out_b_bits_resp;
	input auto_out_ar_ready;
	output wire auto_out_ar_valid;
	output wire [3:0] auto_out_ar_bits_id;
	output wire [31:0] auto_out_ar_bits_addr;
	output wire [7:0] auto_out_ar_bits_len;
	output wire [2:0] auto_out_ar_bits_size;
	output wire auto_out_r_ready;
	input auto_out_r_valid;
	input [3:0] auto_out_r_bits_id;
	input [63:0] auto_out_r_bits_data;
	input [1:0] auto_out_r_bits_resp;
	input auto_out_r_bits_last;
	wire _Queue_31_io_enq_ready;
	wire _Queue_31_io_deq_valid;
	wire _Queue_31_io_deq_bits_real_last;
	wire _Queue_30_io_enq_ready;
	wire _Queue_30_io_deq_valid;
	wire _Queue_30_io_deq_bits_real_last;
	wire _Queue_29_io_enq_ready;
	wire _Queue_29_io_deq_valid;
	wire _Queue_29_io_deq_bits_real_last;
	wire _Queue_28_io_enq_ready;
	wire _Queue_28_io_deq_valid;
	wire _Queue_28_io_deq_bits_real_last;
	wire _Queue_27_io_enq_ready;
	wire _Queue_27_io_deq_valid;
	wire _Queue_27_io_deq_bits_real_last;
	wire _Queue_26_io_enq_ready;
	wire _Queue_26_io_deq_valid;
	wire _Queue_26_io_deq_bits_real_last;
	wire _Queue_25_io_enq_ready;
	wire _Queue_25_io_deq_valid;
	wire _Queue_25_io_deq_bits_real_last;
	wire _Queue_24_io_enq_ready;
	wire _Queue_24_io_deq_valid;
	wire _Queue_24_io_deq_bits_real_last;
	wire _Queue_23_io_enq_ready;
	wire _Queue_23_io_deq_valid;
	wire _Queue_23_io_deq_bits_real_last;
	wire _Queue_22_io_enq_ready;
	wire _Queue_22_io_deq_valid;
	wire _Queue_22_io_deq_bits_real_last;
	wire _Queue_21_io_enq_ready;
	wire _Queue_21_io_deq_valid;
	wire _Queue_21_io_deq_bits_real_last;
	wire _Queue_20_io_enq_ready;
	wire _Queue_20_io_deq_valid;
	wire _Queue_20_io_deq_bits_real_last;
	wire _Queue_19_io_enq_ready;
	wire _Queue_19_io_deq_valid;
	wire _Queue_19_io_deq_bits_real_last;
	wire _Queue_18_io_enq_ready;
	wire _Queue_18_io_deq_valid;
	wire _Queue_18_io_deq_bits_real_last;
	wire _Queue_17_io_enq_ready;
	wire _Queue_17_io_deq_valid;
	wire _Queue_17_io_deq_bits_real_last;
	wire _Queue_16_io_enq_ready;
	wire _Queue_16_io_deq_valid;
	wire _Queue_16_io_deq_bits_real_last;
	wire _Queue_15_io_enq_ready;
	wire _Queue_15_io_deq_valid;
	wire _Queue_15_io_deq_bits_real_last;
	wire _Queue_14_io_enq_ready;
	wire _Queue_14_io_deq_valid;
	wire _Queue_14_io_deq_bits_real_last;
	wire _Queue_13_io_enq_ready;
	wire _Queue_13_io_deq_valid;
	wire _Queue_13_io_deq_bits_real_last;
	wire _Queue_12_io_enq_ready;
	wire _Queue_12_io_deq_valid;
	wire _Queue_12_io_deq_bits_real_last;
	wire _Queue_11_io_enq_ready;
	wire _Queue_11_io_deq_valid;
	wire _Queue_11_io_deq_bits_real_last;
	wire _Queue_10_io_enq_ready;
	wire _Queue_10_io_deq_valid;
	wire _Queue_10_io_deq_bits_real_last;
	wire _Queue_9_io_enq_ready;
	wire _Queue_9_io_deq_valid;
	wire _Queue_9_io_deq_bits_real_last;
	wire _Queue_8_io_enq_ready;
	wire _Queue_8_io_deq_valid;
	wire _Queue_8_io_deq_bits_real_last;
	wire _Queue_7_io_enq_ready;
	wire _Queue_7_io_deq_valid;
	wire _Queue_7_io_deq_bits_real_last;
	wire _Queue_6_io_enq_ready;
	wire _Queue_6_io_deq_valid;
	wire _Queue_6_io_deq_bits_real_last;
	wire _Queue_5_io_enq_ready;
	wire _Queue_5_io_deq_valid;
	wire _Queue_5_io_deq_bits_real_last;
	wire _Queue_4_io_enq_ready;
	wire _Queue_4_io_deq_valid;
	wire _Queue_4_io_deq_bits_real_last;
	wire _Queue_3_io_enq_ready;
	wire _Queue_3_io_deq_valid;
	wire _Queue_3_io_deq_bits_real_last;
	wire _Queue_2_io_enq_ready;
	wire _Queue_2_io_deq_valid;
	wire _Queue_2_io_deq_bits_real_last;
	wire _Queue_1_io_enq_ready;
	wire _Queue_1_io_deq_valid;
	wire _Queue_1_io_deq_bits_real_last;
	wire _Queue_io_enq_ready;
	wire _Queue_io_deq_valid;
	wire _Queue_io_deq_bits_real_last;
	wire [15:0] _GEN = {_Queue_15_io_enq_ready, _Queue_14_io_enq_ready, _Queue_13_io_enq_ready, _Queue_12_io_enq_ready, _Queue_11_io_enq_ready, _Queue_10_io_enq_ready, _Queue_9_io_enq_ready, _Queue_8_io_enq_ready, _Queue_7_io_enq_ready, _Queue_6_io_enq_ready, _Queue_5_io_enq_ready, _Queue_4_io_enq_ready, _Queue_3_io_enq_ready, _Queue_2_io_enq_ready, _Queue_1_io_enq_ready, _Queue_io_enq_ready};
	wire [15:0] _GEN_0 = {_Queue_15_io_deq_bits_real_last, _Queue_14_io_deq_bits_real_last, _Queue_13_io_deq_bits_real_last, _Queue_12_io_deq_bits_real_last, _Queue_11_io_deq_bits_real_last, _Queue_10_io_deq_bits_real_last, _Queue_9_io_deq_bits_real_last, _Queue_8_io_deq_bits_real_last, _Queue_7_io_deq_bits_real_last, _Queue_6_io_deq_bits_real_last, _Queue_5_io_deq_bits_real_last, _Queue_4_io_deq_bits_real_last, _Queue_3_io_deq_bits_real_last, _Queue_2_io_deq_bits_real_last, _Queue_1_io_deq_bits_real_last, _Queue_io_deq_bits_real_last};
	wire _GEN_1 = auto_out_r_valid & auto_in_r_ready;
	wire _GEN_2 = auto_in_ar_valid & auto_out_ar_ready;
	wire [15:0] _GEN_3 = {_Queue_31_io_enq_ready, _Queue_30_io_enq_ready, _Queue_29_io_enq_ready, _Queue_28_io_enq_ready, _Queue_27_io_enq_ready, _Queue_26_io_enq_ready, _Queue_25_io_enq_ready, _Queue_24_io_enq_ready, _Queue_23_io_enq_ready, _Queue_22_io_enq_ready, _Queue_21_io_enq_ready, _Queue_20_io_enq_ready, _Queue_19_io_enq_ready, _Queue_18_io_enq_ready, _Queue_17_io_enq_ready, _Queue_16_io_enq_ready};
	wire [15:0] _GEN_4 = {_Queue_15_io_deq_valid, _Queue_14_io_deq_valid, _Queue_13_io_deq_valid, _Queue_12_io_deq_valid, _Queue_11_io_deq_valid, _Queue_10_io_deq_valid, _Queue_9_io_deq_valid, _Queue_8_io_deq_valid, _Queue_7_io_deq_valid, _Queue_6_io_deq_valid, _Queue_5_io_deq_valid, _Queue_4_io_deq_valid, _Queue_3_io_deq_valid, _Queue_2_io_deq_valid, _Queue_1_io_deq_valid, _Queue_io_deq_valid};
	wire [15:0] _GEN_5 = {_Queue_31_io_deq_valid, _Queue_30_io_deq_valid, _Queue_29_io_deq_valid, _Queue_28_io_deq_valid, _Queue_27_io_deq_valid, _Queue_26_io_deq_valid, _Queue_25_io_deq_valid, _Queue_24_io_deq_valid, _Queue_23_io_deq_valid, _Queue_22_io_deq_valid, _Queue_21_io_deq_valid, _Queue_20_io_deq_valid, _Queue_19_io_deq_valid, _Queue_18_io_deq_valid, _Queue_17_io_deq_valid, _Queue_16_io_deq_valid};
	always @(posedge clock) begin
		if (~reset & ~(~auto_out_r_valid | _GEN_4[auto_out_r_bits_id])) begin
			$error("Assertion failed\n    at UserYanker.scala:66 assert (!out.r.valid || r_valid) // Q must be ready faster than the response\n");
			$fatal;
		end
		if (~reset & ~(~auto_out_b_valid | _GEN_5[auto_out_b_bits_id])) begin
			$error("Assertion failed\n    at UserYanker.scala:95 assert (!out.b.valid || b_valid) // Q must be ready faster than the response\n");
			$fatal;
		end
	end
	wire [15:0] _GEN_6 = {_Queue_31_io_deq_bits_real_last, _Queue_30_io_deq_bits_real_last, _Queue_29_io_deq_bits_real_last, _Queue_28_io_deq_bits_real_last, _Queue_27_io_deq_bits_real_last, _Queue_26_io_deq_bits_real_last, _Queue_25_io_deq_bits_real_last, _Queue_24_io_deq_bits_real_last, _Queue_23_io_deq_bits_real_last, _Queue_22_io_deq_bits_real_last, _Queue_21_io_deq_bits_real_last, _Queue_20_io_deq_bits_real_last, _Queue_19_io_deq_bits_real_last, _Queue_18_io_deq_bits_real_last, _Queue_17_io_deq_bits_real_last, _Queue_16_io_deq_bits_real_last};
	wire _GEN_7 = auto_out_b_valid & auto_in_b_ready;
	wire _GEN_8 = auto_in_aw_valid & auto_out_aw_ready;
	Queue_56 Queue(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h0)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h0)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_io_deq_valid),
		.io_deq_bits_real_last(_Queue_io_deq_bits_real_last)
	);
	Queue_56 Queue_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_1_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h1)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h1)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_1_io_deq_valid),
		.io_deq_bits_real_last(_Queue_1_io_deq_bits_real_last)
	);
	Queue_56 Queue_2(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_2_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h2)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h2)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_2_io_deq_valid),
		.io_deq_bits_real_last(_Queue_2_io_deq_bits_real_last)
	);
	Queue_56 Queue_3(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_3_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h3)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h3)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_3_io_deq_valid),
		.io_deq_bits_real_last(_Queue_3_io_deq_bits_real_last)
	);
	Queue_56 Queue_4(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_4_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h4)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h4)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_4_io_deq_valid),
		.io_deq_bits_real_last(_Queue_4_io_deq_bits_real_last)
	);
	Queue_56 Queue_5(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_5_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h5)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h5)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_5_io_deq_valid),
		.io_deq_bits_real_last(_Queue_5_io_deq_bits_real_last)
	);
	Queue_56 Queue_6(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_6_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h6)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h6)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_6_io_deq_valid),
		.io_deq_bits_real_last(_Queue_6_io_deq_bits_real_last)
	);
	Queue_56 Queue_7(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_7_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h7)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h7)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_7_io_deq_valid),
		.io_deq_bits_real_last(_Queue_7_io_deq_bits_real_last)
	);
	Queue_56 Queue_8(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_8_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h8)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h8)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_8_io_deq_valid),
		.io_deq_bits_real_last(_Queue_8_io_deq_bits_real_last)
	);
	Queue_56 Queue_9(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_9_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'h9)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'h9)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_9_io_deq_valid),
		.io_deq_bits_real_last(_Queue_9_io_deq_bits_real_last)
	);
	Queue_56 Queue_10(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_10_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'ha)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'ha)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_10_io_deq_valid),
		.io_deq_bits_real_last(_Queue_10_io_deq_bits_real_last)
	);
	Queue_56 Queue_11(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_11_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'hb)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'hb)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_11_io_deq_valid),
		.io_deq_bits_real_last(_Queue_11_io_deq_bits_real_last)
	);
	Queue_56 Queue_12(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_12_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'hc)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'hc)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_12_io_deq_valid),
		.io_deq_bits_real_last(_Queue_12_io_deq_bits_real_last)
	);
	Queue_56 Queue_13(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_13_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'hd)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'hd)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_13_io_deq_valid),
		.io_deq_bits_real_last(_Queue_13_io_deq_bits_real_last)
	);
	Queue_56 Queue_14(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_14_io_enq_ready),
		.io_enq_valid(_GEN_2 & (auto_in_ar_bits_id == 4'he)),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & (auto_out_r_bits_id == 4'he)) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_14_io_deq_valid),
		.io_deq_bits_real_last(_Queue_14_io_deq_bits_real_last)
	);
	Queue_56 Queue_15(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_15_io_enq_ready),
		.io_enq_valid(_GEN_2 & &auto_in_ar_bits_id),
		.io_enq_bits_real_last(auto_in_ar_bits_echo_real_last),
		.io_deq_ready((_GEN_1 & &auto_out_r_bits_id) & auto_out_r_bits_last),
		.io_deq_valid(_Queue_15_io_deq_valid),
		.io_deq_bits_real_last(_Queue_15_io_deq_bits_real_last)
	);
	Queue_56 Queue_16(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_16_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h0)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h0)),
		.io_deq_valid(_Queue_16_io_deq_valid),
		.io_deq_bits_real_last(_Queue_16_io_deq_bits_real_last)
	);
	Queue_56 Queue_17(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_17_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h1)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h1)),
		.io_deq_valid(_Queue_17_io_deq_valid),
		.io_deq_bits_real_last(_Queue_17_io_deq_bits_real_last)
	);
	Queue_56 Queue_18(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_18_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h2)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h2)),
		.io_deq_valid(_Queue_18_io_deq_valid),
		.io_deq_bits_real_last(_Queue_18_io_deq_bits_real_last)
	);
	Queue_56 Queue_19(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_19_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h3)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h3)),
		.io_deq_valid(_Queue_19_io_deq_valid),
		.io_deq_bits_real_last(_Queue_19_io_deq_bits_real_last)
	);
	Queue_56 Queue_20(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_20_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h4)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h4)),
		.io_deq_valid(_Queue_20_io_deq_valid),
		.io_deq_bits_real_last(_Queue_20_io_deq_bits_real_last)
	);
	Queue_56 Queue_21(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_21_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h5)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h5)),
		.io_deq_valid(_Queue_21_io_deq_valid),
		.io_deq_bits_real_last(_Queue_21_io_deq_bits_real_last)
	);
	Queue_56 Queue_22(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_22_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h6)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h6)),
		.io_deq_valid(_Queue_22_io_deq_valid),
		.io_deq_bits_real_last(_Queue_22_io_deq_bits_real_last)
	);
	Queue_56 Queue_23(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_23_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h7)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h7)),
		.io_deq_valid(_Queue_23_io_deq_valid),
		.io_deq_bits_real_last(_Queue_23_io_deq_bits_real_last)
	);
	Queue_56 Queue_24(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_24_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h8)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h8)),
		.io_deq_valid(_Queue_24_io_deq_valid),
		.io_deq_bits_real_last(_Queue_24_io_deq_bits_real_last)
	);
	Queue_56 Queue_25(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_25_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'h9)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'h9)),
		.io_deq_valid(_Queue_25_io_deq_valid),
		.io_deq_bits_real_last(_Queue_25_io_deq_bits_real_last)
	);
	Queue_56 Queue_26(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_26_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'ha)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'ha)),
		.io_deq_valid(_Queue_26_io_deq_valid),
		.io_deq_bits_real_last(_Queue_26_io_deq_bits_real_last)
	);
	Queue_56 Queue_27(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_27_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'hb)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'hb)),
		.io_deq_valid(_Queue_27_io_deq_valid),
		.io_deq_bits_real_last(_Queue_27_io_deq_bits_real_last)
	);
	Queue_56 Queue_28(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_28_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'hc)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'hc)),
		.io_deq_valid(_Queue_28_io_deq_valid),
		.io_deq_bits_real_last(_Queue_28_io_deq_bits_real_last)
	);
	Queue_56 Queue_29(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_29_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'hd)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'hd)),
		.io_deq_valid(_Queue_29_io_deq_valid),
		.io_deq_bits_real_last(_Queue_29_io_deq_bits_real_last)
	);
	Queue_56 Queue_30(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_30_io_enq_ready),
		.io_enq_valid(_GEN_8 & (auto_in_aw_bits_id == 4'he)),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & (auto_out_b_bits_id == 4'he)),
		.io_deq_valid(_Queue_30_io_deq_valid),
		.io_deq_bits_real_last(_Queue_30_io_deq_bits_real_last)
	);
	Queue_56 Queue_31(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(_Queue_31_io_enq_ready),
		.io_enq_valid(_GEN_8 & &auto_in_aw_bits_id),
		.io_enq_bits_real_last(auto_in_aw_bits_echo_real_last),
		.io_deq_ready(_GEN_7 & &auto_out_b_bits_id),
		.io_deq_valid(_Queue_31_io_deq_valid),
		.io_deq_bits_real_last(_Queue_31_io_deq_bits_real_last)
	);
	assign auto_in_aw_ready = auto_out_aw_ready & _GEN_3[auto_in_aw_bits_id];
	assign auto_in_w_ready = auto_out_w_ready;
	assign auto_in_b_valid = auto_out_b_valid;
	assign auto_in_b_bits_id = auto_out_b_bits_id;
	assign auto_in_b_bits_resp = auto_out_b_bits_resp;
	assign auto_in_b_bits_echo_real_last = _GEN_6[auto_out_b_bits_id];
	assign auto_in_ar_ready = auto_out_ar_ready & _GEN[auto_in_ar_bits_id];
	assign auto_in_r_valid = auto_out_r_valid;
	assign auto_in_r_bits_id = auto_out_r_bits_id;
	assign auto_in_r_bits_data = auto_out_r_bits_data;
	assign auto_in_r_bits_resp = auto_out_r_bits_resp;
	assign auto_in_r_bits_echo_real_last = _GEN_0[auto_out_r_bits_id];
	assign auto_in_r_bits_last = auto_out_r_bits_last;
	assign auto_out_aw_valid = auto_in_aw_valid & _GEN_3[auto_in_aw_bits_id];
	assign auto_out_aw_bits_id = auto_in_aw_bits_id;
	assign auto_out_aw_bits_addr = auto_in_aw_bits_addr;
	assign auto_out_aw_bits_len = auto_in_aw_bits_len;
	assign auto_out_aw_bits_size = auto_in_aw_bits_size;
	assign auto_out_w_valid = auto_in_w_valid;
	assign auto_out_w_bits_data = auto_in_w_bits_data;
	assign auto_out_w_bits_strb = auto_in_w_bits_strb;
	assign auto_out_w_bits_last = auto_in_w_bits_last;
	assign auto_out_b_ready = auto_in_b_ready;
	assign auto_out_ar_valid = auto_in_ar_valid & _GEN[auto_in_ar_bits_id];
	assign auto_out_ar_bits_id = auto_in_ar_bits_id;
	assign auto_out_ar_bits_addr = auto_in_ar_bits_addr;
	assign auto_out_ar_bits_len = auto_in_ar_bits_len;
	assign auto_out_ar_bits_size = auto_in_ar_bits_size;
	assign auto_out_r_ready = auto_in_r_ready;
endmodule
module Queue_88 (
	clock,
	reset,
	io_enq_ready,
	io_enq_valid,
	io_enq_bits_id,
	io_enq_bits_addr,
	io_enq_bits_len,
	io_enq_bits_size,
	io_enq_bits_burst,
	io_deq_ready,
	io_deq_valid,
	io_deq_bits_id,
	io_deq_bits_addr,
	io_deq_bits_len,
	io_deq_bits_size,
	io_deq_bits_burst
);
	input clock;
	input reset;
	output wire io_enq_ready;
	input io_enq_valid;
	input [3:0] io_enq_bits_id;
	input [31:0] io_enq_bits_addr;
	input [7:0] io_enq_bits_len;
	input [2:0] io_enq_bits_size;
	input [1:0] io_enq_bits_burst;
	input io_deq_ready;
	output wire io_deq_valid;
	output wire [3:0] io_deq_bits_id;
	output wire [31:0] io_deq_bits_addr;
	output wire [7:0] io_deq_bits_len;
	output wire [2:0] io_deq_bits_size;
	output wire [1:0] io_deq_bits_burst;
	reg [1:0] ram_burst;
	reg [2:0] ram_size;
	reg [7:0] ram_len;
	reg [31:0] ram_addr;
	reg [3:0] ram_id;
	reg full;
	wire _io_deq_valid_output = io_enq_valid | full;
	wire do_enq = (~(~full & io_deq_ready) & ~full) & io_enq_valid;
	always @(posedge clock) begin
		if (do_enq) begin
			ram_burst <= io_enq_bits_burst;
			ram_size <= io_enq_bits_size;
			ram_len <= io_enq_bits_len;
			ram_addr <= io_enq_bits_addr;
			ram_id <= io_enq_bits_id;
		end
		if (reset)
			full <= 1'h0;
		else if (~(do_enq == ((full & io_deq_ready) & _io_deq_valid_output)))
			full <= do_enq;
	end
	wire [31:0] _RANDOM [0:1];
	assign io_enq_ready = ~full;
	assign io_deq_valid = _io_deq_valid_output;
	assign io_deq_bits_id = (full ? ram_id : io_enq_bits_id);
	assign io_deq_bits_addr = (full ? ram_addr : io_enq_bits_addr);
	assign io_deq_bits_len = (full ? ram_len : io_enq_bits_len);
	assign io_deq_bits_size = (full ? ram_size : io_enq_bits_size);
	assign io_deq_bits_burst = (full ? ram_burst : io_enq_bits_burst);
endmodule
module AXI4Fragmenter (
	clock,
	reset,
	auto_in_aw_ready,
	auto_in_aw_valid,
	auto_in_aw_bits_id,
	auto_in_aw_bits_addr,
	auto_in_aw_bits_len,
	auto_in_aw_bits_size,
	auto_in_aw_bits_burst,
	auto_in_w_ready,
	auto_in_w_valid,
	auto_in_w_bits_data,
	auto_in_w_bits_strb,
	auto_in_w_bits_last,
	auto_in_b_ready,
	auto_in_b_valid,
	auto_in_b_bits_id,
	auto_in_b_bits_resp,
	auto_in_ar_ready,
	auto_in_ar_valid,
	auto_in_ar_bits_id,
	auto_in_ar_bits_addr,
	auto_in_ar_bits_len,
	auto_in_ar_bits_size,
	auto_in_ar_bits_burst,
	auto_in_r_ready,
	auto_in_r_valid,
	auto_in_r_bits_id,
	auto_in_r_bits_data,
	auto_in_r_bits_resp,
	auto_in_r_bits_last,
	auto_out_aw_ready,
	auto_out_aw_valid,
	auto_out_aw_bits_id,
	auto_out_aw_bits_addr,
	auto_out_aw_bits_len,
	auto_out_aw_bits_size,
	auto_out_aw_bits_echo_real_last,
	auto_out_w_ready,
	auto_out_w_valid,
	auto_out_w_bits_data,
	auto_out_w_bits_strb,
	auto_out_w_bits_last,
	auto_out_b_ready,
	auto_out_b_valid,
	auto_out_b_bits_id,
	auto_out_b_bits_resp,
	auto_out_b_bits_echo_real_last,
	auto_out_ar_ready,
	auto_out_ar_valid,
	auto_out_ar_bits_id,
	auto_out_ar_bits_addr,
	auto_out_ar_bits_len,
	auto_out_ar_bits_size,
	auto_out_ar_bits_echo_real_last,
	auto_out_r_ready,
	auto_out_r_valid,
	auto_out_r_bits_id,
	auto_out_r_bits_data,
	auto_out_r_bits_resp,
	auto_out_r_bits_echo_real_last,
	auto_out_r_bits_last
);
	input clock;
	input reset;
	output wire auto_in_aw_ready;
	input auto_in_aw_valid;
	input [3:0] auto_in_aw_bits_id;
	input [31:0] auto_in_aw_bits_addr;
	input [7:0] auto_in_aw_bits_len;
	input [2:0] auto_in_aw_bits_size;
	input [1:0] auto_in_aw_bits_burst;
	output wire auto_in_w_ready;
	input auto_in_w_valid;
	input [63:0] auto_in_w_bits_data;
	input [7:0] auto_in_w_bits_strb;
	input auto_in_w_bits_last;
	input auto_in_b_ready;
	output wire auto_in_b_valid;
	output wire [3:0] auto_in_b_bits_id;
	output wire [1:0] auto_in_b_bits_resp;
	output wire auto_in_ar_ready;
	input auto_in_ar_valid;
	input [3:0] auto_in_ar_bits_id;
	input [31:0] auto_in_ar_bits_addr;
	input [7:0] auto_in_ar_bits_len;
	input [2:0] auto_in_ar_bits_size;
	input [1:0] auto_in_ar_bits_burst;
	input auto_in_r_ready;
	output wire auto_in_r_valid;
	output wire [3:0] auto_in_r_bits_id;
	output wire [63:0] auto_in_r_bits_data;
	output wire [1:0] auto_in_r_bits_resp;
	output wire auto_in_r_bits_last;
	input auto_out_aw_ready;
	output wire auto_out_aw_valid;
	output wire [3:0] auto_out_aw_bits_id;
	output wire [31:0] auto_out_aw_bits_addr;
	output wire [7:0] auto_out_aw_bits_len;
	output wire [2:0] auto_out_aw_bits_size;
	output wire auto_out_aw_bits_echo_real_last;
	input auto_out_w_ready;
	output wire auto_out_w_valid;
	output wire [63:0] auto_out_w_bits_data;
	output wire [7:0] auto_out_w_bits_strb;
	output wire auto_out_w_bits_last;
	output wire auto_out_b_ready;
	input auto_out_b_valid;
	input [3:0] auto_out_b_bits_id;
	input [1:0] auto_out_b_bits_resp;
	input auto_out_b_bits_echo_real_last;
	input auto_out_ar_ready;
	output wire auto_out_ar_valid;
	output wire [3:0] auto_out_ar_bits_id;
	output wire [31:0] auto_out_ar_bits_addr;
	output wire [7:0] auto_out_ar_bits_len;
	output wire [2:0] auto_out_ar_bits_size;
	output wire auto_out_ar_bits_echo_real_last;
	output wire auto_out_r_ready;
	input auto_out_r_valid;
	input [3:0] auto_out_r_bits_id;
	input [63:0] auto_out_r_bits_data;
	input [1:0] auto_out_r_bits_resp;
	input auto_out_r_bits_echo_real_last;
	input auto_out_r_bits_last;
	wire nodeOut_w_valid;
	wire wbeats_ready;
	wire in_aw_ready;
	wire _in_w_deq_q_io_deq_valid;
	wire _in_w_deq_q_io_deq_bits_last;
	wire _deq_q_1_io_deq_valid;
	wire [31:0] _deq_q_1_io_deq_bits_addr;
	wire [7:0] _deq_q_1_io_deq_bits_len;
	wire [2:0] _deq_q_1_io_deq_bits_size;
	wire [1:0] _deq_q_1_io_deq_bits_burst;
	wire _deq_q_io_deq_valid;
	wire [31:0] _deq_q_io_deq_bits_addr;
	wire [7:0] _deq_q_io_deq_bits_len;
	wire [2:0] _deq_q_io_deq_bits_size;
	wire [1:0] _deq_q_io_deq_bits_burst;
	reg busy;
	reg [31:0] r_addr;
	reg [7:0] r_len;
	wire [7:0] len = (busy ? r_len : _deq_q_io_deq_bits_len);
	wire [31:0] addr = (busy ? r_addr : _deq_q_io_deq_bits_addr);
	wire [5:0] _GEN = len[6:1] | len[7:2];
	wire [4:0] _GEN_0 = _GEN[4:0] | {len[7], _GEN[5:2]};
	wire [7:0] _wipeHigh_T = ~len;
	wire [7:0] _wipeHigh_T_3 = _wipeHigh_T | {_wipeHigh_T[6:0], 1'h0};
	wire [7:0] _wipeHigh_T_6 = _wipeHigh_T_3 | {_wipeHigh_T_3[5:0], 2'h0};
	wire [7:0] _align1_T_2 = addr[10:3] | {addr[9:3], 1'h0};
	wire [7:0] _align1_T_5 = _align1_T_2 | {_align1_T_2[5:0], 2'h0};
	wire fixed = _deq_q_io_deq_bits_burst == 2'h0;
	wire [7:0] in_ar_bits_len = (fixed | (_deq_q_io_deq_bits_size != 3'h3) ? 8'h00 : (({1'h0, len[7], _GEN[5], _GEN_0[4:3], _GEN_0[2:0] | {len[7], _GEN[5], _GEN_0[4]}} | ~(_wipeHigh_T_6 | {_wipeHigh_T_6[3:0], 4'h0})) & ~(_align1_T_5 | {_align1_T_5[3:0], 4'h0})) & ({5'h00, {3 {((((((({addr[31], addr[28:27], addr[25], addr[16], addr[13]} == 6'h00) | ({addr[31], addr[28:27], ~addr[16], addr[13:12]} == 6'h00)) | ({addr[31], addr[28:27], addr[25], ~addr[16]} == 5'h00)) | ({addr[31], addr[28:27], ~addr[25], addr[16]} == 5'h00)) | ({addr[31], addr[28], ~addr[27]} == 3'h0)) | ({addr[31], addr[28], ~addr[27], addr[25], addr[16]} == 5'h00)) | ({addr[31], addr[28:27] ^ 2'h2, addr[25], addr[16], addr[13:12]} == 7'h00)) | ({~addr[31], addr[28]} == 2'h0)}}} | {8 {{addr[31], addr[28:27], addr[25], addr[16], ~addr[13:12]} == 7'h00}}));
	wire nodeOut_ar_bits_echo_real_last = in_ar_bits_len == len;
	wire [31:0] _out_bits_addr_T = ~addr;
	wire [9:0] _out_bits_addr_T_2 = 10'h007 << _deq_q_io_deq_bits_size;
	reg busy_1;
	reg [31:0] r_addr_1;
	reg [7:0] r_len_1;
	wire [7:0] len_1 = (busy_1 ? r_len_1 : _deq_q_1_io_deq_bits_len);
	wire [31:0] addr_1 = (busy_1 ? r_addr_1 : _deq_q_1_io_deq_bits_addr);
	wire [5:0] _GEN_1 = len_1[6:1] | len_1[7:2];
	wire [4:0] _GEN_2 = _GEN_1[4:0] | {len_1[7], _GEN_1[5:2]};
	wire [7:0] _wipeHigh_T_11 = ~len_1;
	wire [7:0] _wipeHigh_T_14 = _wipeHigh_T_11 | {_wipeHigh_T_11[6:0], 1'h0};
	wire [7:0] _wipeHigh_T_17 = _wipeHigh_T_14 | {_wipeHigh_T_14[5:0], 2'h0};
	wire [7:0] _align1_T_12 = addr_1[10:3] | {addr_1[9:3], 1'h0};
	wire [7:0] _align1_T_15 = _align1_T_12 | {_align1_T_12[5:0], 2'h0};
	wire fixed_1 = _deq_q_1_io_deq_bits_burst == 2'h0;
	wire [7:0] in_aw_bits_len = (fixed_1 | (_deq_q_1_io_deq_bits_size != 3'h3) ? 8'h00 : (({1'h0, len_1[7], _GEN_1[5], _GEN_2[4:3], _GEN_2[2:0] | {len_1[7], _GEN_1[5], _GEN_2[4]}} | ~(_wipeHigh_T_17 | {_wipeHigh_T_17[3:0], 4'h0})) & ~(_align1_T_15 | {_align1_T_15[3:0], 4'h0})) & ({5'h00, {3 {(((((({addr_1[31], addr_1[27], addr_1[25], addr_1[20], addr_1[13]} == 5'h00) | ({addr_1[31], addr_1[27], addr_1[25], ~addr_1[20], addr_1[13:12]} == 6'h00)) | ({addr_1[31], addr_1[27], ~addr_1[25], addr_1[20]} == 4'h0)) | ({addr_1[31], addr_1[27], ~addr_1[25], addr_1[20], addr_1[13:12]} == 6'h00)) | ({addr_1[31], ~addr_1[27]} == 2'h0)) | ({addr_1[31], ~addr_1[27], addr_1[25], addr_1[20]} == 4'h0)) | addr_1[31]}}} | {8 {{addr_1[31], addr_1[27], addr_1[25], addr_1[20], ~addr_1[13:12]} == 6'h00}}));
	wire [8:0] w_beats = {in_aw_bits_len, 1'h1} & {1'h1, ~in_aw_bits_len};
	wire nodeOut_aw_bits_echo_real_last = in_aw_bits_len == len_1;
	wire [31:0] _out_bits_addr_T_7 = ~addr_1;
	wire [9:0] _out_bits_addr_T_9 = 10'h007 << _deq_q_1_io_deq_bits_size;
	reg wbeats_latched;
	wire _in_aw_ready_T = wbeats_ready | wbeats_latched;
	wire nodeOut_aw_valid = _deq_q_1_io_deq_valid & _in_aw_ready_T;
	assign in_aw_ready = auto_out_aw_ready & _in_aw_ready_T;
	wire wbeats_valid = _deq_q_1_io_deq_valid & ~wbeats_latched;
	reg [8:0] w_counter;
	assign wbeats_ready = w_counter == 9'h000;
	wire [8:0] w_todo = (wbeats_ready ? (wbeats_valid ? w_beats : 9'h000) : w_counter);
	wire nodeOut_w_bits_last = w_todo == 9'h001;
	wire _w_counter_T = auto_out_w_ready & nodeOut_w_valid;
	assign nodeOut_w_valid = _in_w_deq_q_io_deq_valid & (~wbeats_ready | wbeats_valid);
	always @(posedge clock) begin
		if (~reset & ~(~_w_counter_T | |w_todo)) begin
			$error("Assertion failed\n    at Fragmenter.scala:177 assert (!out.w.fire || w_todo =/= 0.U) // underflow impossible\n");
			$fatal;
		end
		if (~reset & ~((~nodeOut_w_valid | ~_in_w_deq_q_io_deq_bits_last) | nodeOut_w_bits_last)) begin
			$error("Assertion failed\n    at Fragmenter.scala:186 assert (!out.w.valid || !in_w.bits.last || w_last)\n");
			$fatal;
		end
	end
	wire nodeOut_b_ready = auto_in_b_ready | ~auto_out_b_bits_echo_real_last;
	reg [1:0] error_0;
	reg [1:0] error_1;
	reg [1:0] error_2;
	reg [1:0] error_3;
	reg [1:0] error_4;
	reg [1:0] error_5;
	reg [1:0] error_6;
	reg [1:0] error_7;
	reg [1:0] error_8;
	reg [1:0] error_9;
	reg [1:0] error_10;
	reg [1:0] error_11;
	reg [1:0] error_12;
	reg [1:0] error_13;
	reg [1:0] error_14;
	reg [1:0] error_15;
	wire [31:0] _GEN_3 = {error_15, error_14, error_13, error_12, error_11, error_10, error_9, error_8, error_7, error_6, error_5, error_4, error_3, error_2, error_1, error_0};
	wire _GEN_4 = nodeOut_b_ready & auto_out_b_valid;
	wire [22:0] _wrapMask_T_1 = {7'h00, _deq_q_io_deq_bits_len, 8'hff} << _deq_q_io_deq_bits_size;
	wire [31:0] _mux_addr_T_1 = ~_deq_q_io_deq_bits_addr;
	wire [8:0] beats = {in_ar_bits_len, 1'h1} & {1'h1, ~in_ar_bits_len};
	wire [31:0] _inc_addr_T_1 = addr + {16'h0000, {7'h00, beats} << _deq_q_io_deq_bits_size};
	wire [22:0] _wrapMask_T_3 = {7'h00, _deq_q_1_io_deq_bits_len, 8'hff} << _deq_q_1_io_deq_bits_size;
	wire [31:0] _mux_addr_T_6 = ~_deq_q_1_io_deq_bits_addr;
	wire [31:0] _inc_addr_T_3 = addr_1 + {16'h0000, {7'h00, w_beats} << _deq_q_1_io_deq_bits_size};
	wire _GEN_5 = auto_out_ar_ready & _deq_q_io_deq_valid;
	wire _GEN_6 = in_aw_ready & _deq_q_1_io_deq_valid;
	always @(posedge clock) begin
		if (reset) begin
			busy <= 1'h0;
			busy_1 <= 1'h0;
			wbeats_latched <= 1'h0;
			w_counter <= 9'h000;
			error_0 <= 2'h0;
			error_1 <= 2'h0;
			error_2 <= 2'h0;
			error_3 <= 2'h0;
			error_4 <= 2'h0;
			error_5 <= 2'h0;
			error_6 <= 2'h0;
			error_7 <= 2'h0;
			error_8 <= 2'h0;
			error_9 <= 2'h0;
			error_10 <= 2'h0;
			error_11 <= 2'h0;
			error_12 <= 2'h0;
			error_13 <= 2'h0;
			error_14 <= 2'h0;
			error_15 <= 2'h0;
		end
		else begin
			if (_GEN_5)
				busy <= ~nodeOut_ar_bits_echo_real_last;
			if (_GEN_6)
				busy_1 <= ~nodeOut_aw_bits_echo_real_last;
			wbeats_latched <= ~(auto_out_aw_ready & nodeOut_aw_valid) & ((wbeats_valid & wbeats_ready) | wbeats_latched);
			w_counter <= w_todo - {8'h00, _w_counter_T};
			if ((auto_out_b_bits_id == 4'h0) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_0 <= 2'h0;
				else
					error_0 <= error_0 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h1) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_1 <= 2'h0;
				else
					error_1 <= error_1 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h2) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_2 <= 2'h0;
				else
					error_2 <= error_2 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h3) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_3 <= 2'h0;
				else
					error_3 <= error_3 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h4) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_4 <= 2'h0;
				else
					error_4 <= error_4 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h5) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_5 <= 2'h0;
				else
					error_5 <= error_5 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h6) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_6 <= 2'h0;
				else
					error_6 <= error_6 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h7) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_7 <= 2'h0;
				else
					error_7 <= error_7 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h8) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_8 <= 2'h0;
				else
					error_8 <= error_8 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'h9) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_9 <= 2'h0;
				else
					error_9 <= error_9 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'ha) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_10 <= 2'h0;
				else
					error_10 <= error_10 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'hb) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_11 <= 2'h0;
				else
					error_11 <= error_11 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'hc) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_12 <= 2'h0;
				else
					error_12 <= error_12 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'hd) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_13 <= 2'h0;
				else
					error_13 <= error_13 | auto_out_b_bits_resp;
			end
			if ((auto_out_b_bits_id == 4'he) & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_14 <= 2'h0;
				else
					error_14 <= error_14 | auto_out_b_bits_resp;
			end
			if (&auto_out_b_bits_id & _GEN_4) begin
				if (auto_out_b_bits_echo_real_last)
					error_15 <= 2'h0;
				else
					error_15 <= error_15 | auto_out_b_bits_resp;
			end
		end
		if (_GEN_5) begin
			if (fixed)
				r_addr <= _deq_q_io_deq_bits_addr;
			else if (_deq_q_io_deq_bits_burst == 2'h2)
				r_addr <= {17'h00000, _inc_addr_T_1[14:0] & _wrapMask_T_1[22:8]} | ~{_mux_addr_T_1[31:15], _mux_addr_T_1[14:0] | _wrapMask_T_1[22:8]};
			else
				r_addr <= _inc_addr_T_1;
			r_len <= len - beats[7:0];
		end
		if (_GEN_6) begin
			if (fixed_1)
				r_addr_1 <= _deq_q_1_io_deq_bits_addr;
			else if (_deq_q_1_io_deq_bits_burst == 2'h2)
				r_addr_1 <= {17'h00000, _inc_addr_T_3[14:0] & _wrapMask_T_3[22:8]} | ~{_mux_addr_T_6[31:15], _mux_addr_T_6[14:0] | _wrapMask_T_3[22:8]};
			else
				r_addr_1 <= _inc_addr_T_3;
			r_len_1 <= len_1 - w_beats[7:0];
		end
	end
	wire [31:0] _RANDOM [0:3];
	Queue_88 deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(auto_in_ar_ready),
		.io_enq_valid(auto_in_ar_valid),
		.io_enq_bits_id(auto_in_ar_bits_id),
		.io_enq_bits_addr(auto_in_ar_bits_addr),
		.io_enq_bits_len(auto_in_ar_bits_len),
		.io_enq_bits_size(auto_in_ar_bits_size),
		.io_enq_bits_burst(auto_in_ar_bits_burst),
		.io_deq_ready(auto_out_ar_ready & nodeOut_ar_bits_echo_real_last),
		.io_deq_valid(_deq_q_io_deq_valid),
		.io_deq_bits_id(auto_out_ar_bits_id),
		.io_deq_bits_addr(_deq_q_io_deq_bits_addr),
		.io_deq_bits_len(_deq_q_io_deq_bits_len),
		.io_deq_bits_size(_deq_q_io_deq_bits_size),
		.io_deq_bits_burst(_deq_q_io_deq_bits_burst)
	);
	Queue_88 deq_q_1(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(auto_in_aw_ready),
		.io_enq_valid(auto_in_aw_valid),
		.io_enq_bits_id(auto_in_aw_bits_id),
		.io_enq_bits_addr(auto_in_aw_bits_addr),
		.io_enq_bits_len(auto_in_aw_bits_len),
		.io_enq_bits_size(auto_in_aw_bits_size),
		.io_enq_bits_burst(auto_in_aw_bits_burst),
		.io_deq_ready(in_aw_ready & nodeOut_aw_bits_echo_real_last),
		.io_deq_valid(_deq_q_1_io_deq_valid),
		.io_deq_bits_id(auto_out_aw_bits_id),
		.io_deq_bits_addr(_deq_q_1_io_deq_bits_addr),
		.io_deq_bits_len(_deq_q_1_io_deq_bits_len),
		.io_deq_bits_size(_deq_q_1_io_deq_bits_size),
		.io_deq_bits_burst(_deq_q_1_io_deq_bits_burst)
	);
	Queue_37 in_w_deq_q(
		.clock(clock),
		.reset(reset),
		.io_enq_ready(auto_in_w_ready),
		.io_enq_valid(auto_in_w_valid),
		.io_enq_bits_data(auto_in_w_bits_data),
		.io_enq_bits_strb(auto_in_w_bits_strb),
		.io_enq_bits_last(auto_in_w_bits_last),
		.io_deq_ready(auto_out_w_ready & (~wbeats_ready | wbeats_valid)),
		.io_deq_valid(_in_w_deq_q_io_deq_valid),
		.io_deq_bits_data(auto_out_w_bits_data),
		.io_deq_bits_strb(auto_out_w_bits_strb),
		.io_deq_bits_last(_in_w_deq_q_io_deq_bits_last)
	);
	assign auto_in_b_valid = auto_out_b_valid & auto_out_b_bits_echo_real_last;
	assign auto_in_b_bits_id = auto_out_b_bits_id;
	assign auto_in_b_bits_resp = auto_out_b_bits_resp | _GEN_3[auto_out_b_bits_id * 2+:2];
	assign auto_in_r_valid = auto_out_r_valid;
	assign auto_in_r_bits_id = auto_out_r_bits_id;
	assign auto_in_r_bits_data = auto_out_r_bits_data;
	assign auto_in_r_bits_resp = auto_out_r_bits_resp;
	assign auto_in_r_bits_last = auto_out_r_bits_last & auto_out_r_bits_echo_real_last;
	assign auto_out_aw_valid = nodeOut_aw_valid;
	assign auto_out_aw_bits_addr = ~{_out_bits_addr_T_7[31:3], _out_bits_addr_T_7[2:0] | ~_out_bits_addr_T_9[2:0]};
	assign auto_out_aw_bits_len = in_aw_bits_len;
	assign auto_out_aw_bits_size = _deq_q_1_io_deq_bits_size;
	assign auto_out_aw_bits_echo_real_last = nodeOut_aw_bits_echo_real_last;
	assign auto_out_w_valid = nodeOut_w_valid;
	assign auto_out_w_bits_last = nodeOut_w_bits_last;
	assign auto_out_b_ready = nodeOut_b_ready;
	assign auto_out_ar_valid = _deq_q_io_deq_valid;
	assign auto_out_ar_bits_addr = ~{_out_bits_addr_T[31:3], _out_bits_addr_T[2:0] | ~_out_bits_addr_T_2[2:0]};
	assign auto_out_ar_bits_len = in_ar_bits_len;
	assign auto_out_ar_bits_size = _deq_q_io_deq_bits_size;
	assign auto_out_ar_bits_echo_real_last = nodeOut_ar_bits_echo_real_last;
	assign auto_out_r_ready = auto_in_r_ready;
endmodule
module CVA6Tile (
	clock,
	reset,
	auto_buffer_out_a_ready,
	auto_buffer_out_a_valid,
	auto_buffer_out_a_bits_opcode,
	auto_buffer_out_a_bits_param,
	auto_buffer_out_a_bits_size,
	auto_buffer_out_a_bits_source,
	auto_buffer_out_a_bits_address,
	auto_buffer_out_a_bits_mask,
	auto_buffer_out_a_bits_data,
	auto_buffer_out_a_bits_corrupt,
	auto_buffer_out_d_ready,
	auto_buffer_out_d_valid,
	auto_buffer_out_d_bits_opcode,
	auto_buffer_out_d_bits_param,
	auto_buffer_out_d_bits_size,
	auto_buffer_out_d_bits_source,
	auto_buffer_out_d_bits_sink,
	auto_buffer_out_d_bits_denied,
	auto_buffer_out_d_bits_data,
	auto_buffer_out_d_bits_corrupt,
	auto_int_local_in_3_0,
	auto_int_local_in_2_0,
	auto_int_local_in_1_0,
	auto_int_local_in_1_1,
	auto_int_local_in_0_0,
	auto_hartid_in
);
	input clock;
	input reset;
	input auto_buffer_out_a_ready;
	output wire auto_buffer_out_a_valid;
	output wire [2:0] auto_buffer_out_a_bits_opcode;
	output wire [2:0] auto_buffer_out_a_bits_param;
	output wire [3:0] auto_buffer_out_a_bits_size;
	output wire [5:0] auto_buffer_out_a_bits_source;
	output wire [31:0] auto_buffer_out_a_bits_address;
	output wire [7:0] auto_buffer_out_a_bits_mask;
	output wire [63:0] auto_buffer_out_a_bits_data;
	output wire auto_buffer_out_a_bits_corrupt;
	output wire auto_buffer_out_d_ready;
	input auto_buffer_out_d_valid;
	input [2:0] auto_buffer_out_d_bits_opcode;
	input [1:0] auto_buffer_out_d_bits_param;
	input [3:0] auto_buffer_out_d_bits_size;
	input [5:0] auto_buffer_out_d_bits_source;
	input [2:0] auto_buffer_out_d_bits_sink;
	input auto_buffer_out_d_bits_denied;
	input [63:0] auto_buffer_out_d_bits_data;
	input auto_buffer_out_d_bits_corrupt;
	input auto_int_local_in_3_0;
	input auto_int_local_in_2_0;
	input auto_int_local_in_1_0;
	input auto_int_local_in_1_1;
	input auto_int_local_in_0_0;
	input auto_hartid_in;
	wire _core_axi_req_o_aw_valid;
	wire [3:0] _core_axi_req_o_aw_bits_id;
	wire [63:0] _core_axi_req_o_aw_bits_addr;
	wire [7:0] _core_axi_req_o_aw_bits_len;
	wire [2:0] _core_axi_req_o_aw_bits_size;
	wire [1:0] _core_axi_req_o_aw_bits_burst;
	wire [3:0] _core_axi_req_o_aw_bits_region;
	wire [5:0] _core_axi_req_o_aw_bits_atop;
	wire _core_axi_req_o_aw_bits_user;
	wire _core_axi_req_o_w_valid;
	wire [63:0] _core_axi_req_o_w_bits_data;
	wire [7:0] _core_axi_req_o_w_bits_strb;
	wire _core_axi_req_o_w_bits_last;
	wire _core_axi_req_o_w_bits_user;
	wire _core_axi_req_o_ar_valid;
	wire [3:0] _core_axi_req_o_ar_bits_id;
	wire [63:0] _core_axi_req_o_ar_bits_addr;
	wire [7:0] _core_axi_req_o_ar_bits_len;
	wire [2:0] _core_axi_req_o_ar_bits_size;
	wire [1:0] _core_axi_req_o_ar_bits_burst;
	wire [3:0] _core_axi_req_o_ar_bits_region;
	wire _core_axi_req_o_ar_bits_user;
	wire _core_axi_req_o_b_ready;
	wire _core_axi_req_o_r_ready;
	wire _axi4frag_auto_in_aw_ready;
	wire _axi4frag_auto_in_w_ready;
	wire _axi4frag_auto_in_b_valid;
	wire [3:0] _axi4frag_auto_in_b_bits_id;
	wire [1:0] _axi4frag_auto_in_b_bits_resp;
	wire _axi4frag_auto_in_ar_ready;
	wire _axi4frag_auto_in_r_valid;
	wire [3:0] _axi4frag_auto_in_r_bits_id;
	wire [63:0] _axi4frag_auto_in_r_bits_data;
	wire [1:0] _axi4frag_auto_in_r_bits_resp;
	wire _axi4frag_auto_in_r_bits_last;
	wire _axi4frag_auto_out_aw_valid;
	wire [3:0] _axi4frag_auto_out_aw_bits_id;
	wire [31:0] _axi4frag_auto_out_aw_bits_addr;
	wire [7:0] _axi4frag_auto_out_aw_bits_len;
	wire [2:0] _axi4frag_auto_out_aw_bits_size;
	wire _axi4frag_auto_out_aw_bits_echo_real_last;
	wire _axi4frag_auto_out_w_valid;
	wire [63:0] _axi4frag_auto_out_w_bits_data;
	wire [7:0] _axi4frag_auto_out_w_bits_strb;
	wire _axi4frag_auto_out_w_bits_last;
	wire _axi4frag_auto_out_b_ready;
	wire _axi4frag_auto_out_ar_valid;
	wire [3:0] _axi4frag_auto_out_ar_bits_id;
	wire [31:0] _axi4frag_auto_out_ar_bits_addr;
	wire [7:0] _axi4frag_auto_out_ar_bits_len;
	wire [2:0] _axi4frag_auto_out_ar_bits_size;
	wire _axi4frag_auto_out_ar_bits_echo_real_last;
	wire _axi4frag_auto_out_r_ready;
	wire _axi4yank_auto_in_aw_ready;
	wire _axi4yank_auto_in_w_ready;
	wire _axi4yank_auto_in_b_valid;
	wire [3:0] _axi4yank_auto_in_b_bits_id;
	wire [1:0] _axi4yank_auto_in_b_bits_resp;
	wire _axi4yank_auto_in_b_bits_echo_real_last;
	wire _axi4yank_auto_in_ar_ready;
	wire _axi4yank_auto_in_r_valid;
	wire [3:0] _axi4yank_auto_in_r_bits_id;
	wire [63:0] _axi4yank_auto_in_r_bits_data;
	wire [1:0] _axi4yank_auto_in_r_bits_resp;
	wire _axi4yank_auto_in_r_bits_echo_real_last;
	wire _axi4yank_auto_in_r_bits_last;
	wire _axi4yank_auto_out_aw_valid;
	wire [3:0] _axi4yank_auto_out_aw_bits_id;
	wire [31:0] _axi4yank_auto_out_aw_bits_addr;
	wire [7:0] _axi4yank_auto_out_aw_bits_len;
	wire [2:0] _axi4yank_auto_out_aw_bits_size;
	wire _axi4yank_auto_out_w_valid;
	wire [63:0] _axi4yank_auto_out_w_bits_data;
	wire [7:0] _axi4yank_auto_out_w_bits_strb;
	wire _axi4yank_auto_out_w_bits_last;
	wire _axi4yank_auto_out_b_ready;
	wire _axi4yank_auto_out_ar_valid;
	wire [3:0] _axi4yank_auto_out_ar_bits_id;
	wire [31:0] _axi4yank_auto_out_ar_bits_addr;
	wire [7:0] _axi4yank_auto_out_ar_bits_len;
	wire [2:0] _axi4yank_auto_out_ar_bits_size;
	wire _axi4yank_auto_out_r_ready;
	wire _axi42tl_auto_in_aw_ready;
	wire _axi42tl_auto_in_w_ready;
	wire _axi42tl_auto_in_b_valid;
	wire [3:0] _axi42tl_auto_in_b_bits_id;
	wire [1:0] _axi42tl_auto_in_b_bits_resp;
	wire _axi42tl_auto_in_ar_ready;
	wire _axi42tl_auto_in_r_valid;
	wire [3:0] _axi42tl_auto_in_r_bits_id;
	wire [63:0] _axi42tl_auto_in_r_bits_data;
	wire [1:0] _axi42tl_auto_in_r_bits_resp;
	wire _axi42tl_auto_in_r_bits_last;
	wire _axi42tl_auto_out_a_valid;
	wire [2:0] _axi42tl_auto_out_a_bits_opcode;
	wire [3:0] _axi42tl_auto_out_a_bits_size;
	wire [5:0] _axi42tl_auto_out_a_bits_source;
	wire [31:0] _axi42tl_auto_out_a_bits_address;
	wire [7:0] _axi42tl_auto_out_a_bits_mask;
	wire [63:0] _axi42tl_auto_out_a_bits_data;
	wire _axi42tl_auto_out_d_ready;
	wire _fixer_auto_in_a_ready;
	wire _fixer_auto_in_d_valid;
	wire [2:0] _fixer_auto_in_d_bits_opcode;
	wire [3:0] _fixer_auto_in_d_bits_size;
	wire [5:0] _fixer_auto_in_d_bits_source;
	wire _fixer_auto_in_d_bits_denied;
	wire [63:0] _fixer_auto_in_d_bits_data;
	wire _fixer_auto_in_d_bits_corrupt;
	wire _fixer_auto_out_a_valid;
	wire [2:0] _fixer_auto_out_a_bits_opcode;
	wire [3:0] _fixer_auto_out_a_bits_size;
	wire [5:0] _fixer_auto_out_a_bits_source;
	wire [31:0] _fixer_auto_out_a_bits_address;
	wire [7:0] _fixer_auto_out_a_bits_mask;
	wire [63:0] _fixer_auto_out_a_bits_data;
	wire _fixer_auto_out_d_ready;
	wire _buffer_auto_in_a_ready;
	wire _buffer_auto_in_d_valid;
	wire [2:0] _buffer_auto_in_d_bits_opcode;
	wire [1:0] _buffer_auto_in_d_bits_param;
	wire [3:0] _buffer_auto_in_d_bits_size;
	wire [5:0] _buffer_auto_in_d_bits_source;
	wire [2:0] _buffer_auto_in_d_bits_sink;
	wire _buffer_auto_in_d_bits_denied;
	wire [63:0] _buffer_auto_in_d_bits_data;
	wire _buffer_auto_in_d_bits_corrupt;
	wire _intXbar_auto_int_out_0;
	wire _intXbar_auto_int_out_1;
	wire _intXbar_auto_int_out_2;
	wire _intXbar_auto_int_out_3;
	wire _intXbar_auto_int_out_4;
	always @(posedge clock) begin
		if (~reset & |_core_axi_req_o_aw_bits_region) begin
			$error("Assertion failed\n    at CVA6Tile.scala:306 assert(core.io.axi_req_o_aw_bits_region === 0.U)\n");
			$fatal;
		end
		if (~reset & |_core_axi_req_o_aw_bits_atop) begin
			$error("Assertion failed\n    at CVA6Tile.scala:307 assert(core.io.axi_req_o_aw_bits_atop === 0.U)\n");
			$fatal;
		end
		if (~reset & _core_axi_req_o_aw_bits_user) begin
			$error("Assertion failed\n    at CVA6Tile.scala:308 assert(core.io.axi_req_o_aw_bits_user === 0.U)\n");
			$fatal;
		end
		if (~reset & _core_axi_req_o_w_bits_user) begin
			$error("Assertion failed\n    at CVA6Tile.scala:316 assert(core.io.axi_req_o_w_bits_user === 0.U)\n");
			$fatal;
		end
		if (~reset & |_core_axi_req_o_ar_bits_region) begin
			$error("Assertion failed\n    at CVA6Tile.scala:336 assert(core.io.axi_req_o_ar_bits_region === 0.U)\n");
			$fatal;
		end
		if (~reset & _core_axi_req_o_ar_bits_user) begin
			$error("Assertion failed\n    at CVA6Tile.scala:337 assert(core.io.axi_req_o_ar_bits_user === 0.U)\n");
			$fatal;
		end
	end
	IntXbar_1 intXbar(
		.auto_int_in_3_0(auto_int_local_in_3_0),
		.auto_int_in_2_0(auto_int_local_in_2_0),
		.auto_int_in_1_0(auto_int_local_in_1_0),
		.auto_int_in_1_1(auto_int_local_in_1_1),
		.auto_int_in_0_0(auto_int_local_in_0_0),
		.auto_int_out_0(_intXbar_auto_int_out_0),
		.auto_int_out_1(_intXbar_auto_int_out_1),
		.auto_int_out_2(_intXbar_auto_int_out_2),
		.auto_int_out_3(_intXbar_auto_int_out_3),
		.auto_int_out_4(_intXbar_auto_int_out_4)
	);
	TLBuffer_14 buffer(
		.clock(clock),
		.reset(reset),
		.auto_in_a_ready(_buffer_auto_in_a_ready),
		.auto_in_a_valid(_fixer_auto_out_a_valid),
		.auto_in_a_bits_opcode(_fixer_auto_out_a_bits_opcode),
		.auto_in_a_bits_size(_fixer_auto_out_a_bits_size),
		.auto_in_a_bits_source(_fixer_auto_out_a_bits_source),
		.auto_in_a_bits_address(_fixer_auto_out_a_bits_address),
		.auto_in_a_bits_mask(_fixer_auto_out_a_bits_mask),
		.auto_in_a_bits_data(_fixer_auto_out_a_bits_data),
		.auto_in_d_ready(_fixer_auto_out_d_ready),
		.auto_in_d_valid(_buffer_auto_in_d_valid),
		.auto_in_d_bits_opcode(_buffer_auto_in_d_bits_opcode),
		.auto_in_d_bits_param(_buffer_auto_in_d_bits_param),
		.auto_in_d_bits_size(_buffer_auto_in_d_bits_size),
		.auto_in_d_bits_source(_buffer_auto_in_d_bits_source),
		.auto_in_d_bits_sink(_buffer_auto_in_d_bits_sink),
		.auto_in_d_bits_denied(_buffer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(_buffer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(auto_buffer_out_a_ready),
		.auto_out_a_valid(auto_buffer_out_a_valid),
		.auto_out_a_bits_opcode(auto_buffer_out_a_bits_opcode),
		.auto_out_a_bits_param(auto_buffer_out_a_bits_param),
		.auto_out_a_bits_size(auto_buffer_out_a_bits_size),
		.auto_out_a_bits_source(auto_buffer_out_a_bits_source),
		.auto_out_a_bits_address(auto_buffer_out_a_bits_address),
		.auto_out_a_bits_mask(auto_buffer_out_a_bits_mask),
		.auto_out_a_bits_data(auto_buffer_out_a_bits_data),
		.auto_out_a_bits_corrupt(auto_buffer_out_a_bits_corrupt),
		.auto_out_d_ready(auto_buffer_out_d_ready),
		.auto_out_d_valid(auto_buffer_out_d_valid),
		.auto_out_d_bits_opcode(auto_buffer_out_d_bits_opcode),
		.auto_out_d_bits_param(auto_buffer_out_d_bits_param),
		.auto_out_d_bits_size(auto_buffer_out_d_bits_size),
		.auto_out_d_bits_source(auto_buffer_out_d_bits_source),
		.auto_out_d_bits_sink(auto_buffer_out_d_bits_sink),
		.auto_out_d_bits_denied(auto_buffer_out_d_bits_denied),
		.auto_out_d_bits_data(auto_buffer_out_d_bits_data),
		.auto_out_d_bits_corrupt(auto_buffer_out_d_bits_corrupt)
	);
	TLFIFOFixer_5 fixer(
		.clock(clock),
		.reset(reset),
		.auto_in_a_ready(_fixer_auto_in_a_ready),
		.auto_in_a_valid(_axi42tl_auto_out_a_valid),
		.auto_in_a_bits_opcode(_axi42tl_auto_out_a_bits_opcode),
		.auto_in_a_bits_size(_axi42tl_auto_out_a_bits_size),
		.auto_in_a_bits_source(_axi42tl_auto_out_a_bits_source),
		.auto_in_a_bits_address(_axi42tl_auto_out_a_bits_address),
		.auto_in_a_bits_mask(_axi42tl_auto_out_a_bits_mask),
		.auto_in_a_bits_data(_axi42tl_auto_out_a_bits_data),
		.auto_in_d_ready(_axi42tl_auto_out_d_ready),
		.auto_in_d_valid(_fixer_auto_in_d_valid),
		.auto_in_d_bits_opcode(_fixer_auto_in_d_bits_opcode),
		.auto_in_d_bits_size(_fixer_auto_in_d_bits_size),
		.auto_in_d_bits_source(_fixer_auto_in_d_bits_source),
		.auto_in_d_bits_denied(_fixer_auto_in_d_bits_denied),
		.auto_in_d_bits_data(_fixer_auto_in_d_bits_data),
		.auto_in_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt),
		.auto_out_a_ready(_buffer_auto_in_a_ready),
		.auto_out_a_valid(_fixer_auto_out_a_valid),
		.auto_out_a_bits_opcode(_fixer_auto_out_a_bits_opcode),
		.auto_out_a_bits_size(_fixer_auto_out_a_bits_size),
		.auto_out_a_bits_source(_fixer_auto_out_a_bits_source),
		.auto_out_a_bits_address(_fixer_auto_out_a_bits_address),
		.auto_out_a_bits_mask(_fixer_auto_out_a_bits_mask),
		.auto_out_a_bits_data(_fixer_auto_out_a_bits_data),
		.auto_out_d_ready(_fixer_auto_out_d_ready),
		.auto_out_d_valid(_buffer_auto_in_d_valid),
		.auto_out_d_bits_opcode(_buffer_auto_in_d_bits_opcode),
		.auto_out_d_bits_param(_buffer_auto_in_d_bits_param),
		.auto_out_d_bits_size(_buffer_auto_in_d_bits_size),
		.auto_out_d_bits_source(_buffer_auto_in_d_bits_source),
		.auto_out_d_bits_sink(_buffer_auto_in_d_bits_sink),
		.auto_out_d_bits_denied(_buffer_auto_in_d_bits_denied),
		.auto_out_d_bits_data(_buffer_auto_in_d_bits_data),
		.auto_out_d_bits_corrupt(_buffer_auto_in_d_bits_corrupt)
	);
	AXI4ToTL axi42tl(
		.clock(clock),
		.reset(reset),
		.auto_in_aw_ready(_axi42tl_auto_in_aw_ready),
		.auto_in_aw_valid(_axi4yank_auto_out_aw_valid),
		.auto_in_aw_bits_id(_axi4yank_auto_out_aw_bits_id),
		.auto_in_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),
		.auto_in_aw_bits_len(_axi4yank_auto_out_aw_bits_len),
		.auto_in_aw_bits_size(_axi4yank_auto_out_aw_bits_size),
		.auto_in_w_ready(_axi42tl_auto_in_w_ready),
		.auto_in_w_valid(_axi4yank_auto_out_w_valid),
		.auto_in_w_bits_data(_axi4yank_auto_out_w_bits_data),
		.auto_in_w_bits_strb(_axi4yank_auto_out_w_bits_strb),
		.auto_in_w_bits_last(_axi4yank_auto_out_w_bits_last),
		.auto_in_b_ready(_axi4yank_auto_out_b_ready),
		.auto_in_b_valid(_axi42tl_auto_in_b_valid),
		.auto_in_b_bits_id(_axi42tl_auto_in_b_bits_id),
		.auto_in_b_bits_resp(_axi42tl_auto_in_b_bits_resp),
		.auto_in_ar_ready(_axi42tl_auto_in_ar_ready),
		.auto_in_ar_valid(_axi4yank_auto_out_ar_valid),
		.auto_in_ar_bits_id(_axi4yank_auto_out_ar_bits_id),
		.auto_in_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),
		.auto_in_ar_bits_len(_axi4yank_auto_out_ar_bits_len),
		.auto_in_ar_bits_size(_axi4yank_auto_out_ar_bits_size),
		.auto_in_r_ready(_axi4yank_auto_out_r_ready),
		.auto_in_r_valid(_axi42tl_auto_in_r_valid),
		.auto_in_r_bits_id(_axi42tl_auto_in_r_bits_id),
		.auto_in_r_bits_data(_axi42tl_auto_in_r_bits_data),
		.auto_in_r_bits_resp(_axi42tl_auto_in_r_bits_resp),
		.auto_in_r_bits_last(_axi42tl_auto_in_r_bits_last),
		.auto_out_a_ready(_fixer_auto_in_a_ready),
		.auto_out_a_valid(_axi42tl_auto_out_a_valid),
		.auto_out_a_bits_opcode(_axi42tl_auto_out_a_bits_opcode),
		.auto_out_a_bits_size(_axi42tl_auto_out_a_bits_size),
		.auto_out_a_bits_source(_axi42tl_auto_out_a_bits_source),
		.auto_out_a_bits_address(_axi42tl_auto_out_a_bits_address),
		.auto_out_a_bits_mask(_axi42tl_auto_out_a_bits_mask),
		.auto_out_a_bits_data(_axi42tl_auto_out_a_bits_data),
		.auto_out_d_ready(_axi42tl_auto_out_d_ready),
		.auto_out_d_valid(_fixer_auto_in_d_valid),
		.auto_out_d_bits_opcode(_fixer_auto_in_d_bits_opcode),
		.auto_out_d_bits_size(_fixer_auto_in_d_bits_size),
		.auto_out_d_bits_source(_fixer_auto_in_d_bits_source),
		.auto_out_d_bits_denied(_fixer_auto_in_d_bits_denied),
		.auto_out_d_bits_data(_fixer_auto_in_d_bits_data),
		.auto_out_d_bits_corrupt(_fixer_auto_in_d_bits_corrupt)
	);
	AXI4UserYanker_1 axi4yank(
		.clock(clock),
		.reset(reset),
		.auto_in_aw_ready(_axi4yank_auto_in_aw_ready),
		.auto_in_aw_valid(_axi4frag_auto_out_aw_valid),
		.auto_in_aw_bits_id(_axi4frag_auto_out_aw_bits_id),
		.auto_in_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),
		.auto_in_aw_bits_len(_axi4frag_auto_out_aw_bits_len),
		.auto_in_aw_bits_size(_axi4frag_auto_out_aw_bits_size),
		.auto_in_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),
		.auto_in_w_ready(_axi4yank_auto_in_w_ready),
		.auto_in_w_valid(_axi4frag_auto_out_w_valid),
		.auto_in_w_bits_data(_axi4frag_auto_out_w_bits_data),
		.auto_in_w_bits_strb(_axi4frag_auto_out_w_bits_strb),
		.auto_in_w_bits_last(_axi4frag_auto_out_w_bits_last),
		.auto_in_b_ready(_axi4frag_auto_out_b_ready),
		.auto_in_b_valid(_axi4yank_auto_in_b_valid),
		.auto_in_b_bits_id(_axi4yank_auto_in_b_bits_id),
		.auto_in_b_bits_resp(_axi4yank_auto_in_b_bits_resp),
		.auto_in_b_bits_echo_real_last(_axi4yank_auto_in_b_bits_echo_real_last),
		.auto_in_ar_ready(_axi4yank_auto_in_ar_ready),
		.auto_in_ar_valid(_axi4frag_auto_out_ar_valid),
		.auto_in_ar_bits_id(_axi4frag_auto_out_ar_bits_id),
		.auto_in_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),
		.auto_in_ar_bits_len(_axi4frag_auto_out_ar_bits_len),
		.auto_in_ar_bits_size(_axi4frag_auto_out_ar_bits_size),
		.auto_in_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),
		.auto_in_r_ready(_axi4frag_auto_out_r_ready),
		.auto_in_r_valid(_axi4yank_auto_in_r_valid),
		.auto_in_r_bits_id(_axi4yank_auto_in_r_bits_id),
		.auto_in_r_bits_data(_axi4yank_auto_in_r_bits_data),
		.auto_in_r_bits_resp(_axi4yank_auto_in_r_bits_resp),
		.auto_in_r_bits_echo_real_last(_axi4yank_auto_in_r_bits_echo_real_last),
		.auto_in_r_bits_last(_axi4yank_auto_in_r_bits_last),
		.auto_out_aw_ready(_axi42tl_auto_in_aw_ready),
		.auto_out_aw_valid(_axi4yank_auto_out_aw_valid),
		.auto_out_aw_bits_id(_axi4yank_auto_out_aw_bits_id),
		.auto_out_aw_bits_addr(_axi4yank_auto_out_aw_bits_addr),
		.auto_out_aw_bits_len(_axi4yank_auto_out_aw_bits_len),
		.auto_out_aw_bits_size(_axi4yank_auto_out_aw_bits_size),
		.auto_out_w_ready(_axi42tl_auto_in_w_ready),
		.auto_out_w_valid(_axi4yank_auto_out_w_valid),
		.auto_out_w_bits_data(_axi4yank_auto_out_w_bits_data),
		.auto_out_w_bits_strb(_axi4yank_auto_out_w_bits_strb),
		.auto_out_w_bits_last(_axi4yank_auto_out_w_bits_last),
		.auto_out_b_ready(_axi4yank_auto_out_b_ready),
		.auto_out_b_valid(_axi42tl_auto_in_b_valid),
		.auto_out_b_bits_id(_axi42tl_auto_in_b_bits_id),
		.auto_out_b_bits_resp(_axi42tl_auto_in_b_bits_resp),
		.auto_out_ar_ready(_axi42tl_auto_in_ar_ready),
		.auto_out_ar_valid(_axi4yank_auto_out_ar_valid),
		.auto_out_ar_bits_id(_axi4yank_auto_out_ar_bits_id),
		.auto_out_ar_bits_addr(_axi4yank_auto_out_ar_bits_addr),
		.auto_out_ar_bits_len(_axi4yank_auto_out_ar_bits_len),
		.auto_out_ar_bits_size(_axi4yank_auto_out_ar_bits_size),
		.auto_out_r_ready(_axi4yank_auto_out_r_ready),
		.auto_out_r_valid(_axi42tl_auto_in_r_valid),
		.auto_out_r_bits_id(_axi42tl_auto_in_r_bits_id),
		.auto_out_r_bits_data(_axi42tl_auto_in_r_bits_data),
		.auto_out_r_bits_resp(_axi42tl_auto_in_r_bits_resp),
		.auto_out_r_bits_last(_axi42tl_auto_in_r_bits_last)
	);
	AXI4Fragmenter axi4frag(
		.clock(clock),
		.reset(reset),
		.auto_in_aw_ready(_axi4frag_auto_in_aw_ready),
		.auto_in_aw_valid(_core_axi_req_o_aw_valid),
		.auto_in_aw_bits_id(_core_axi_req_o_aw_bits_id),
		.auto_in_aw_bits_addr(_core_axi_req_o_aw_bits_addr[31:0]),
		.auto_in_aw_bits_len(_core_axi_req_o_aw_bits_len),
		.auto_in_aw_bits_size(_core_axi_req_o_aw_bits_size),
		.auto_in_aw_bits_burst(_core_axi_req_o_aw_bits_burst),
		.auto_in_w_ready(_axi4frag_auto_in_w_ready),
		.auto_in_w_valid(_core_axi_req_o_w_valid),
		.auto_in_w_bits_data(_core_axi_req_o_w_bits_data),
		.auto_in_w_bits_strb(_core_axi_req_o_w_bits_strb),
		.auto_in_w_bits_last(_core_axi_req_o_w_bits_last),
		.auto_in_b_ready(_core_axi_req_o_b_ready),
		.auto_in_b_valid(_axi4frag_auto_in_b_valid),
		.auto_in_b_bits_id(_axi4frag_auto_in_b_bits_id),
		.auto_in_b_bits_resp(_axi4frag_auto_in_b_bits_resp),
		.auto_in_ar_ready(_axi4frag_auto_in_ar_ready),
		.auto_in_ar_valid(_core_axi_req_o_ar_valid),
		.auto_in_ar_bits_id(_core_axi_req_o_ar_bits_id),
		.auto_in_ar_bits_addr(_core_axi_req_o_ar_bits_addr[31:0]),
		.auto_in_ar_bits_len(_core_axi_req_o_ar_bits_len),
		.auto_in_ar_bits_size(_core_axi_req_o_ar_bits_size),
		.auto_in_ar_bits_burst(_core_axi_req_o_ar_bits_burst),
		.auto_in_r_ready(_core_axi_req_o_r_ready),
		.auto_in_r_valid(_axi4frag_auto_in_r_valid),
		.auto_in_r_bits_id(_axi4frag_auto_in_r_bits_id),
		.auto_in_r_bits_data(_axi4frag_auto_in_r_bits_data),
		.auto_in_r_bits_resp(_axi4frag_auto_in_r_bits_resp),
		.auto_in_r_bits_last(_axi4frag_auto_in_r_bits_last),
		.auto_out_aw_ready(_axi4yank_auto_in_aw_ready),
		.auto_out_aw_valid(_axi4frag_auto_out_aw_valid),
		.auto_out_aw_bits_id(_axi4frag_auto_out_aw_bits_id),
		.auto_out_aw_bits_addr(_axi4frag_auto_out_aw_bits_addr),
		.auto_out_aw_bits_len(_axi4frag_auto_out_aw_bits_len),
		.auto_out_aw_bits_size(_axi4frag_auto_out_aw_bits_size),
		.auto_out_aw_bits_echo_real_last(_axi4frag_auto_out_aw_bits_echo_real_last),
		.auto_out_w_ready(_axi4yank_auto_in_w_ready),
		.auto_out_w_valid(_axi4frag_auto_out_w_valid),
		.auto_out_w_bits_data(_axi4frag_auto_out_w_bits_data),
		.auto_out_w_bits_strb(_axi4frag_auto_out_w_bits_strb),
		.auto_out_w_bits_last(_axi4frag_auto_out_w_bits_last),
		.auto_out_b_ready(_axi4frag_auto_out_b_ready),
		.auto_out_b_valid(_axi4yank_auto_in_b_valid),
		.auto_out_b_bits_id(_axi4yank_auto_in_b_bits_id),
		.auto_out_b_bits_resp(_axi4yank_auto_in_b_bits_resp),
		.auto_out_b_bits_echo_real_last(_axi4yank_auto_in_b_bits_echo_real_last),
		.auto_out_ar_ready(_axi4yank_auto_in_ar_ready),
		.auto_out_ar_valid(_axi4frag_auto_out_ar_valid),
		.auto_out_ar_bits_id(_axi4frag_auto_out_ar_bits_id),
		.auto_out_ar_bits_addr(_axi4frag_auto_out_ar_bits_addr),
		.auto_out_ar_bits_len(_axi4frag_auto_out_ar_bits_len),
		.auto_out_ar_bits_size(_axi4frag_auto_out_ar_bits_size),
		.auto_out_ar_bits_echo_real_last(_axi4frag_auto_out_ar_bits_echo_real_last),
		.auto_out_r_ready(_axi4frag_auto_out_r_ready),
		.auto_out_r_valid(_axi4yank_auto_in_r_valid),
		.auto_out_r_bits_id(_axi4yank_auto_in_r_bits_id),
		.auto_out_r_bits_data(_axi4yank_auto_in_r_bits_data),
		.auto_out_r_bits_resp(_axi4yank_auto_in_r_bits_resp),
		.auto_out_r_bits_echo_real_last(_axi4yank_auto_in_r_bits_echo_real_last),
		.auto_out_r_bits_last(_axi4yank_auto_in_r_bits_last)
	);
	CVA6CoreBlackbox #(
		.AXI_ADDRESS_WIDTH(64),
		.AXI_DATA_WIDTH(64),
		.AXI_ID_WIDTH(4),
		.AXI_USER_WIDTH(1),
		.BHT_ENTRIES(16),
		.BTB_ENTRIES(16),
		.CACHE_REG_BASE_0(40'd2147487872),
		.CACHE_REG_BASE_1(40'd2147483648),
		.CACHE_REG_BASE_2(0),
		.CACHE_REG_BASE_3(0),
		.CACHE_REG_BASE_4(0),
		.CACHE_REG_CNT(5),
		.CACHE_REG_SZ_0(268431232),
		.CACHE_REG_SZ_1(4096),
		.CACHE_REG_SZ_2(0),
		.CACHE_REG_SZ_3(0),
		.CACHE_REG_SZ_4(0),
		.DEBUG_BASE(0),
		.EXEC_REG_BASE_0(40'd2147483648),
		.EXEC_REG_BASE_1(65536),
		.EXEC_REG_BASE_2(0),
		.EXEC_REG_BASE_3(0),
		.EXEC_REG_BASE_4(0),
		.EXEC_REG_CNT(5),
		.EXEC_REG_SZ_0(268435456),
		.EXEC_REG_SZ_1(65536),
		.EXEC_REG_SZ_2(4096),
		.EXEC_REG_SZ_3(0),
		.EXEC_REG_SZ_4(0),
		.PMP_ENTRIES(4),
		.RAS_ENTRIES(4),
		.TRACEPORT_SZ(368),
		.XLEN(64)
	) core(
		.clk_i(clock),
		.rst_ni(~reset),
		.boot_addr_i(64'h0000000000010000),
		.hart_id_i({63'h0000000000000000, auto_hartid_in}),
		.irq_i({_intXbar_auto_int_out_4, _intXbar_auto_int_out_3}),
		.ipi_i(_intXbar_auto_int_out_1),
		.time_irq_i(_intXbar_auto_int_out_2),
		.debug_req_i(_intXbar_auto_int_out_0),
		.trace_o(),
		.axi_resp_i_aw_ready(_axi4frag_auto_in_aw_ready),
		.axi_req_o_aw_valid(_core_axi_req_o_aw_valid),
		.axi_req_o_aw_bits_id(_core_axi_req_o_aw_bits_id),
		.axi_req_o_aw_bits_addr(_core_axi_req_o_aw_bits_addr),
		.axi_req_o_aw_bits_len(_core_axi_req_o_aw_bits_len),
		.axi_req_o_aw_bits_size(_core_axi_req_o_aw_bits_size),
		.axi_req_o_aw_bits_burst(_core_axi_req_o_aw_bits_burst),
		.axi_req_o_aw_bits_lock(),
		.axi_req_o_aw_bits_cache(),
		.axi_req_o_aw_bits_prot(),
		.axi_req_o_aw_bits_qos(),
		.axi_req_o_aw_bits_region(_core_axi_req_o_aw_bits_region),
		.axi_req_o_aw_bits_atop(_core_axi_req_o_aw_bits_atop),
		.axi_req_o_aw_bits_user(_core_axi_req_o_aw_bits_user),
		.axi_resp_i_w_ready(_axi4frag_auto_in_w_ready),
		.axi_req_o_w_valid(_core_axi_req_o_w_valid),
		.axi_req_o_w_bits_data(_core_axi_req_o_w_bits_data),
		.axi_req_o_w_bits_strb(_core_axi_req_o_w_bits_strb),
		.axi_req_o_w_bits_last(_core_axi_req_o_w_bits_last),
		.axi_req_o_w_bits_user(_core_axi_req_o_w_bits_user),
		.axi_resp_i_ar_ready(_axi4frag_auto_in_ar_ready),
		.axi_req_o_ar_valid(_core_axi_req_o_ar_valid),
		.axi_req_o_ar_bits_id(_core_axi_req_o_ar_bits_id),
		.axi_req_o_ar_bits_addr(_core_axi_req_o_ar_bits_addr),
		.axi_req_o_ar_bits_len(_core_axi_req_o_ar_bits_len),
		.axi_req_o_ar_bits_size(_core_axi_req_o_ar_bits_size),
		.axi_req_o_ar_bits_burst(_core_axi_req_o_ar_bits_burst),
		.axi_req_o_ar_bits_lock(),
		.axi_req_o_ar_bits_cache(),
		.axi_req_o_ar_bits_prot(),
		.axi_req_o_ar_bits_qos(),
		.axi_req_o_ar_bits_region(_core_axi_req_o_ar_bits_region),
		.axi_req_o_ar_bits_user(_core_axi_req_o_ar_bits_user),
		.axi_req_o_b_ready(_core_axi_req_o_b_ready),
		.axi_resp_i_b_valid(_axi4frag_auto_in_b_valid),
		.axi_resp_i_b_bits_id(_axi4frag_auto_in_b_bits_id),
		.axi_resp_i_b_bits_resp(_axi4frag_auto_in_b_bits_resp),
		.axi_resp_i_b_bits_user(1'h0),
		.axi_req_o_r_ready(_core_axi_req_o_r_ready),
		.axi_resp_i_r_valid(_axi4frag_auto_in_r_valid),
		.axi_resp_i_r_bits_id(_axi4frag_auto_in_r_bits_id),
		.axi_resp_i_r_bits_data(_axi4frag_auto_in_r_bits_data),
		.axi_resp_i_r_bits_resp(_axi4frag_auto_in_r_bits_resp),
		.axi_resp_i_r_bits_last(_axi4frag_auto_in_r_bits_last),
		.axi_resp_i_r_bits_user(1'h0)
	);
endmodule
module plusarg_reader (out);
	parameter FORMAT = "borked=%d";
	parameter WIDTH = 1;
	parameter [WIDTH - 1:0] DEFAULT = 0;
	output wire [WIDTH - 1:0] out;
	reg [WIDTH - 1:0] myplus;
	assign out = myplus;
	initial if (!$value$plusargs(FORMAT, myplus))
		myplus = DEFAULT;
endmodule
module alu (
	clk_i,
	rst_ni,
	fu_data_i,
	result_o,
	alu_branch_res_o
);
	input wire clk_i;
	input wire rst_ni;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	output reg [63:0] result_o;
	output reg alu_branch_res_o;
	wire [63:0] operand_a_rev;
	wire [31:0] operand_a_rev32;
	wire [riscv_XLEN:0] operand_b_neg;
	wire [65:0] adder_result_ext_o;
	reg less;
	genvar k;
	generate
		for (k = 0; k < riscv_XLEN; k = k + 1) begin : genblk1
			assign operand_a_rev[k] = fu_data_i[194 - (0 + k)];
		end
		for (k = 0; k < 32; k = k + 1) begin : genblk2
			assign operand_a_rev32[k] = fu_data_i[194 - (32 + k)];
		end
	endgenerate
	reg adder_op_b_negate;
	wire adder_z_flag;
	wire [riscv_XLEN:0] adder_in_a;
	wire [riscv_XLEN:0] adder_in_b;
	wire [63:0] adder_result;
	always @(*) begin
		adder_op_b_negate = 1'b0;
		case (fu_data_i[201-:7])
			7'd17, 7'd18, 7'd1, 7'd3: adder_op_b_negate = 1'b1;
			default:
				;
		endcase
	end
	assign adder_in_a = {fu_data_i[194-:64], 1'b1};
	assign operand_b_neg = {fu_data_i[130-:64], 1'b0} ^ {65 {adder_op_b_negate}};
	assign adder_in_b = operand_b_neg;
	assign adder_result_ext_o = $unsigned(adder_in_a) + $unsigned(adder_in_b);
	assign adder_result = adder_result_ext_o[riscv_XLEN:1];
	assign adder_z_flag = ~|adder_result;
	always @(*) begin : branch_resolve
		alu_branch_res_o = 1'b1;
		case (fu_data_i[201-:7])
			7'd17: alu_branch_res_o = adder_z_flag;
			7'd18: alu_branch_res_o = ~adder_z_flag;
			7'd13, 7'd14: alu_branch_res_o = less;
			7'd15, 7'd16: alu_branch_res_o = ~less;
			default: alu_branch_res_o = 1'b1;
		endcase
	end
	wire shift_left;
	wire shift_arithmetic;
	wire [63:0] shift_amt;
	wire [63:0] shift_op_a;
	wire [31:0] shift_op_a32;
	wire [63:0] shift_result;
	wire [31:0] shift_result32;
	wire [riscv_XLEN:0] shift_right_result;
	wire [32:0] shift_right_result32;
	wire [63:0] shift_left_result;
	wire [31:0] shift_left_result32;
	assign shift_amt = fu_data_i[130-:64];
	assign shift_left = (fu_data_i[201-:7] == 7'd9) | (fu_data_i[201-:7] == 7'd11);
	assign shift_arithmetic = (fu_data_i[201-:7] == 7'd7) | (fu_data_i[201-:7] == 7'd12);
	wire [riscv_XLEN:0] shift_op_a_64;
	wire [32:0] shift_op_a_32;
	assign shift_op_a = (shift_left ? operand_a_rev : fu_data_i[194-:64]);
	assign shift_op_a32 = (shift_left ? operand_a_rev32 : fu_data_i[162:131]);
	assign shift_op_a_64 = {shift_arithmetic & shift_op_a[63], shift_op_a};
	assign shift_op_a_32 = {shift_arithmetic & shift_op_a[31], shift_op_a32};
	assign shift_right_result = $unsigned($signed(shift_op_a_64) >>> shift_amt[5:0]);
	assign shift_right_result32 = $unsigned($signed(shift_op_a_32) >>> shift_amt[4:0]);
	genvar j;
	generate
		for (j = 0; j < riscv_XLEN; j = j + 1) begin : genblk3
			assign shift_left_result[j] = shift_right_result[63 - j];
		end
		for (j = 0; j < 32; j = j + 1) begin : genblk4
			assign shift_left_result32[j] = shift_right_result32[31 - j];
		end
	endgenerate
	assign shift_result = (shift_left ? shift_left_result : shift_right_result[63:0]);
	assign shift_result32 = (shift_left ? shift_left_result32 : shift_right_result32[31:0]);
	always @(*) begin : sv2v_autoblock_1
		reg sgn;
		sgn = 1'b0;
		if (((fu_data_i[201-:7] == 7'd21) || (fu_data_i[201-:7] == 7'd13)) || (fu_data_i[201-:7] == 7'd15))
			sgn = 1'b1;
		less = $signed({sgn & fu_data_i[194], fu_data_i[194-:64]}) < $signed({sgn & fu_data_i[130], fu_data_i[130-:64]});
	end
	always @(*) begin
		result_o = 1'sb0;
		case (fu_data_i[201-:7])
			7'd6: result_o = fu_data_i[194-:64] & fu_data_i[130-:64];
			7'd5: result_o = fu_data_i[194-:64] | fu_data_i[130-:64];
			7'd4: result_o = fu_data_i[194-:64] ^ fu_data_i[130-:64];
			7'd0, 7'd1: result_o = adder_result;
			7'd2, 7'd3: result_o = {{32 {adder_result[31]}}, adder_result[31:0]};
			7'd9, 7'd8, 7'd7: result_o = shift_result;
			7'd11, 7'd10, 7'd12: result_o = {{32 {shift_result32[31]}}, shift_result32[31:0]};
			7'd21, 7'd22: result_o = {{63 {1'b0}}, less};
			default:
				;
		endcase
	end
endmodule
module amo_buffer (
	clk_i,
	rst_ni,
	flush_i,
	valid_i,
	ready_o,
	amo_op_i,
	paddr_i,
	data_i,
	data_size_i,
	amo_req_o,
	amo_resp_i,
	amo_valid_commit_i,
	no_st_pending_i
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire valid_i;
	output wire ready_o;
	input wire [3:0] amo_op_i;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	input wire [55:0] paddr_i;
	input wire [63:0] data_i;
	input wire [1:0] data_size_i;
	output wire [134:0] amo_req_o;
	input wire [64:0] amo_resp_i;
	input wire amo_valid_commit_i;
	input wire no_st_pending_i;
	wire flush_amo_buffer;
	wire amo_valid;
	wire [125:0] amo_data_in;
	wire [125:0] amo_data_out;
	assign amo_req_o[134] = (no_st_pending_i & amo_valid_commit_i) & amo_valid;
	assign amo_req_o[133-:4] = amo_data_out[125-:4];
	assign amo_req_o[129-:2] = amo_data_out[1-:2];
	assign amo_req_o[127-:64] = {{8 {1'b0}}, amo_data_out[121-:56]};
	assign amo_req_o[63-:64] = {amo_data_out[65-:64]};
	assign amo_data_in[125-:4] = amo_op_i;
	assign amo_data_in[65-:64] = data_i;
	assign amo_data_in[121-:56] = paddr_i;
	assign amo_data_in[1-:2] = data_size_i;
	assign flush_amo_buffer = flush_i & !amo_valid_commit_i;
	fifo_v3_4F30F_AEF03 #(
		.dtype_riscv_PLEN(riscv_PLEN),
		.dtype_riscv_XLEN(riscv_XLEN),
		.DEPTH(1)
	) i_amo_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_amo_buffer),
		.testmode_i(1'b0),
		.full_o(amo_valid),
		.empty_o(ready_o),
		.usage_o(),
		.data_i(amo_data_in),
		.push_i(valid_i),
		.data_o(amo_data_out),
		.pop_i(amo_resp_i[64])
	);
endmodule
module ariane_regfile (
	clk_i,
	rst_ni,
	test_en_i,
	raddr_i,
	rdata_o,
	waddr_i,
	wdata_i,
	we_i
);
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] NR_READ_PORTS = 2;
	parameter [31:0] NR_WRITE_PORTS = 2;
	parameter [0:0] ZERO_REG_ZERO = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire test_en_i;
	input wire [(NR_READ_PORTS * 5) - 1:0] raddr_i;
	output wire [(NR_READ_PORTS * DATA_WIDTH) - 1:0] rdata_o;
	input wire [(NR_WRITE_PORTS * 5) - 1:0] waddr_i;
	input wire [(NR_WRITE_PORTS * DATA_WIDTH) - 1:0] wdata_i;
	input wire [NR_WRITE_PORTS - 1:0] we_i;
	localparam ADDR_WIDTH = 5;
	localparam NUM_WORDS = 32;
	reg [(32 * DATA_WIDTH) - 1:0] mem;
	reg [(NR_WRITE_PORTS * 32) - 1:0] we_dec;
	always @(*) begin : we_decoder
		begin : sv2v_autoblock_1
			reg [31:0] j;
			for (j = 0; j < NR_WRITE_PORTS; j = j + 1)
				begin : sv2v_autoblock_2
					reg [31:0] i;
					for (i = 0; i < NUM_WORDS; i = i + 1)
						if (waddr_i[j * 5+:5] == i)
							we_dec[(j * 32) + i] = we_i[j];
						else
							we_dec[(j * 32) + i] = 1'b0;
				end
		end
	end
	function automatic [DATA_WIDTH - 1:0] sv2v_cast_9134D;
		input reg [DATA_WIDTH - 1:0] inp;
		sv2v_cast_9134D = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : register_write_behavioral
		if (~rst_ni)
			mem <= {NUM_WORDS {sv2v_cast_9134D(1'sb0)}};
		else begin : sv2v_autoblock_3
			reg [31:0] j;
			for (j = 0; j < NR_WRITE_PORTS; j = j + 1)
				begin
					begin : sv2v_autoblock_4
						reg [31:0] i;
						for (i = 0; i < NUM_WORDS; i = i + 1)
							if (we_dec[(j * 32) + i])
								mem[i * DATA_WIDTH+:DATA_WIDTH] <= wdata_i[j * DATA_WIDTH+:DATA_WIDTH];
					end
					if (ZERO_REG_ZERO)
						mem[0+:DATA_WIDTH] <= 1'sb0;
				end
		end
	end
	genvar i;
	generate
		for (i = 0; i < NR_READ_PORTS; i = i + 1) begin : genblk1
			assign rdata_o[i * DATA_WIDTH+:DATA_WIDTH] = mem[raddr_i[i * 5+:5] * DATA_WIDTH+:DATA_WIDTH];
		end
	endgenerate
endmodule
module ariane (
	clk_i,
	rst_ni,
	boot_addr_i,
	hart_id_i,
	irq_i,
	ipi_i,
	time_irq_i,
	debug_req_i,
	axi_req_o,
	axi_resp_i
);
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire [63:0] boot_addr_i;
	input wire [63:0] hart_id_i;
	input wire [1:0] irq_i;
	input wire ipi_i;
	input wire time_irq_i;
	input wire debug_req_i;
	localparam ariane_axi_AddrWidth = 64;
	localparam ariane_axi_IdWidth = 4;
	localparam ariane_axi_UserWidth = 1;
	localparam ariane_axi_DataWidth = 64;
	localparam ariane_axi_StrbWidth = 8;
	output wire [280:0] axi_req_o;
	input wire [83:0] axi_resp_i;
	wire [1:0] priv_lvl;
	localparam riscv_XLEN = 64;
	wire [128:0] ex_commit;
	localparam riscv_VLEN = 64;
	wire [133:0] resolved_branch;
	wire [63:0] pc_commit;
	wire eret;
	localparam ariane_pkg_NR_COMMIT_PORTS = 2;
	wire [1:0] commit_ack;
	wire [63:0] trap_vector_base_commit_pcgen;
	wire [63:0] epc_commit_pcgen;
	wire [291:0] fetch_entry_if_id;
	wire fetch_valid_if_id;
	wire fetch_ready_id_if;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	wire [360:0] issue_entry_id_issue;
	wire issue_entry_valid_id_issue;
	wire is_ctrl_fow_id_issue;
	wire issue_instr_issue_id;
	wire [63:0] rs1_forwarding_id_ex;
	wire [63:0] rs2_forwarding_id_ex;
	wire [205:0] fu_data_id_ex;
	wire [63:0] pc_id_ex;
	wire is_compressed_instr_id_ex;
	wire flu_ready_ex_id;
	wire [2:0] flu_trans_id_ex_id;
	wire flu_valid_ex_id;
	wire [63:0] flu_result_ex_id;
	wire [128:0] flu_exception_ex_id;
	wire alu_valid_id_ex;
	wire branch_valid_id_ex;
	wire [66:0] branch_predict_id_ex;
	wire resolve_branch_ex_id;
	wire lsu_valid_id_ex;
	wire lsu_ready_ex_id;
	wire [2:0] load_trans_id_ex_id;
	wire [63:0] load_result_ex_id;
	wire load_valid_ex_id;
	wire [128:0] load_exception_ex_id;
	wire [63:0] store_result_ex_id;
	wire [2:0] store_trans_id_ex_id;
	wire store_valid_ex_id;
	wire [128:0] store_exception_ex_id;
	wire mult_valid_id_ex;
	wire fpu_ready_ex_id;
	wire fpu_valid_id_ex;
	wire [1:0] fpu_fmt_id_ex;
	wire [2:0] fpu_rm_id_ex;
	wire [2:0] fpu_trans_id_ex_id;
	wire [63:0] fpu_result_ex_id;
	wire fpu_valid_ex_id;
	wire [128:0] fpu_exception_ex_id;
	wire csr_valid_id_ex;
	wire csr_commit_commit_ex;
	wire dirty_fp_state;
	wire lsu_commit_commit_ex;
	wire lsu_commit_ready_ex_commit;
	wire [2:0] lsu_commit_trans_id;
	wire no_st_pending_ex;
	wire no_st_pending_commit;
	wire amo_valid_commit;
	wire [721:0] commit_instr_id_commit;
	wire [9:0] waddr_commit_id;
	wire [127:0] wdata_commit_id;
	wire [1:0] we_gpr_commit_id;
	wire [1:0] we_fpr_commit_id;
	wire [4:0] fflags_csr_commit;
	wire [1:0] fs;
	wire [2:0] frm_csr_id_issue_ex;
	wire [6:0] fprec_csr_ex;
	wire enable_translation_csr_ex;
	wire en_ld_st_translation_csr_ex;
	wire [1:0] ld_st_priv_lvl_csr_ex;
	wire sum_csr_ex;
	wire mxr_csr_ex;
	localparam riscv_PPNW = 44;
	wire [43:0] satp_ppn_csr_ex;
	localparam ariane_pkg_ASID_WIDTH = 16;
	wire [15:0] asid_csr_ex;
	wire [11:0] csr_addr_ex_csr;
	wire [6:0] csr_op_commit_csr;
	wire [63:0] csr_wdata_commit_csr;
	wire [63:0] csr_rdata_csr_commit;
	wire [128:0] csr_exception_csr_commit;
	wire tvm_csr_id;
	wire tw_csr_id;
	wire tsr_csr_id;
	wire [193:0] irq_ctrl_csr_id;
	wire dcache_en_csr_nbdcache;
	wire csr_write_fflags_commit_cs;
	wire icache_en_csr;
	wire debug_mode;
	wire single_step_csr_commit;
	wire [127:0] pmpcfg;
	localparam riscv_PLEN = 56;
	wire [863:0] pmpaddr;
	wire [4:0] addr_csr_perf;
	wire [63:0] data_csr_perf;
	wire [63:0] data_perf_csr;
	wire we_csr_perf;
	wire icache_flush_ctrl_cache;
	wire itlb_miss_ex_perf;
	wire dtlb_miss_ex_perf;
	wire dcache_miss_cache_perf;
	wire icache_miss_cache_perf;
	wire set_pc_ctrl_pcgen;
	wire flush_csr_ctrl;
	wire flush_unissued_instr_ctrl_id;
	wire flush_ctrl_if;
	wire flush_ctrl_id;
	wire flush_ctrl_ex;
	wire flush_ctrl_bp;
	wire flush_tlb_ctrl_ex;
	wire fence_i_commit_controller;
	wire fence_commit_controller;
	wire sfence_vma_commit_controller;
	wire halt_ctrl;
	wire halt_csr_ctrl;
	wire dcache_flush_ctrl_cache;
	wire dcache_flush_ack_cache_ctrl;
	wire set_debug_pc;
	wire flush_commit;
	wire [185:0] icache_areq_ex_cache;
	wire [64:0] icache_areq_cache_ex;
	wire [67:0] icache_dreq_if_cache;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	wire [226:0] icache_dreq_cache_if;
	wire [134:0] amo_req;
	wire [64:0] amo_resp;
	wire sb_full;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (3 * ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78)) - 1 : (3 * (1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 76)):(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)] dcache_req_ports_ex_cache;
	wire [197:0] dcache_req_ports_cache_ex;
	wire dcache_commit_wbuffer_empty;
	wire dcache_commit_wbuffer_not_ni;
	frontend #(.ArianeCfg(ArianeCfg)) i_frontend(
		.flush_i(flush_ctrl_if),
		.flush_bp_i(1'b0),
		.debug_mode_i(debug_mode),
		.boot_addr_i(boot_addr_i[63:0]),
		.icache_dreq_i(icache_dreq_cache_if),
		.icache_dreq_o(icache_dreq_if_cache),
		.resolved_branch_i(resolved_branch),
		.pc_commit_i(pc_commit),
		.set_pc_commit_i(set_pc_ctrl_pcgen),
		.set_debug_pc_i(set_debug_pc),
		.epc_i(epc_commit_pcgen),
		.eret_i(eret),
		.trap_vector_base_i(trap_vector_base_commit_pcgen),
		.ex_valid_i(ex_commit[0]),
		.fetch_entry_o(fetch_entry_if_id),
		.fetch_entry_valid_o(fetch_valid_if_id),
		.fetch_entry_ready_i(fetch_ready_id_if),
		.clk_i(clk_i),
		.rst_ni(rst_ni)
	);
	id_stage id_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_ctrl_if),
		.debug_req_i(debug_req_i),
		.fetch_entry_i(fetch_entry_if_id),
		.fetch_entry_valid_i(fetch_valid_if_id),
		.fetch_entry_ready_o(fetch_ready_id_if),
		.issue_entry_o(issue_entry_id_issue),
		.issue_entry_valid_o(issue_entry_valid_id_issue),
		.is_ctrl_flow_o(is_ctrl_fow_id_issue),
		.issue_instr_ack_i(issue_instr_issue_id),
		.priv_lvl_i(priv_lvl),
		.fs_i(fs),
		.frm_i(frm_csr_id_issue_ex),
		.irq_i(irq_i),
		.irq_ctrl_i(irq_ctrl_csr_id),
		.debug_mode_i(debug_mode),
		.tvm_i(tvm_csr_id),
		.tw_i(tw_csr_id),
		.tsr_i(tsr_csr_id)
	);
	localparam ariane_pkg_NR_WB_PORTS = 4;
	issue_stage #(
		.NR_ENTRIES(ariane_pkg_NR_SB_ENTRIES),
		.NR_WB_PORTS(ariane_pkg_NR_WB_PORTS),
		.NR_COMMIT_PORTS(ariane_pkg_NR_COMMIT_PORTS)
	) issue_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.sb_full_o(sb_full),
		.flush_unissued_instr_i(flush_unissued_instr_ctrl_id),
		.flush_i(flush_ctrl_id),
		.decoded_instr_i(issue_entry_id_issue),
		.decoded_instr_valid_i(issue_entry_valid_id_issue),
		.is_ctrl_flow_i(is_ctrl_fow_id_issue),
		.decoded_instr_ack_o(issue_instr_issue_id),
		.rs1_forwarding_o(rs1_forwarding_id_ex),
		.rs2_forwarding_o(rs2_forwarding_id_ex),
		.fu_data_o(fu_data_id_ex),
		.pc_o(pc_id_ex),
		.is_compressed_instr_o(is_compressed_instr_id_ex),
		.flu_ready_i(flu_ready_ex_id),
		.alu_valid_o(alu_valid_id_ex),
		.branch_valid_o(branch_valid_id_ex),
		.branch_predict_o(branch_predict_id_ex),
		.resolve_branch_i(resolve_branch_ex_id),
		.lsu_ready_i(lsu_ready_ex_id),
		.lsu_valid_o(lsu_valid_id_ex),
		.mult_valid_o(mult_valid_id_ex),
		.fpu_ready_i(fpu_ready_ex_id),
		.fpu_valid_o(fpu_valid_id_ex),
		.fpu_fmt_o(fpu_fmt_id_ex),
		.fpu_rm_o(fpu_rm_id_ex),
		.csr_valid_o(csr_valid_id_ex),
		.resolved_branch_i(resolved_branch),
		.trans_id_i({flu_trans_id_ex_id, load_trans_id_ex_id, store_trans_id_ex_id, fpu_trans_id_ex_id}),
		.wbdata_i({flu_result_ex_id, load_result_ex_id, store_result_ex_id, fpu_result_ex_id}),
		.ex_ex_i({flu_exception_ex_id, load_exception_ex_id, store_exception_ex_id, fpu_exception_ex_id}),
		.wt_valid_i({flu_valid_ex_id, load_valid_ex_id, store_valid_ex_id, fpu_valid_ex_id}),
		.waddr_i(waddr_commit_id),
		.wdata_i(wdata_commit_id),
		.we_gpr_i(we_gpr_commit_id),
		.we_fpr_i(we_fpr_commit_id),
		.commit_instr_o(commit_instr_id_commit),
		.commit_ack_i(commit_ack)
	);
	ex_stage #(
		.ASID_WIDTH(ariane_pkg_ASID_WIDTH),
		.ArianeCfg(ArianeCfg)
	) ex_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.debug_mode_i(debug_mode),
		.flush_i(flush_ctrl_ex),
		.rs1_forwarding_i(rs1_forwarding_id_ex),
		.rs2_forwarding_i(rs2_forwarding_id_ex),
		.fu_data_i(fu_data_id_ex),
		.pc_i(pc_id_ex),
		.is_compressed_instr_i(is_compressed_instr_id_ex),
		.flu_result_o(flu_result_ex_id),
		.flu_trans_id_o(flu_trans_id_ex_id),
		.flu_valid_o(flu_valid_ex_id),
		.flu_exception_o(flu_exception_ex_id),
		.flu_ready_o(flu_ready_ex_id),
		.alu_valid_i(alu_valid_id_ex),
		.branch_valid_i(branch_valid_id_ex),
		.branch_predict_i(branch_predict_id_ex),
		.resolved_branch_o(resolved_branch),
		.resolve_branch_o(resolve_branch_ex_id),
		.csr_valid_i(csr_valid_id_ex),
		.csr_addr_o(csr_addr_ex_csr),
		.csr_commit_i(csr_commit_commit_ex),
		.mult_valid_i(mult_valid_id_ex),
		.lsu_ready_o(lsu_ready_ex_id),
		.lsu_valid_i(lsu_valid_id_ex),
		.load_result_o(load_result_ex_id),
		.load_trans_id_o(load_trans_id_ex_id),
		.load_valid_o(load_valid_ex_id),
		.load_exception_o(load_exception_ex_id),
		.store_result_o(store_result_ex_id),
		.store_trans_id_o(store_trans_id_ex_id),
		.store_valid_o(store_valid_ex_id),
		.store_exception_o(store_exception_ex_id),
		.lsu_commit_i(lsu_commit_commit_ex),
		.lsu_commit_ready_o(lsu_commit_ready_ex_commit),
		.commit_tran_id_i(lsu_commit_trans_id),
		.no_st_pending_o(no_st_pending_ex),
		.fpu_ready_o(fpu_ready_ex_id),
		.fpu_valid_i(fpu_valid_id_ex),
		.fpu_fmt_i(fpu_fmt_id_ex),
		.fpu_rm_i(fpu_rm_id_ex),
		.fpu_frm_i(frm_csr_id_issue_ex),
		.fpu_prec_i(fprec_csr_ex),
		.fpu_trans_id_o(fpu_trans_id_ex_id),
		.fpu_result_o(fpu_result_ex_id),
		.fpu_valid_o(fpu_valid_ex_id),
		.fpu_exception_o(fpu_exception_ex_id),
		.amo_valid_commit_i(amo_valid_commit),
		.amo_req_o(amo_req),
		.amo_resp_i(amo_resp),
		.itlb_miss_o(itlb_miss_ex_perf),
		.dtlb_miss_o(dtlb_miss_ex_perf),
		.enable_translation_i(enable_translation_csr_ex),
		.en_ld_st_translation_i(en_ld_st_translation_csr_ex),
		.flush_tlb_i(flush_tlb_ctrl_ex),
		.priv_lvl_i(priv_lvl),
		.ld_st_priv_lvl_i(ld_st_priv_lvl_csr_ex),
		.sum_i(sum_csr_ex),
		.mxr_i(mxr_csr_ex),
		.satp_ppn_i(satp_ppn_csr_ex),
		.asid_i(asid_csr_ex),
		.icache_areq_i(icache_areq_cache_ex),
		.icache_areq_o(icache_areq_ex_cache),
		.dcache_req_ports_i(dcache_req_ports_cache_ex),
		.dcache_req_ports_o(dcache_req_ports_ex_cache),
		.dcache_wbuffer_empty_i(dcache_commit_wbuffer_empty),
		.dcache_wbuffer_not_ni_i(dcache_commit_wbuffer_not_ni),
		.pmpcfg_i(pmpcfg),
		.pmpaddr_i(pmpaddr)
	);
	assign no_st_pending_commit = no_st_pending_ex & dcache_commit_wbuffer_empty;
	commit_stage #(.NR_COMMIT_PORTS(ariane_pkg_NR_COMMIT_PORTS)) commit_stage_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.halt_i(halt_ctrl),
		.flush_dcache_i(dcache_flush_ctrl_cache),
		.exception_o(ex_commit),
		.dirty_fp_state_o(dirty_fp_state),
		.single_step_i(single_step_csr_commit),
		.commit_instr_i(commit_instr_id_commit),
		.commit_ack_o(commit_ack),
		.no_st_pending_i(no_st_pending_commit),
		.waddr_o(waddr_commit_id),
		.wdata_o(wdata_commit_id),
		.we_gpr_o(we_gpr_commit_id),
		.we_fpr_o(we_fpr_commit_id),
		.commit_lsu_o(lsu_commit_commit_ex),
		.commit_lsu_ready_i(lsu_commit_ready_ex_commit),
		.commit_tran_id_o(lsu_commit_trans_id),
		.amo_valid_commit_o(amo_valid_commit),
		.amo_resp_i(amo_resp),
		.commit_csr_o(csr_commit_commit_ex),
		.pc_o(pc_commit),
		.csr_op_o(csr_op_commit_csr),
		.csr_wdata_o(csr_wdata_commit_csr),
		.csr_rdata_i(csr_rdata_csr_commit),
		.csr_write_fflags_o(csr_write_fflags_commit_cs),
		.csr_exception_i(csr_exception_csr_commit),
		.fence_i_o(fence_i_commit_controller),
		.fence_o(fence_commit_controller),
		.sfence_vma_o(sfence_vma_commit_controller),
		.flush_commit_o(flush_commit)
	);
	csr_regfile #(
		.AsidWidth(ariane_pkg_ASID_WIDTH),
		.DmBaseAddress(ArianeCfg[95-:64]),
		.NrCommitPorts(ariane_pkg_NR_COMMIT_PORTS),
		.NrPMPEntries(ArianeCfg[31-:32])
	) csr_regfile_i(
		.flush_o(flush_csr_ctrl),
		.halt_csr_o(halt_csr_ctrl),
		.commit_instr_i(commit_instr_id_commit),
		.commit_ack_i(commit_ack),
		.boot_addr_i(boot_addr_i[63:0]),
		.hart_id_i(hart_id_i[63:0]),
		.ex_i(ex_commit),
		.csr_op_i(csr_op_commit_csr),
		.csr_write_fflags_i(csr_write_fflags_commit_cs),
		.dirty_fp_state_i(dirty_fp_state),
		.csr_addr_i(csr_addr_ex_csr),
		.csr_wdata_i(csr_wdata_commit_csr),
		.csr_rdata_o(csr_rdata_csr_commit),
		.pc_i(pc_commit),
		.csr_exception_o(csr_exception_csr_commit),
		.epc_o(epc_commit_pcgen),
		.eret_o(eret),
		.set_debug_pc_o(set_debug_pc),
		.trap_vector_base_o(trap_vector_base_commit_pcgen),
		.priv_lvl_o(priv_lvl),
		.fs_o(fs),
		.fflags_o(fflags_csr_commit),
		.frm_o(frm_csr_id_issue_ex),
		.fprec_o(fprec_csr_ex),
		.irq_ctrl_o(irq_ctrl_csr_id),
		.ld_st_priv_lvl_o(ld_st_priv_lvl_csr_ex),
		.en_translation_o(enable_translation_csr_ex),
		.en_ld_st_translation_o(en_ld_st_translation_csr_ex),
		.sum_o(sum_csr_ex),
		.mxr_o(mxr_csr_ex),
		.satp_ppn_o(satp_ppn_csr_ex),
		.asid_o(asid_csr_ex),
		.tvm_o(tvm_csr_id),
		.tw_o(tw_csr_id),
		.tsr_o(tsr_csr_id),
		.debug_mode_o(debug_mode),
		.single_step_o(single_step_csr_commit),
		.dcache_en_o(dcache_en_csr_nbdcache),
		.icache_en_o(icache_en_csr),
		.perf_addr_o(addr_csr_perf),
		.perf_data_o(data_csr_perf),
		.perf_data_i(data_perf_csr),
		.perf_we_o(we_csr_perf),
		.pmpcfg_o(pmpcfg),
		.pmpaddr_o(pmpaddr),
		.debug_req_i(debug_req_i),
		.ipi_i(ipi_i),
		.irq_i(irq_i),
		.time_irq_i(time_irq_i),
		.clk_i(clk_i),
		.rst_ni(rst_ni)
	);
	perf_counters i_perf_counters(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.debug_mode_i(debug_mode),
		.addr_i(addr_csr_perf),
		.we_i(we_csr_perf),
		.data_i(data_csr_perf),
		.data_o(data_perf_csr),
		.commit_instr_i(commit_instr_id_commit),
		.commit_ack_i(commit_ack),
		.l1_icache_miss_i(icache_miss_cache_perf),
		.l1_dcache_miss_i(dcache_miss_cache_perf),
		.itlb_miss_i(itlb_miss_ex_perf),
		.dtlb_miss_i(dtlb_miss_ex_perf),
		.sb_full_i(sb_full),
		.if_empty_i(~fetch_valid_if_id),
		.ex_i(ex_commit),
		.eret_i(eret),
		.resolved_branch_i(resolved_branch)
	);
	controller controller_i(
		.set_pc_commit_o(set_pc_ctrl_pcgen),
		.flush_unissued_instr_o(flush_unissued_instr_ctrl_id),
		.flush_if_o(flush_ctrl_if),
		.flush_id_o(flush_ctrl_id),
		.flush_ex_o(flush_ctrl_ex),
		.flush_bp_o(flush_ctrl_bp),
		.flush_tlb_o(flush_tlb_ctrl_ex),
		.flush_dcache_o(dcache_flush_ctrl_cache),
		.flush_dcache_ack_i(dcache_flush_ack_cache_ctrl),
		.halt_csr_i(halt_csr_ctrl),
		.halt_o(halt_ctrl),
		.eret_i(eret),
		.ex_valid_i(ex_commit[0]),
		.set_debug_pc_i(set_debug_pc),
		.flush_csr_i(flush_csr_ctrl),
		.resolved_branch_i(resolved_branch),
		.fence_i_i(fence_i_commit_controller),
		.fence_i(fence_commit_controller),
		.sfence_vma_i(sfence_vma_commit_controller),
		.flush_commit_i(flush_commit),
		.flush_icache_o(icache_flush_ctrl_cache),
		.clk_i(clk_i),
		.rst_ni(rst_ni)
	);
	wt_cache_subsystem #(.ArianeCfg(ArianeCfg)) i_cache_subsystem(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.icache_en_i(icache_en_csr),
		.icache_flush_i(icache_flush_ctrl_cache),
		.icache_miss_o(icache_miss_cache_perf),
		.icache_areq_i(icache_areq_ex_cache),
		.icache_areq_o(icache_areq_cache_ex),
		.icache_dreq_i(icache_dreq_if_cache),
		.icache_dreq_o(icache_dreq_cache_if),
		.dcache_enable_i(dcache_en_csr_nbdcache),
		.dcache_flush_i(dcache_flush_ctrl_cache),
		.dcache_flush_ack_o(dcache_flush_ack_cache_ctrl),
		.dcache_amo_req_i(amo_req),
		.dcache_amo_resp_o(amo_resp),
		.dcache_miss_o(dcache_miss_cache_perf),
		.dcache_req_ports_i(dcache_req_ports_ex_cache),
		.dcache_req_ports_o(dcache_req_ports_cache_ex),
		.wbuffer_empty_o(dcache_commit_wbuffer_empty),
		.wbuffer_not_ni_o(dcache_commit_wbuffer_not_ni),
		.axi_req_o(axi_req_o),
		.axi_resp_i(axi_resp_i)
	);
	reg signed [31:0] f;
	reg [63:0] cycles;
	initial f = $fopen("trace_hart_00.dasm", "w");
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			cycles <= 0;
		else begin : sv2v_autoblock_1
			reg signed [7:0] mode;
			mode = "";
			if (debug_mode)
				mode = "D";
			else
				case (priv_lvl)
					2'b11: mode = "M";
					2'b01: mode = "S";
					2'b00: mode = "U";
				endcase
			begin : sv2v_autoblock_2
				reg signed [31:0] i;
				for (i = 0; i < ariane_pkg_NR_COMMIT_PORTS; i = i + 1)
					if (commit_ack[i] && !commit_instr_id_commit[(i * 361) + 68])
						$fwrite(f, "%d 0x%0h %s (0x%h) DASM(%h)\n", cycles, commit_instr_id_commit[(i * 361) + 360-:64], mode, commit_instr_id_commit[(i * 361) + 100-:32], commit_instr_id_commit[(i * 361) + 100-:32]);
					else if (commit_ack[i] && commit_instr_id_commit[(i * 361) + 68]) begin
						if (commit_instr_id_commit[(i * 361) + 196-:64] == 2)
							$fwrite(f, "Exception Cause: Illegal Instructions, DASM(%h) PC=%h\n", commit_instr_id_commit[(i * 361) + 100-:32], commit_instr_id_commit[(i * 361) + 360-:64]);
						else if (debug_mode)
							$fwrite(f, "%d 0x%0h %s (0x%h) DASM(%h)\n", cycles, commit_instr_id_commit[(i * 361) + 360-:64], mode, commit_instr_id_commit[(i * 361) + 100-:32], commit_instr_id_commit[(i * 361) + 100-:32]);
						else
							$fwrite(f, "Exception Cause: %5d, DASM(%h) PC=%h\n", commit_instr_id_commit[(i * 361) + 196-:64], commit_instr_id_commit[(i * 361) + 100-:32], commit_instr_id_commit[(i * 361) + 360-:64]);
					end
			end
			cycles <= cycles + 1;
		end
	// final $fclose(f);
endmodule
module axi_shim (
	clk_i,
	rst_ni,
	rd_req_i,
	rd_gnt_o,
	rd_addr_i,
	rd_blen_i,
	rd_size_i,
	rd_id_i,
	rd_lock_i,
	rd_rdy_i,
	rd_last_o,
	rd_valid_o,
	rd_data_o,
	rd_id_o,
	rd_exokay_o,
	wr_req_i,
	wr_gnt_o,
	wr_addr_i,
	wr_data_i,
	wr_be_i,
	wr_blen_i,
	wr_size_i,
	wr_id_i,
	wr_lock_i,
	wr_atop_i,
	wr_rdy_i,
	wr_valid_o,
	wr_id_o,
	wr_exokay_o,
	axi_req_o,
	axi_resp_i
);
	parameter [31:0] AxiNumWords = 4;
	parameter [31:0] AxiIdWidth = 4;
	input wire clk_i;
	input wire rst_ni;
	input wire rd_req_i;
	output wire rd_gnt_o;
	input wire [63:0] rd_addr_i;
	input wire [$clog2(AxiNumWords) - 1:0] rd_blen_i;
	input wire [1:0] rd_size_i;
	input wire [AxiIdWidth - 1:0] rd_id_i;
	input wire rd_lock_i;
	input wire rd_rdy_i;
	output wire rd_last_o;
	output wire rd_valid_o;
	output wire [63:0] rd_data_o;
	output wire [AxiIdWidth - 1:0] rd_id_o;
	output wire rd_exokay_o;
	input wire wr_req_i;
	output reg wr_gnt_o;
	input wire [63:0] wr_addr_i;
	input wire [(AxiNumWords * 64) - 1:0] wr_data_i;
	input wire [(AxiNumWords * 8) - 1:0] wr_be_i;
	input wire [$clog2(AxiNumWords) - 1:0] wr_blen_i;
	input wire [1:0] wr_size_i;
	input wire [AxiIdWidth - 1:0] wr_id_i;
	input wire wr_lock_i;
	input wire [5:0] wr_atop_i;
	input wire wr_rdy_i;
	output wire wr_valid_o;
	output wire [AxiIdWidth - 1:0] wr_id_o;
	output wire wr_exokay_o;
	localparam ariane_axi_AddrWidth = 64;
	localparam ariane_axi_IdWidth = 4;
	localparam ariane_axi_UserWidth = 1;
	localparam ariane_axi_DataWidth = 64;
	localparam ariane_axi_StrbWidth = 8;
	output reg [280:0] axi_req_o;
	input wire [83:0] axi_resp_i;
	localparam AddrIndex = ($clog2(AxiNumWords) > 0 ? $clog2(AxiNumWords) : 1);
	reg [3:0] wr_state_q;
	reg [3:0] wr_state_d;
	wire [AddrIndex - 1:0] wr_cnt_d;
	reg [AddrIndex - 1:0] wr_cnt_q;
	wire wr_single_req;
	wire wr_cnt_done;
	reg wr_cnt_clr;
	reg wr_cnt_en;
	assign wr_single_req = wr_blen_i == 0;
	localparam axi_pkg_BURST_INCR = 2'b01;
	wire [2:1] sv2v_tmp_6E9DC;
	assign sv2v_tmp_6E9DC = axi_pkg_BURST_INCR;
	always @(*) axi_req_o[201-:2] = sv2v_tmp_6E9DC;
	wire [64:1] sv2v_tmp_930DC;
	assign sv2v_tmp_930DC = wr_addr_i;
	always @(*) axi_req_o[276-:64] = sv2v_tmp_930DC;
	wire [3:1] sv2v_tmp_448EB;
	assign sv2v_tmp_448EB = wr_size_i;
	always @(*) axi_req_o[204-:3] = sv2v_tmp_448EB;
	wire [8:1] sv2v_tmp_8D74F;
	assign sv2v_tmp_8D74F = wr_blen_i;
	always @(*) axi_req_o[212-:8] = sv2v_tmp_8D74F;
	wire [4:1] sv2v_tmp_96550;
	assign sv2v_tmp_96550 = wr_id_i;
	always @(*) axi_req_o[280-:4] = sv2v_tmp_96550;
	wire [3:1] sv2v_tmp_B8D42;
	assign sv2v_tmp_B8D42 = 3'b000;
	always @(*) axi_req_o[194-:3] = sv2v_tmp_B8D42;
	wire [4:1] sv2v_tmp_88B04;
	assign sv2v_tmp_88B04 = 4'b0000;
	always @(*) axi_req_o[187-:4] = sv2v_tmp_88B04;
	wire [1:1] sv2v_tmp_2B037;
	assign sv2v_tmp_2B037 = wr_lock_i;
	always @(*) axi_req_o[199] = sv2v_tmp_2B037;
	wire [4:1] sv2v_tmp_D3810;
	assign sv2v_tmp_D3810 = 4'b0000;
	always @(*) axi_req_o[198-:4] = sv2v_tmp_D3810;
	wire [4:1] sv2v_tmp_32328;
	assign sv2v_tmp_32328 = 4'b0000;
	always @(*) axi_req_o[191-:4] = sv2v_tmp_32328;
	wire [6:1] sv2v_tmp_FD09F;
	assign sv2v_tmp_FD09F = wr_atop_i;
	always @(*) axi_req_o[183-:6] = sv2v_tmp_FD09F;
	wire [64:1] sv2v_tmp_96288;
	assign sv2v_tmp_96288 = wr_data_i[wr_cnt_q * 64+:64];
	always @(*) axi_req_o[175-:64] = sv2v_tmp_96288;
	wire [8:1] sv2v_tmp_CF23C;
	assign sv2v_tmp_CF23C = wr_be_i[wr_cnt_q * 8+:8];
	always @(*) axi_req_o[111-:8] = sv2v_tmp_CF23C;
	wire [1:1] sv2v_tmp_1AB64;
	assign sv2v_tmp_1AB64 = wr_cnt_done;
	always @(*) axi_req_o[103] = sv2v_tmp_1AB64;
	localparam axi_pkg_RESP_EXOKAY = 2'b01;
	assign wr_exokay_o = axi_resp_i[75-:2] == axi_pkg_RESP_EXOKAY;
	wire [1:1] sv2v_tmp_3E233;
	assign sv2v_tmp_3E233 = wr_rdy_i;
	always @(*) axi_req_o[100] = sv2v_tmp_3E233;
	assign wr_valid_o = axi_resp_i[80];
	assign wr_id_o = axi_resp_i[79-:4];
	assign wr_cnt_done = wr_cnt_q == wr_blen_i;
	assign wr_cnt_d = (wr_cnt_clr ? {AddrIndex {1'sb0}} : (wr_cnt_en ? wr_cnt_q + 1 : wr_cnt_q));
	always @(*) begin : p_axi_write_fsm
		wr_state_d = wr_state_q;
		axi_req_o[176] = 1'b0;
		axi_req_o[101] = 1'b0;
		wr_gnt_o = 1'b0;
		wr_cnt_en = 1'b0;
		wr_cnt_clr = 1'b0;
		case (wr_state_q)
			4'd0:
				if (wr_req_i) begin
					axi_req_o[176] = 1'b1;
					axi_req_o[101] = 1'b1;
					if (wr_single_req) begin
						wr_cnt_clr = 1'b1;
						wr_gnt_o = axi_resp_i[83] & axi_resp_i[81];
						case ({axi_resp_i[83], axi_resp_i[81]})
							2'b01: wr_state_d = 4'd1;
							2'b10: wr_state_d = 4'd2;
							default: wr_state_d = 4'd0;
						endcase
					end
					else begin
						wr_cnt_en = axi_resp_i[81];
						case ({axi_resp_i[83], axi_resp_i[81]})
							2'b11: wr_state_d = 4'd2;
							2'b01: wr_state_d = 4'd3;
							2'b10: wr_state_d = 4'd2;
							default:
								;
						endcase
					end
				end
			4'd1: begin
				axi_req_o[176] = 1'b1;
				if (axi_resp_i[83]) begin
					wr_state_d = 4'd0;
					wr_gnt_o = 1'b1;
				end
			end
			4'd3: begin
				axi_req_o[101] = 1'b1;
				axi_req_o[176] = 1'b1;
				case ({axi_resp_i[83], axi_resp_i[81]})
					2'b01:
						if (wr_cnt_done) begin
							wr_state_d = 4'd4;
							wr_cnt_clr = 1'b1;
						end
						else
							wr_cnt_en = 1'b1;
					2'b10: wr_state_d = 4'd2;
					2'b11:
						if (wr_cnt_done) begin
							wr_state_d = 4'd0;
							wr_gnt_o = 1'b1;
							wr_cnt_clr = 1'b1;
						end
						else begin
							wr_state_d = 4'd2;
							wr_cnt_en = 1'b1;
						end
					default:
						;
				endcase
			end
			4'd4: begin
				axi_req_o[176] = 1'b1;
				if (axi_resp_i[83]) begin
					wr_state_d = 4'd0;
					wr_gnt_o = 1'b1;
				end
			end
			4'd2: begin
				axi_req_o[101] = 1'b1;
				if (wr_cnt_done) begin
					if (axi_resp_i[81]) begin
						wr_state_d = 4'd0;
						wr_cnt_clr = 1'b1;
						wr_gnt_o = 1'b1;
					end
				end
				else if (axi_resp_i[81])
					wr_cnt_en = 1'b1;
			end
			default: wr_state_d = 4'd0;
		endcase
	end
	wire [2:1] sv2v_tmp_20CF9;
	assign sv2v_tmp_20CF9 = axi_pkg_BURST_INCR;
	always @(*) axi_req_o[20-:2] = sv2v_tmp_20CF9;
	wire [64:1] sv2v_tmp_975D7;
	assign sv2v_tmp_975D7 = rd_addr_i;
	always @(*) axi_req_o[95-:64] = sv2v_tmp_975D7;
	wire [3:1] sv2v_tmp_2B990;
	assign sv2v_tmp_2B990 = rd_size_i;
	always @(*) axi_req_o[23-:3] = sv2v_tmp_2B990;
	wire [8:1] sv2v_tmp_E0E65;
	assign sv2v_tmp_E0E65 = rd_blen_i;
	always @(*) axi_req_o[31-:8] = sv2v_tmp_E0E65;
	wire [4:1] sv2v_tmp_7B90C;
	assign sv2v_tmp_7B90C = rd_id_i;
	always @(*) axi_req_o[99-:4] = sv2v_tmp_7B90C;
	wire [3:1] sv2v_tmp_A8AC6;
	assign sv2v_tmp_A8AC6 = 3'b000;
	always @(*) axi_req_o[13-:3] = sv2v_tmp_A8AC6;
	wire [4:1] sv2v_tmp_49C20;
	assign sv2v_tmp_49C20 = 4'b0000;
	always @(*) axi_req_o[6-:4] = sv2v_tmp_49C20;
	wire [1:1] sv2v_tmp_99F91;
	assign sv2v_tmp_99F91 = rd_lock_i;
	always @(*) axi_req_o[18] = sv2v_tmp_99F91;
	wire [4:1] sv2v_tmp_042AF;
	assign sv2v_tmp_042AF = 4'b0000;
	always @(*) axi_req_o[17-:4] = sv2v_tmp_042AF;
	wire [4:1] sv2v_tmp_F01FC;
	assign sv2v_tmp_F01FC = 4'b0000;
	always @(*) axi_req_o[10-:4] = sv2v_tmp_F01FC;
	wire [1:1] sv2v_tmp_8FD7F;
	assign sv2v_tmp_8FD7F = rd_req_i;
	always @(*) axi_req_o[1] = sv2v_tmp_8FD7F;
	assign rd_gnt_o = rd_req_i & axi_resp_i[82];
	wire [1:1] sv2v_tmp_967F1;
	assign sv2v_tmp_967F1 = rd_rdy_i;
	always @(*) axi_req_o[0] = sv2v_tmp_967F1;
	assign rd_data_o = axi_resp_i[67-:64];
	assign rd_last_o = axi_resp_i[1];
	assign rd_valid_o = axi_resp_i[72];
	assign rd_id_o = axi_resp_i[71-:4];
	assign rd_exokay_o = axi_resp_i[3-:2] == axi_pkg_RESP_EXOKAY;
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			wr_state_q <= 4'd0;
			wr_cnt_q <= 1'sb0;
		end
		else begin
			wr_state_q <= wr_state_d;
			wr_cnt_q <= wr_cnt_d;
		end
endmodule
module branch_unit (
	clk_i,
	rst_ni,
	debug_mode_i,
	fu_data_i,
	pc_i,
	is_compressed_instr_i,
	fu_valid_i,
	branch_valid_i,
	branch_comp_res_i,
	branch_result_o,
	branch_predict_i,
	resolved_branch_o,
	resolve_branch_o,
	branch_exception_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire debug_mode_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	localparam riscv_VLEN = 64;
	input wire [63:0] pc_i;
	input wire is_compressed_instr_i;
	input wire fu_valid_i;
	input wire branch_valid_i;
	input wire branch_comp_res_i;
	output reg [63:0] branch_result_o;
	input wire [66:0] branch_predict_i;
	output reg [133:0] resolved_branch_o;
	output reg resolve_branch_o;
	output reg [128:0] branch_exception_o;
	reg [63:0] target_address;
	reg [63:0] next_pc;
	function automatic ariane_pkg_op_is_branch;
		input reg [6:0] op;
		if (|{op == 7'd17, op == 7'd18, op == 7'd13, op == 7'd15, op == 7'd14, op == 7'd16})
			ariane_pkg_op_is_branch = 1'b1;
		else
			ariane_pkg_op_is_branch = 1'b0;
	endfunction
	always @(*) begin : mispredict_handler
		reg [63:0] jump_base;
		jump_base = (fu_data_i[201-:7] == 7'd19 ? fu_data_i[194:131] : pc_i);
		target_address = {riscv_VLEN {1'b0}};
		resolve_branch_o = 1'b0;
		resolved_branch_o[68-:64] = {riscv_VLEN {1'b0}};
		resolved_branch_o[3] = 1'b0;
		resolved_branch_o[133] = branch_valid_i;
		resolved_branch_o[4] = 1'b0;
		resolved_branch_o[2-:3] = branch_predict_i[66-:3];
		next_pc = pc_i + (is_compressed_instr_i ? {{62 {1'b0}}, 2'h2} : {{61 {1'b0}}, 3'h4});
		target_address = $unsigned($signed(jump_base) + $signed(fu_data_i[66:3]));
		if (fu_data_i[201-:7] == 7'd19)
			target_address[0] = 1'b0;
		branch_result_o = next_pc;
		resolved_branch_o[132-:64] = pc_i;
		if (branch_valid_i) begin
			resolved_branch_o[68-:64] = (branch_comp_res_i ? target_address : next_pc);
			resolved_branch_o[3] = branch_comp_res_i;
			if (ariane_pkg_op_is_branch(fu_data_i[201-:7]) && (branch_comp_res_i != (branch_predict_i[66-:3] == 3'd1))) begin
				resolved_branch_o[4] = 1'b1;
				resolved_branch_o[2-:3] = 3'd1;
			end
			if ((fu_data_i[201-:7] == 7'd19) && ((branch_predict_i[66-:3] == 3'd0) || (target_address != branch_predict_i[63-:riscv_VLEN]))) begin
				resolved_branch_o[4] = 1'b1;
				if (branch_predict_i[66-:3] != 3'd4)
					resolved_branch_o[2-:3] = 3'd3;
			end
			resolve_branch_o = 1'b1;
		end
	end
	localparam [63:0] riscv_INSTR_ADDR_MISALIGNED = 0;
	always @(*) begin : exception_handling
		branch_exception_o[128-:64] = riscv_INSTR_ADDR_MISALIGNED;
		branch_exception_o[0] = 1'b0;
		branch_exception_o[64-:64] = {pc_i};
		if (branch_valid_i && (target_address[0] != 1'b0))
			branch_exception_o[0] = 1'b1;
	end
endmodule
module commit_stage (
	clk_i,
	rst_ni,
	halt_i,
	flush_dcache_i,
	exception_o,
	dirty_fp_state_o,
	single_step_i,
	commit_instr_i,
	commit_ack_o,
	waddr_o,
	wdata_o,
	we_gpr_o,
	we_fpr_o,
	amo_resp_i,
	pc_o,
	csr_op_o,
	csr_wdata_o,
	csr_rdata_i,
	csr_exception_i,
	csr_write_fflags_o,
	commit_lsu_o,
	commit_lsu_ready_i,
	commit_tran_id_o,
	amo_valid_commit_o,
	no_st_pending_i,
	commit_csr_o,
	fence_i_o,
	fence_o,
	flush_commit_o,
	sfence_vma_o
);
	parameter [31:0] NR_COMMIT_PORTS = 2;
	input wire clk_i;
	input wire rst_ni;
	input wire halt_i;
	input wire flush_dcache_i;
	localparam riscv_XLEN = 64;
	output reg [128:0] exception_o;
	output reg dirty_fp_state_o;
	input wire single_step_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_VLEN = 64;
	input wire [(NR_COMMIT_PORTS * 361) - 1:0] commit_instr_i;
	output reg [NR_COMMIT_PORTS - 1:0] commit_ack_o;
	output wire [(NR_COMMIT_PORTS * 5) - 1:0] waddr_o;
	output reg [(NR_COMMIT_PORTS * 64) - 1:0] wdata_o;
	output reg [NR_COMMIT_PORTS - 1:0] we_gpr_o;
	output reg [NR_COMMIT_PORTS - 1:0] we_fpr_o;
	input wire [64:0] amo_resp_i;
	output wire [63:0] pc_o;
	output reg [6:0] csr_op_o;
	output reg [63:0] csr_wdata_o;
	input wire [63:0] csr_rdata_i;
	input wire [128:0] csr_exception_i;
	output reg csr_write_fflags_o;
	output reg commit_lsu_o;
	input wire commit_lsu_ready_i;
	output wire [2:0] commit_tran_id_o;
	output reg amo_valid_commit_o;
	input wire no_st_pending_i;
	output reg commit_csr_o;
	output reg fence_i_o;
	output reg fence_o;
	output reg flush_commit_o;
	output reg sfence_vma_o;
	genvar i;
	generate
		for (i = 0; i < NR_COMMIT_PORTS; i = i + 1) begin : gen_waddr
			assign waddr_o[i * 5+:5] = commit_instr_i[(i * 361) + 269-:5];
		end
	endgenerate
	assign pc_o = commit_instr_i[360-:64];
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	function automatic ariane_pkg_is_rd_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd81 <= op) && (7'd84 >= op), (7'd89 <= op) && (7'd98 >= op), op == 7'd100, op == 7'd101, op == 7'd102, op == 7'd104, (7'd107 <= op) && (7'd111 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rd_fpr = 1'b1;
			else
				ariane_pkg_is_rd_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rd_fpr = 1'b0;
	endfunction
	always @(*) begin : dirty_fp_state
		dirty_fp_state_o = 1'b0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < NR_COMMIT_PORTS; i = i + 1)
				dirty_fp_state_o = dirty_fp_state_o | (commit_ack_o[i] & (|{commit_instr_i[(i * 361) + 293-:4] == 4'd7, commit_instr_i[(i * 361) + 293-:4] == 4'd8} || ariane_pkg_is_rd_fpr(commit_instr_i[(i * 361) + 289-:7])));
		end
	end
	assign commit_tran_id_o = commit_instr_i[296-:3];
	wire instr_0_is_amo;
	function automatic ariane_pkg_is_amo;
		input reg [6:0] op;
		if ((7'd46 <= op) && (7'd67 >= op))
			ariane_pkg_is_amo = 1'b1;
		else
			ariane_pkg_is_amo = 1'b0;
	endfunction
	assign instr_0_is_amo = ariane_pkg_is_amo(commit_instr_i[289-:7]);
	localparam [0:0] ariane_pkg_RVA = 1'b1;
	always @(*) begin : commit
		commit_ack_o[0] = 1'b0;
		commit_ack_o[1] = 1'b0;
		amo_valid_commit_o = 1'b0;
		we_gpr_o[0] = 1'b0;
		we_gpr_o[1] = 1'b0;
		we_fpr_o = {NR_COMMIT_PORTS {1'b0}};
		commit_lsu_o = 1'b0;
		commit_csr_o = 1'b0;
		wdata_o[0+:64] = (amo_resp_i[64] ? amo_resp_i[63:0] : commit_instr_i[264-:64]);
		wdata_o[64+:64] = commit_instr_i[625-:64];
		csr_op_o = 7'd0;
		csr_wdata_o = {riscv_XLEN {1'b0}};
		fence_i_o = 1'b0;
		fence_o = 1'b0;
		sfence_vma_o = 1'b0;
		csr_write_fflags_o = 1'b0;
		flush_commit_o = 1'b0;
		if ((commit_instr_i[200] && !commit_instr_i[68]) && !halt_i) begin
			commit_ack_o[0] = 1'b1;
			if (ariane_pkg_is_rd_fpr(commit_instr_i[289-:7]))
				we_fpr_o[0] = 1'b1;
			else
				we_gpr_o[0] = 1'b1;
			if ((commit_instr_i[293-:4] == 4'd2) && !instr_0_is_amo) begin
				if (commit_lsu_ready_i) begin
					commit_ack_o[0] = 1'b1;
					commit_lsu_o = 1'b1;
				end
				else
					commit_ack_o[0] = 1'b0;
			end
			if (|{commit_instr_i[293-:4] == 4'd7, commit_instr_i[293-:4] == 4'd8}) begin
				csr_wdata_o = {{59 {1'b0}}, commit_instr_i[137-:5]};
				csr_write_fflags_o = 1'b1;
				commit_ack_o[0] = 1'b1;
			end
			if (commit_instr_i[293-:4] == 4'd6) begin
				csr_op_o = commit_instr_i[289-:7];
				csr_wdata_o = commit_instr_i[264-:64];
				if (!csr_exception_i[0]) begin
					commit_csr_o = 1'b1;
					wdata_o[0+:64] = csr_rdata_i;
					commit_ack_o[0] = 1'b1;
				end
				else begin
					commit_ack_o[0] = 1'b0;
					we_gpr_o[0] = 1'b0;
				end
			end
			if (commit_instr_i[289-:7] == 7'd30) begin
				sfence_vma_o = no_st_pending_i;
				commit_ack_o[0] = no_st_pending_i;
			end
			if ((commit_instr_i[289-:7] == 7'd29) || (flush_dcache_i && (commit_instr_i[293-:4] != 4'd2))) begin
				commit_ack_o[0] = no_st_pending_i;
				fence_i_o = no_st_pending_i;
			end
			if (commit_instr_i[289-:7] == 7'd28) begin
				commit_ack_o[0] = no_st_pending_i;
				fence_o = no_st_pending_i;
			end
			if (ariane_pkg_RVA && instr_0_is_amo) begin
				commit_ack_o[0] = amo_resp_i[64];
				flush_commit_o = amo_resp_i[64];
				amo_valid_commit_o = 1'b1;
				we_gpr_o[0] = amo_resp_i[64];
			end
		end
		if (NR_COMMIT_PORTS > 1) begin
			if ((((((commit_ack_o[0] && commit_instr_i[561]) && !halt_i) && (commit_instr_i[293-:4] != 4'd6)) && !flush_dcache_i) && !instr_0_is_amo) && !single_step_i) begin
				if ((!exception_o[0] && !commit_instr_i[429]) && |{commit_instr_i[654-:4] == 4'd3, commit_instr_i[654-:4] == 4'd1, commit_instr_i[654-:4] == 4'd4, commit_instr_i[654-:4] == 4'd5, commit_instr_i[654-:4] == 4'd7, commit_instr_i[654-:4] == 4'd8}) begin
					if (ariane_pkg_is_rd_fpr(commit_instr_i[650-:7]))
						we_fpr_o[1] = 1'b1;
					else
						we_gpr_o[1] = 1'b1;
					commit_ack_o[1] = 1'b1;
					if (|{commit_instr_i[654-:4] == 4'd7, commit_instr_i[654-:4] == 4'd8}) begin
						if (csr_write_fflags_o)
							csr_wdata_o = {{59 {1'b0}}, commit_instr_i[137-:5] | commit_instr_i[498-:5]};
						else
							csr_wdata_o = {{59 {1'b0}}, commit_instr_i[498-:5]};
						csr_write_fflags_o = 1'b1;
					end
				end
			end
		end
	end
	always @(*) begin : exception_handling
		exception_o[0] = 1'b0;
		exception_o[128-:64] = 1'sb0;
		exception_o[64-:64] = 1'sb0;
		if (commit_instr_i[200]) begin
			if (csr_exception_i[0]) begin
				exception_o = csr_exception_i;
				exception_o[64-:64] = commit_instr_i[132-:64];
			end
			if (commit_instr_i[68])
				exception_o = commit_instr_i[196-:129];
		end
		if (halt_i)
			exception_o[0] = 1'b0;
	end
endmodule
module compressed_decoder (
	instr_i,
	instr_o,
	illegal_instr_o,
	is_compressed_o
);
	input wire [31:0] instr_i;
	output reg [31:0] instr_o;
	output reg illegal_instr_o;
	output reg is_compressed_o;
	localparam riscv_OpcodeBranch = 7'b1100011;
	localparam riscv_OpcodeC0 = 2'b00;
	localparam riscv_OpcodeC0Addi4spn = 3'b000;
	localparam riscv_OpcodeC0Fld = 3'b001;
	localparam riscv_OpcodeC0Fsd = 3'b101;
	localparam riscv_OpcodeC0Ld = 3'b011;
	localparam riscv_OpcodeC0Lw = 3'b010;
	localparam riscv_OpcodeC0Sd = 3'b111;
	localparam riscv_OpcodeC0Sw = 3'b110;
	localparam riscv_OpcodeC1 = 2'b01;
	localparam riscv_OpcodeC1Addi = 3'b000;
	localparam riscv_OpcodeC1Addiw = 3'b001;
	localparam riscv_OpcodeC1Beqz = 3'b110;
	localparam riscv_OpcodeC1Bnez = 3'b111;
	localparam riscv_OpcodeC1J = 3'b101;
	localparam riscv_OpcodeC1Li = 3'b010;
	localparam riscv_OpcodeC1LuiAddi16sp = 3'b011;
	localparam riscv_OpcodeC1MiscAlu = 3'b100;
	localparam riscv_OpcodeC2 = 2'b10;
	localparam riscv_OpcodeC2Fldsp = 3'b001;
	localparam riscv_OpcodeC2Fsdsp = 3'b101;
	localparam riscv_OpcodeC2JalrMvAdd = 3'b100;
	localparam riscv_OpcodeC2Ldsp = 3'b011;
	localparam riscv_OpcodeC2Lwsp = 3'b010;
	localparam riscv_OpcodeC2Sdsp = 3'b111;
	localparam riscv_OpcodeC2Slli = 3'b000;
	localparam riscv_OpcodeC2Swsp = 3'b110;
	localparam riscv_OpcodeJal = 7'b1101111;
	localparam riscv_OpcodeJalr = 7'b1100111;
	localparam riscv_OpcodeLoad = 7'b0000011;
	localparam riscv_OpcodeLoadFp = 7'b0000111;
	localparam riscv_OpcodeLui = 7'b0110111;
	localparam riscv_OpcodeOp = 7'b0110011;
	localparam riscv_OpcodeOp32 = 7'b0111011;
	localparam riscv_OpcodeOpImm = 7'b0010011;
	localparam riscv_OpcodeOpImm32 = 7'b0011011;
	localparam riscv_OpcodeStore = 7'b0100011;
	localparam riscv_OpcodeStoreFp = 7'b0100111;
	localparam riscv_XLEN = 64;
	always @(*) begin
		illegal_instr_o = 1'b0;
		instr_o = 1'sb0;
		is_compressed_o = 1'b1;
		instr_o = instr_i;
		case (instr_i[1:0])
			riscv_OpcodeC0:
				case (instr_i[15:13])
					riscv_OpcodeC0Addi4spn: begin
						instr_o = {2'b00, instr_i[10:7], instr_i[12:11], instr_i[5], instr_i[6], 12'h041, instr_i[4:2], riscv_OpcodeOpImm};
						if (instr_i[12:5] == 8'b00000000)
							illegal_instr_o = 1'b1;
					end
					riscv_OpcodeC0Fld: instr_o = {4'b0000, instr_i[6:5], instr_i[12:10], 5'b00001, instr_i[9:7], 5'b01101, instr_i[4:2], riscv_OpcodeLoadFp};
					riscv_OpcodeC0Lw: instr_o = {5'b00000, instr_i[5], instr_i[12:10], instr_i[6], 4'b0001, instr_i[9:7], 5'b01001, instr_i[4:2], riscv_OpcodeLoad};
					riscv_OpcodeC0Ld: instr_o = {4'b0000, instr_i[6:5], instr_i[12:10], 5'b00001, instr_i[9:7], 5'b01101, instr_i[4:2], riscv_OpcodeLoad};
					riscv_OpcodeC0Fsd: instr_o = {4'b0000, instr_i[6:5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b011, instr_i[11:10], 3'b000, riscv_OpcodeStoreFp};
					riscv_OpcodeC0Sw: instr_o = {5'b00000, instr_i[5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b010, instr_i[11:10], instr_i[6], 2'b00, riscv_OpcodeStore};
					riscv_OpcodeC0Sd: instr_o = {4'b0000, instr_i[6:5], instr_i[12], 2'b01, instr_i[4:2], 2'b01, instr_i[9:7], 3'b011, instr_i[11:10], 3'b000, riscv_OpcodeStore};
					default: illegal_instr_o = 1'b1;
				endcase
			riscv_OpcodeC1:
				case (instr_i[15:13])
					riscv_OpcodeC1Addi: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], riscv_OpcodeOpImm};
					riscv_OpcodeC1Addiw:
						if (instr_i[11:7] != 5'h00)
							instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], riscv_OpcodeOpImm32};
						else
							illegal_instr_o = 1'b1;
					riscv_OpcodeC1Li: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 8'b00000000, instr_i[11:7], riscv_OpcodeOpImm};
					riscv_OpcodeC1LuiAddi16sp: begin
						instr_o = {{15 {instr_i[12]}}, instr_i[6:2], instr_i[11:7], riscv_OpcodeLui};
						if (instr_i[11:7] == 5'h02)
							instr_o = {{3 {instr_i[12]}}, instr_i[4:3], instr_i[5], instr_i[2], instr_i[6], 17'h00202, riscv_OpcodeOpImm};
						if ({instr_i[12], instr_i[6:2]} == 6'b000000)
							illegal_instr_o = 1'b1;
					end
					riscv_OpcodeC1MiscAlu:
						case (instr_i[11:10])
							2'b00, 2'b01: instr_o = {1'b0, instr_i[10], 4'b0000, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 5'b10101, instr_i[9:7], riscv_OpcodeOpImm};
							2'b10: instr_o = {{6 {instr_i[12]}}, instr_i[12], instr_i[6:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], riscv_OpcodeOpImm};
							2'b11:
								case ({instr_i[12], instr_i[6:5]})
									3'b000: instr_o = {9'b010000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b00001, instr_i[9:7], riscv_OpcodeOp};
									3'b001: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b10001, instr_i[9:7], riscv_OpcodeOp};
									3'b010: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11001, instr_i[9:7], riscv_OpcodeOp};
									3'b011: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b11101, instr_i[9:7], riscv_OpcodeOp};
									3'b100: instr_o = {9'b010000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b00001, instr_i[9:7], riscv_OpcodeOp32};
									3'b101: instr_o = {9'b000000001, instr_i[4:2], 2'b01, instr_i[9:7], 5'b00001, instr_i[9:7], riscv_OpcodeOp32};
									3'b110, 3'b111: begin
										illegal_instr_o = 1'b1;
										instr_o = {16'b0000000000000000, instr_i};
									end
								endcase
						endcase
					riscv_OpcodeC1J: instr_o = {instr_i[12], instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], {9 {instr_i[12]}}, 4'b0000, ~instr_i[15], riscv_OpcodeJal};
					riscv_OpcodeC1Beqz, riscv_OpcodeC1Bnez: instr_o = {{4 {instr_i[12]}}, instr_i[6:5], instr_i[2], 7'b0000001, instr_i[9:7], 2'b00, instr_i[13], instr_i[11:10], instr_i[4:3], instr_i[12], riscv_OpcodeBranch};
				endcase
			riscv_OpcodeC2:
				case (instr_i[15:13])
					riscv_OpcodeC2Slli: instr_o = {6'b000000, instr_i[12], instr_i[6:2], instr_i[11:7], 3'b001, instr_i[11:7], riscv_OpcodeOpImm};
					riscv_OpcodeC2Fldsp: instr_o = {3'b000, instr_i[4:2], instr_i[12], instr_i[6:5], 11'h013, instr_i[11:7], riscv_OpcodeLoadFp};
					riscv_OpcodeC2Lwsp: begin
						instr_o = {4'b0000, instr_i[3:2], instr_i[12], instr_i[6:4], 10'h012, instr_i[11:7], riscv_OpcodeLoad};
						if (instr_i[11:7] == 5'b00000)
							illegal_instr_o = 1'b1;
					end
					riscv_OpcodeC2Ldsp: begin
						instr_o = {3'b000, instr_i[4:2], instr_i[12], instr_i[6:5], 11'h013, instr_i[11:7], riscv_OpcodeLoad};
						if (instr_i[11:7] == 5'b00000)
							illegal_instr_o = 1'b1;
					end
					riscv_OpcodeC2JalrMvAdd:
						if (instr_i[12] == 1'b0) begin
							instr_o = {7'b0000000, instr_i[6:2], 8'b00000000, instr_i[11:7], riscv_OpcodeOp};
							if (instr_i[6:2] == 5'b00000) begin
								instr_o = {12'b000000000000, instr_i[11:7], 8'b00000000, riscv_OpcodeJalr};
								illegal_instr_o = (instr_i[11:7] != {5 {1'sb0}} ? 1'b0 : 1'b1);
							end
						end
						else begin
							instr_o = {7'b0000000, instr_i[6:2], instr_i[11:7], 3'b000, instr_i[11:7], riscv_OpcodeOp};
							if ((instr_i[11:7] == 5'b00000) && (instr_i[6:2] == 5'b00000))
								instr_o = 32'h00100073;
							else if ((instr_i[11:7] != 5'b00000) && (instr_i[6:2] == 5'b00000))
								instr_o = {12'b000000000000, instr_i[11:7], 8'b00000001, riscv_OpcodeJalr};
						end
					riscv_OpcodeC2Fsdsp: instr_o = {3'b000, instr_i[9:7], instr_i[12], instr_i[6:2], 8'h13, instr_i[11:10], 3'b000, riscv_OpcodeStoreFp};
					riscv_OpcodeC2Swsp: instr_o = {4'b0000, instr_i[8:7], instr_i[12], instr_i[6:2], 8'h12, instr_i[11:9], 2'b00, riscv_OpcodeStore};
					riscv_OpcodeC2Sdsp: instr_o = {3'b000, instr_i[9:7], instr_i[12], instr_i[6:2], 8'h13, instr_i[11:10], 3'b000, riscv_OpcodeStore};
					default: illegal_instr_o = 1'b1;
				endcase
			default: is_compressed_o = 1'b0;
		endcase
		if (illegal_instr_o && is_compressed_o)
			instr_o = instr_i;
	end
endmodule
module controller (
	clk_i,
	rst_ni,
	set_pc_commit_o,
	flush_if_o,
	flush_unissued_instr_o,
	flush_id_o,
	flush_ex_o,
	flush_bp_o,
	flush_icache_o,
	flush_dcache_o,
	flush_dcache_ack_i,
	flush_tlb_o,
	halt_csr_i,
	halt_o,
	eret_i,
	ex_valid_i,
	set_debug_pc_i,
	resolved_branch_i,
	flush_csr_i,
	fence_i_i,
	fence_i,
	sfence_vma_i,
	flush_commit_i
);
	input wire clk_i;
	input wire rst_ni;
	output reg set_pc_commit_o;
	output reg flush_if_o;
	output reg flush_unissued_instr_o;
	output reg flush_id_o;
	output reg flush_ex_o;
	output reg flush_bp_o;
	output reg flush_icache_o;
	output reg flush_dcache_o;
	input wire flush_dcache_ack_i;
	output reg flush_tlb_o;
	input wire halt_csr_i;
	output reg halt_o;
	input wire eret_i;
	input wire ex_valid_i;
	input wire set_debug_pc_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [133:0] resolved_branch_i;
	input wire flush_csr_i;
	input wire fence_i_i;
	input wire fence_i;
	input wire sfence_vma_i;
	input wire flush_commit_i;
	reg fence_active_d;
	reg fence_active_q;
	reg flush_dcache;
	always @(*) begin : flush_ctrl
		fence_active_d = fence_active_q;
		set_pc_commit_o = 1'b0;
		flush_if_o = 1'b0;
		flush_unissued_instr_o = 1'b0;
		flush_id_o = 1'b0;
		flush_ex_o = 1'b0;
		flush_dcache = 1'b0;
		flush_icache_o = 1'b0;
		flush_tlb_o = 1'b0;
		flush_bp_o = 1'b0;
		if (resolved_branch_i[4]) begin
			flush_unissued_instr_o = 1'b1;
			flush_if_o = 1'b1;
		end
		if (fence_i) begin
			set_pc_commit_o = 1'b1;
			flush_if_o = 1'b1;
			flush_unissued_instr_o = 1'b1;
			flush_id_o = 1'b1;
			flush_ex_o = 1'b1;
		end
		if (fence_i_i) begin
			set_pc_commit_o = 1'b1;
			flush_if_o = 1'b1;
			flush_unissued_instr_o = 1'b1;
			flush_id_o = 1'b1;
			flush_ex_o = 1'b1;
			flush_icache_o = 1'b1;
		end
		if (sfence_vma_i) begin
			set_pc_commit_o = 1'b1;
			flush_if_o = 1'b1;
			flush_unissued_instr_o = 1'b1;
			flush_id_o = 1'b1;
			flush_ex_o = 1'b1;
			flush_tlb_o = 1'b1;
		end
		if (flush_csr_i || flush_commit_i) begin
			set_pc_commit_o = 1'b1;
			flush_if_o = 1'b1;
			flush_unissued_instr_o = 1'b1;
			flush_id_o = 1'b1;
			flush_ex_o = 1'b1;
		end
		if ((ex_valid_i || eret_i) || set_debug_pc_i) begin
			set_pc_commit_o = 1'b0;
			flush_if_o = 1'b1;
			flush_unissued_instr_o = 1'b1;
			flush_id_o = 1'b1;
			flush_ex_o = 1'b1;
			flush_bp_o = 1'b1;
		end
	end
	always @(*) halt_o = halt_csr_i || fence_active_q;
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			fence_active_q <= 1'b0;
			flush_dcache_o <= 1'b0;
		end
		else begin
			fence_active_q <= fence_active_d;
			flush_dcache_o <= flush_dcache;
		end
endmodule
module csr_buffer (
	clk_i,
	rst_ni,
	flush_i,
	fu_data_i,
	csr_ready_o,
	csr_valid_i,
	csr_result_o,
	csr_commit_i,
	csr_addr_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	output reg csr_ready_o;
	input wire csr_valid_i;
	output wire [63:0] csr_result_o;
	input wire csr_commit_i;
	output wire [11:0] csr_addr_o;
	reg [12:0] csr_reg_n;
	reg [12:0] csr_reg_q;
	assign csr_result_o = fu_data_i[194-:64];
	assign csr_addr_o = csr_reg_q[12-:12];
	always @(*) begin : write
		csr_reg_n = csr_reg_q;
		csr_ready_o = 1'b1;
		if ((csr_reg_q[0] || csr_valid_i) && ~csr_commit_i)
			csr_ready_o = 1'b0;
		if (csr_valid_i) begin
			csr_reg_n[12-:12] = fu_data_i[78:67];
			csr_reg_n[0] = 1'b1;
		end
		if (csr_commit_i && ~csr_valid_i)
			csr_reg_n[0] = 1'b0;
		if (flush_i)
			csr_reg_n[0] = 1'b0;
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			csr_reg_q <= 13'h0000;
		else
			csr_reg_q <= csr_reg_n;
endmodule
module csr_regfile (
	clk_i,
	rst_ni,
	time_irq_i,
	flush_o,
	halt_csr_o,
	commit_instr_i,
	commit_ack_i,
	boot_addr_i,
	hart_id_i,
	ex_i,
	csr_op_i,
	csr_addr_i,
	csr_wdata_i,
	csr_rdata_o,
	dirty_fp_state_i,
	csr_write_fflags_i,
	pc_i,
	csr_exception_o,
	epc_o,
	eret_o,
	trap_vector_base_o,
	priv_lvl_o,
	fs_o,
	fflags_o,
	frm_o,
	fprec_o,
	irq_ctrl_o,
	en_translation_o,
	en_ld_st_translation_o,
	ld_st_priv_lvl_o,
	sum_o,
	mxr_o,
	satp_ppn_o,
	asid_o,
	irq_i,
	ipi_i,
	debug_req_i,
	set_debug_pc_o,
	tvm_o,
	tw_o,
	tsr_o,
	debug_mode_o,
	single_step_o,
	icache_en_o,
	dcache_en_o,
	perf_addr_o,
	perf_data_o,
	perf_data_i,
	perf_we_o,
	pmpcfg_o,
	pmpaddr_o
);
	parameter [63:0] DmBaseAddress = 64'h0000000000000000;
	parameter signed [31:0] AsidWidth = 1;
	parameter [31:0] NrCommitPorts = 2;
	parameter [31:0] NrPMPEntries = 8;
	input wire clk_i;
	input wire rst_ni;
	input wire time_irq_i;
	output reg flush_o;
	output wire halt_csr_o;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [(NrCommitPorts * 361) - 1:0] commit_instr_i;
	input wire [NrCommitPorts - 1:0] commit_ack_i;
	input wire [63:0] boot_addr_i;
	input wire [63:0] hart_id_i;
	input wire [128:0] ex_i;
	input wire [6:0] csr_op_i;
	input wire [11:0] csr_addr_i;
	input wire [63:0] csr_wdata_i;
	output reg [63:0] csr_rdata_o;
	input wire dirty_fp_state_i;
	input wire csr_write_fflags_i;
	input wire [63:0] pc_i;
	output reg [128:0] csr_exception_o;
	output reg [63:0] epc_o;
	output reg eret_o;
	output reg [63:0] trap_vector_base_o;
	output wire [1:0] priv_lvl_o;
	output wire [1:0] fs_o;
	output wire [4:0] fflags_o;
	output wire [2:0] frm_o;
	output wire [6:0] fprec_o;
	output wire [193:0] irq_ctrl_o;
	output wire en_translation_o;
	output reg en_ld_st_translation_o;
	output reg [1:0] ld_st_priv_lvl_o;
	output wire sum_o;
	output wire mxr_o;
	localparam riscv_PPNW = 44;
	output wire [43:0] satp_ppn_o;
	output wire [AsidWidth - 1:0] asid_o;
	input wire [1:0] irq_i;
	input wire ipi_i;
	input wire debug_req_i;
	output reg set_debug_pc_o;
	output wire tvm_o;
	output wire tw_o;
	output wire tsr_o;
	output wire debug_mode_o;
	output wire single_step_o;
	output wire icache_en_o;
	output wire dcache_en_o;
	output reg [4:0] perf_addr_o;
	output reg [63:0] perf_data_o;
	input wire [63:0] perf_data_i;
	output reg perf_we_o;
	output wire [127:0] pmpcfg_o;
	localparam riscv_PLEN = 56;
	output wire [863:0] pmpaddr_o;
	reg read_access_exception;
	reg update_access_exception;
	reg privilege_violation;
	reg csr_we;
	reg csr_read;
	reg [63:0] csr_wdata;
	reg [63:0] csr_rdata;
	reg [1:0] trap_to_priv_lvl;
	reg en_ld_st_translation_d;
	reg en_ld_st_translation_q;
	wire mprv;
	reg mret;
	reg sret;
	reg dret;
	reg dirty_fp_state_csr;
	reg [63:0] mstatus_q;
	reg [63:0] mstatus_d;
	wire [63:0] mstatus_extended;
	localparam riscv_ASIDW = 16;
	localparam riscv_ModeW = 4;
	reg [63:0] satp_q;
	reg [63:0] satp_d;
	reg [31:0] dcsr_q;
	reg [31:0] dcsr_d;
	wire [11:0] csr_addr;
	reg [1:0] priv_lvl_d;
	reg [1:0] priv_lvl_q;
	reg debug_mode_q;
	reg debug_mode_d;
	reg mtvec_rst_load_q;
	reg [63:0] dpc_q;
	reg [63:0] dpc_d;
	reg [63:0] dscratch0_q;
	reg [63:0] dscratch0_d;
	reg [63:0] dscratch1_q;
	reg [63:0] dscratch1_d;
	reg [63:0] mtvec_q;
	reg [63:0] mtvec_d;
	reg [63:0] medeleg_q;
	reg [63:0] medeleg_d;
	reg [63:0] mideleg_q;
	reg [63:0] mideleg_d;
	reg [63:0] mip_q;
	reg [63:0] mip_d;
	reg [63:0] mie_q;
	reg [63:0] mie_d;
	reg [63:0] mcounteren_q;
	reg [63:0] mcounteren_d;
	reg [63:0] mscratch_q;
	reg [63:0] mscratch_d;
	reg [63:0] mepc_q;
	reg [63:0] mepc_d;
	reg [63:0] mcause_q;
	reg [63:0] mcause_d;
	reg [63:0] mtval_q;
	reg [63:0] mtval_d;
	reg [63:0] stvec_q;
	reg [63:0] stvec_d;
	reg [63:0] scounteren_q;
	reg [63:0] scounteren_d;
	reg [63:0] sscratch_q;
	reg [63:0] sscratch_d;
	reg [63:0] sepc_q;
	reg [63:0] sepc_d;
	reg [63:0] scause_q;
	reg [63:0] scause_d;
	reg [63:0] stval_q;
	reg [63:0] stval_d;
	reg [63:0] dcache_q;
	reg [63:0] dcache_d;
	reg [63:0] icache_q;
	reg [63:0] icache_d;
	reg wfi_d;
	reg wfi_q;
	reg [63:0] cycle_q;
	reg [63:0] cycle_d;
	reg [63:0] instret_q;
	reg [63:0] instret_d;
	reg [127:0] pmpcfg_q;
	reg [127:0] pmpcfg_d;
	reg [863:0] pmpaddr_q;
	reg [863:0] pmpaddr_d;
	assign pmpcfg_o = pmpcfg_q[0+:128];
	assign pmpaddr_o = pmpaddr_q;
	reg [31:0] fcsr_q;
	reg [31:0] fcsr_d;
	assign csr_addr = csr_addr_i;
	assign fs_o = mstatus_q[14-:2];
	localparam riscv_IS_XLEN64 = 1'b1;
	assign mstatus_extended = (riscv_IS_XLEN64 ? mstatus_q[63:0] : {mstatus_q[63], mstatus_q[30:23], mstatus_q[22:0]});
	localparam [63:0] ariane_pkg_ARIANE_MARCHID = {{32 {1'b0}}, 32'd3};
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam [0:0] ariane_pkg_XFVEC = 1'b0;
	localparam [0:0] ariane_pkg_NSX = ((ariane_pkg_XF16 | ariane_pkg_XF16ALT) | ariane_pkg_XF8) | ariane_pkg_XFVEC;
	localparam [0:0] ariane_pkg_RVA = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [63:0] ariane_pkg_ISA_CODE = ((((((((((ariane_pkg_RVA << 0) | 4) | (ariane_pkg_RVD << 3)) | (ariane_pkg_RVF << 5)) | 256) | 4096) | 0) | 262144) | 1048576) | (ariane_pkg_NSX << 23)) | 65'sd9223372036854775808;
	localparam [63:0] riscv_SSTATUS_FS = 'h6000;
	localparam [63:0] riscv_SSTATUS_MXR = 'h80000;
	localparam [63:0] riscv_SSTATUS_SD = {riscv_IS_XLEN64, 31'h00000000, ~riscv_IS_XLEN64, 31'h00000000};
	localparam [63:0] riscv_SSTATUS_SIE = 'h2;
	localparam [63:0] riscv_SSTATUS_SPIE = 'h20;
	localparam [63:0] riscv_SSTATUS_SPP = 'h100;
	localparam [63:0] riscv_SSTATUS_SUM = 'h40000;
	localparam [63:0] riscv_SSTATUS_UIE = 'h1;
	localparam [63:0] riscv_SSTATUS_UPIE = 'h10;
	localparam [63:0] riscv_SSTATUS_UXL = 64'h0000000300000000;
	localparam [63:0] riscv_SSTATUS_XS = 'h18000;
	localparam [63:0] ariane_pkg_SMODE_STATUS_READ_MASK = ((((((((((riscv_SSTATUS_UIE | riscv_SSTATUS_SIE) | riscv_SSTATUS_SPIE) | riscv_SSTATUS_SPP) | riscv_SSTATUS_FS) | riscv_SSTATUS_XS) | riscv_SSTATUS_SUM) | riscv_SSTATUS_MXR) | riscv_SSTATUS_UPIE) | riscv_SSTATUS_SPIE) | riscv_SSTATUS_UXL) | riscv_SSTATUS_SD;
	always @(*) begin : csr_read_process
		read_access_exception = 1'b0;
		csr_rdata = 1'sb0;
		perf_addr_o = csr_addr[4:0];
		if (csr_read)
			case (csr_addr[11-:12])
				12'h001:
					if (mstatus_q[14-:2] == 2'b00)
						read_access_exception = 1'b1;
					else
						csr_rdata = {{59 {1'b0}}, fcsr_q[4-:5]};
				12'h002:
					if (mstatus_q[14-:2] == 2'b00)
						read_access_exception = 1'b1;
					else
						csr_rdata = {{61 {1'b0}}, fcsr_q[7-:3]};
				12'h003:
					if (mstatus_q[14-:2] == 2'b00)
						read_access_exception = 1'b1;
					else
						csr_rdata = {{56 {1'b0}}, fcsr_q[7-:3], fcsr_q[4-:5]};
				12'h800:
					if (mstatus_q[14-:2] == 2'b00)
						read_access_exception = 1'b1;
					else
						csr_rdata = {{57 {1'b0}}, fcsr_q[14-:7]};
				12'h7b0: csr_rdata = {{32 {1'b0}}, dcsr_q};
				12'h7b1: csr_rdata = dpc_q;
				12'h7b2: csr_rdata = dscratch0_q;
				12'h7b3: csr_rdata = dscratch1_q;
				12'h7a0:
					;
				12'h7a1:
					;
				12'h7a2:
					;
				12'h7a3:
					;
				12'h100: csr_rdata = mstatus_extended & ariane_pkg_SMODE_STATUS_READ_MASK[63:0];
				12'h104: csr_rdata = mie_q & mideleg_q;
				12'h144: csr_rdata = mip_q & mideleg_q;
				12'h105: csr_rdata = stvec_q;
				12'h106: csr_rdata = scounteren_q;
				12'h140: csr_rdata = sscratch_q;
				12'h141: csr_rdata = sepc_q;
				12'h142: csr_rdata = scause_q;
				12'h143: csr_rdata = stval_q;
				12'h180:
					if ((priv_lvl_o == 2'b01) && mstatus_q[20])
						read_access_exception = 1'b1;
					else
						csr_rdata = satp_q;
				12'h300: csr_rdata = mstatus_extended;
				12'h301: csr_rdata = ariane_pkg_ISA_CODE;
				12'h302: csr_rdata = medeleg_q;
				12'h303: csr_rdata = mideleg_q;
				12'h304: csr_rdata = mie_q;
				12'h305: csr_rdata = mtvec_q;
				12'h306: csr_rdata = mcounteren_q;
				12'h340: csr_rdata = mscratch_q;
				12'h341: csr_rdata = mepc_q;
				12'h342: csr_rdata = mcause_q;
				12'h343: csr_rdata = mtval_q;
				12'h344: csr_rdata = mip_q;
				12'hf11: csr_rdata = 1'sb0;
				12'hf12: csr_rdata = ariane_pkg_ARIANE_MARCHID;
				12'hf13: csr_rdata = 1'sb0;
				12'hf14: csr_rdata = hart_id_i;
				12'hb00: csr_rdata = cycle_q;
				12'hb02: csr_rdata = instret_q;
				12'hc00: csr_rdata = cycle_q;
				12'hc02: csr_rdata = instret_q;
				12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f: csr_rdata = perf_data_i;
				12'h701: csr_rdata = dcache_q;
				12'h700: csr_rdata = icache_q;
				12'h3a0: csr_rdata = pmpcfg_q[0+:64];
				12'h3a2: csr_rdata = pmpcfg_q[64+:64];
				12'h3b0: csr_rdata = {10'b0000000000, pmpaddr_q[53-:53], (pmpcfg_q[4] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b1: csr_rdata = {10'b0000000000, pmpaddr_q[107-:53], (pmpcfg_q[12] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b2: csr_rdata = {10'b0000000000, pmpaddr_q[161-:53], (pmpcfg_q[20] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b3: csr_rdata = {10'b0000000000, pmpaddr_q[215-:53], (pmpcfg_q[28] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b4: csr_rdata = {10'b0000000000, pmpaddr_q[269-:53], (pmpcfg_q[36] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b5: csr_rdata = {10'b0000000000, pmpaddr_q[323-:53], (pmpcfg_q[44] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b6: csr_rdata = {10'b0000000000, pmpaddr_q[377-:53], (pmpcfg_q[52] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b7: csr_rdata = {10'b0000000000, pmpaddr_q[431-:53], (pmpcfg_q[60] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b8: csr_rdata = {10'b0000000000, pmpaddr_q[485-:53], (pmpcfg_q[68] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3b9: csr_rdata = {10'b0000000000, pmpaddr_q[539-:53], (pmpcfg_q[76] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3ba: csr_rdata = {10'b0000000000, pmpaddr_q[593-:53], (pmpcfg_q[84] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3bb: csr_rdata = {10'b0000000000, pmpaddr_q[647-:53], (pmpcfg_q[92] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3bc: csr_rdata = {10'b0000000000, pmpaddr_q[701-:53], (pmpcfg_q[100] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3bd: csr_rdata = {10'b0000000000, pmpaddr_q[755-:53], (pmpcfg_q[108] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3be: csr_rdata = {10'b0000000000, pmpaddr_q[809-:53], (pmpcfg_q[116] == 1'b1 ? 1'b1 : 1'b0)};
				12'h3bf: csr_rdata = {10'b0000000000, pmpaddr_q[863-:53], (pmpcfg_q[124] == 1'b1 ? 1'b1 : 1'b0)};
				default: read_access_exception = 1'b1;
			endcase
	end
	reg [63:0] mask;
	localparam [0:0] ariane_pkg_ENABLE_CYCLE_COUNT = 1'b1;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	localparam [63:0] ariane_pkg_SMODE_STATUS_WRITE_MASK = ((((riscv_SSTATUS_SIE | riscv_SSTATUS_SPIE) | riscv_SSTATUS_SPP) | riscv_SSTATUS_FS) | riscv_SSTATUS_SUM) | riscv_SSTATUS_MXR;
	localparam [0:0] ariane_pkg_ZERO_TVAL = 1'b0;
	localparam [2:0] dm_CauseBreakpoint = 3'h1;
	localparam [2:0] dm_CauseRequest = 3'h3;
	localparam [2:0] dm_CauseSingleStep = 3'h4;
	localparam [63:0] riscv_BREAKPOINT = 3;
	localparam [63:0] riscv_DEBUG_REQUEST = 24;
	localparam [63:0] riscv_ENV_CALL_MMODE = 11;
	localparam [63:0] riscv_ENV_CALL_SMODE = 9;
	localparam [63:0] riscv_ENV_CALL_UMODE = 8;
	localparam [63:0] riscv_ILLEGAL_INSTR = 2;
	localparam [63:0] riscv_INSTR_ADDR_MISALIGNED = 0;
	localparam [63:0] riscv_INSTR_PAGE_FAULT = 12;
	localparam [31:0] riscv_IRQ_M_EXT = 11;
	localparam [31:0] riscv_IRQ_M_SOFT = 3;
	localparam [31:0] riscv_IRQ_M_TIMER = 7;
	localparam [63:0] riscv_LOAD_PAGE_FAULT = 13;
	localparam [63:0] riscv_MIP_MEIP = 2048;
	localparam [63:0] riscv_MIP_MSIP = 8;
	localparam [63:0] riscv_MIP_MTIP = 128;
	localparam [31:0] riscv_IRQ_S_EXT = 9;
	localparam [63:0] riscv_MIP_SEIP = 512;
	localparam [31:0] riscv_IRQ_S_SOFT = 1;
	localparam [63:0] riscv_MIP_SSIP = 2;
	localparam [31:0] riscv_IRQ_S_TIMER = 5;
	localparam [63:0] riscv_MIP_STIP = 32;
	localparam [3:0] riscv_MODE_SV = 4'd8;
	localparam [63:0] riscv_STORE_PAGE_FAULT = 15;
	function automatic [63:0] sv2v_cast_3DFE6;
		input reg [63:0] inp;
		sv2v_cast_3DFE6 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	always @(*) begin : csr_update
		reg [63:0] satp;
		reg [63:0] instret;
		satp = satp_q;
		instret = instret_q;
		cycle_d = cycle_q;
		instret_d = instret_q;
		if (!debug_mode_q) begin
			begin : sv2v_autoblock_1
				reg signed [31:0] i;
				for (i = 0; i < NrCommitPorts; i = i + 1)
					if (commit_ack_i[i] && !ex_i[0])
						instret = instret + 1;
			end
			instret_d = instret;
			if (ariane_pkg_ENABLE_CYCLE_COUNT)
				cycle_d = cycle_q + 1'b1;
			else
				cycle_d = instret;
		end
		eret_o = 1'b0;
		flush_o = 1'b0;
		update_access_exception = 1'b0;
		set_debug_pc_o = 1'b0;
		perf_we_o = 1'b0;
		perf_data_o = 'b0;
		fcsr_d = fcsr_q;
		priv_lvl_d = priv_lvl_q;
		debug_mode_d = debug_mode_q;
		dcsr_d = dcsr_q;
		dpc_d = dpc_q;
		dscratch0_d = dscratch0_q;
		dscratch1_d = dscratch1_q;
		mstatus_d = mstatus_q;
		if (mtvec_rst_load_q)
			mtvec_d = {boot_addr_i} + 'h40;
		else
			mtvec_d = mtvec_q;
		medeleg_d = medeleg_q;
		mideleg_d = mideleg_q;
		mip_d = mip_q;
		mie_d = mie_q;
		mepc_d = mepc_q;
		mcause_d = mcause_q;
		mcounteren_d = mcounteren_q;
		mscratch_d = mscratch_q;
		mtval_d = mtval_q;
		dcache_d = dcache_q;
		icache_d = icache_q;
		sepc_d = sepc_q;
		scause_d = scause_q;
		stvec_d = stvec_q;
		scounteren_d = scounteren_q;
		sscratch_d = sscratch_q;
		stval_d = stval_q;
		satp_d = satp_q;
		en_ld_st_translation_d = en_ld_st_translation_q;
		dirty_fp_state_csr = 1'b0;
		pmpcfg_d = pmpcfg_q;
		pmpaddr_d = pmpaddr_q;
		if (csr_we)
			case (csr_addr[11-:12])
				12'h001:
					if (mstatus_q[14-:2] == 2'b00)
						update_access_exception = 1'b1;
					else begin
						dirty_fp_state_csr = 1'b1;
						fcsr_d[4-:5] = csr_wdata[4:0];
						flush_o = 1'b1;
					end
				12'h002:
					if (mstatus_q[14-:2] == 2'b00)
						update_access_exception = 1'b1;
					else begin
						dirty_fp_state_csr = 1'b1;
						fcsr_d[7-:3] = csr_wdata[2:0];
						flush_o = 1'b1;
					end
				12'h003:
					if (mstatus_q[14-:2] == 2'b00)
						update_access_exception = 1'b1;
					else begin
						dirty_fp_state_csr = 1'b1;
						fcsr_d[7:0] = csr_wdata[7:0];
						flush_o = 1'b1;
					end
				12'h800:
					if (mstatus_q[14-:2] == 2'b00)
						update_access_exception = 1'b1;
					else begin
						dirty_fp_state_csr = 1'b1;
						fcsr_d[14-:7] = csr_wdata[6:0];
						flush_o = 1'b1;
					end
				12'h7b0: begin
					dcsr_d = csr_wdata[31:0];
					dcsr_d[31-:4] = 4'h4;
					dcsr_d[3] = 1'b0;
					dcsr_d[10] = 1'b0;
					dcsr_d[9] = 1'b0;
				end
				12'h7b1: dpc_d = csr_wdata;
				12'h7b2: dscratch0_d = csr_wdata;
				12'h7b3: dscratch1_d = csr_wdata;
				12'h7a0:
					;
				12'h7a1:
					;
				12'h7a2:
					;
				12'h7a3:
					;
				12'h100: begin
					mask = ariane_pkg_SMODE_STATUS_WRITE_MASK[63:0];
					mstatus_d = (mstatus_q & ~{mask}) | {csr_wdata & mask};
					if (!ariane_pkg_FP_PRESENT)
						mstatus_d[14-:2] = 2'b00;
					flush_o = 1'b1;
				end
				12'h104: mie_d = (mie_q & ~mideleg_q) | (csr_wdata & mideleg_q);
				12'h144: begin
					mask = riscv_MIP_SSIP & mideleg_q;
					mip_d = (mip_q & ~mask) | (csr_wdata & mask);
				end
				12'h105: stvec_d = {csr_wdata[63:2], 1'b0, csr_wdata[0]};
				12'h106: scounteren_d = {{32 {1'b0}}, csr_wdata[31:0]};
				12'h140: sscratch_d = csr_wdata;
				12'h141: sepc_d = {csr_wdata[63:1], 1'b0};
				12'h142: scause_d = csr_wdata;
				12'h143: stval_d = csr_wdata;
				12'h180: begin
					if ((priv_lvl_o == 2'b01) && mstatus_q[20])
						update_access_exception = 1'b1;
					else begin
						satp = sv2v_cast_3DFE6(csr_wdata);
						satp[59-:16] = satp[59-:16] & {{riscv_ASIDW - AsidWidth {1'b0}}, {AsidWidth {1'b1}}};
						if ((sv2v_cast_4(satp[63-:4]) == 4'd0) || (sv2v_cast_4(satp[63-:4]) == riscv_MODE_SV))
							satp_d = satp;
					end
					flush_o = 1'b1;
				end
				12'h300: begin
					mstatus_d = {csr_wdata};
					mstatus_d[16-:2] = 2'b00;
					if (!ariane_pkg_FP_PRESENT)
						mstatus_d[14-:2] = 2'b00;
					mstatus_d[4] = 1'b0;
					mstatus_d[0] = 1'b0;
					flush_o = 1'b1;
				end
				12'h301:
					;
				12'h302: begin
					mask = 45321;
					medeleg_d = (medeleg_q & ~mask) | (csr_wdata & mask);
				end
				12'h303: begin
					mask = (riscv_MIP_SSIP | riscv_MIP_STIP) | riscv_MIP_SEIP;
					mideleg_d = (mideleg_q & ~mask) | (csr_wdata & mask);
				end
				12'h304: begin
					mask = ((((riscv_MIP_SSIP | riscv_MIP_STIP) | riscv_MIP_SEIP) | riscv_MIP_MSIP) | riscv_MIP_MTIP) | riscv_MIP_MEIP;
					mie_d = (mie_q & ~mask) | (csr_wdata & mask);
				end
				12'h305: begin
					mtvec_d = {csr_wdata[63:2], 1'b0, csr_wdata[0]};
					if (csr_wdata[0])
						mtvec_d = {csr_wdata[63:8], 7'b0000000, csr_wdata[0]};
				end
				12'h306: mcounteren_d = {{32 {1'b0}}, csr_wdata[31:0]};
				12'h340: mscratch_d = csr_wdata;
				12'h341: mepc_d = {csr_wdata[63:1], 1'b0};
				12'h342: mcause_d = csr_wdata;
				12'h343: mtval_d = csr_wdata;
				12'h344: begin
					mask = (riscv_MIP_SSIP | riscv_MIP_STIP) | riscv_MIP_SEIP;
					mip_d = (mip_q & ~mask) | (csr_wdata & mask);
				end
				12'hb00: cycle_d = csr_wdata;
				12'hb02: instret = csr_wdata;
				12'hb03, 12'hb04, 12'hb05, 12'hb06, 12'hb07, 12'hb08, 12'hb09, 12'hb0a, 12'hb0b, 12'hb0c, 12'hb0d, 12'hb0e, 12'hb0f, 12'hb10, 12'hb11, 12'hb12, 12'hb13, 12'hb14, 12'hb15, 12'hb16, 12'hb17, 12'hb18, 12'hb19, 12'hb1a, 12'hb1b, 12'hb1c, 12'hb1d, 12'hb1e, 12'hb1f: begin
					perf_data_o = csr_wdata;
					perf_we_o = 1'b1;
				end
				12'h701: dcache_d = {{63 {1'b0}}, csr_wdata[0]};
				12'h700: icache_d = {{63 {1'b0}}, csr_wdata[0]};
				12'h3a0: begin : sv2v_autoblock_2
					reg signed [31:0] i;
					for (i = 0; i < 8; i = i + 1)
						if (!pmpcfg_q[(i * 8) + 7])
							pmpcfg_d[i * 8+:8] = csr_wdata[i * 8+:8];
				end
				12'h3a1:
					;
				12'h3a2: begin : sv2v_autoblock_3
					reg signed [31:0] i;
					for (i = 0; i < 8; i = i + 1)
						if (!pmpcfg_q[((i + 8) * 8) + 7])
							pmpcfg_d[(i + 8) * 8+:8] = csr_wdata[i * 8+:8];
				end
				12'h3a3:
					;
				12'h3b0:
					if (!pmpcfg_q[7] && !(pmpcfg_q[15] && (pmpcfg_q[12-:2] == 2'b01)))
						pmpaddr_d[0+:54] = csr_wdata[53:0];
				12'h3b1:
					if (!pmpcfg_q[15] && !(pmpcfg_q[23] && (pmpcfg_q[20-:2] == 2'b01)))
						pmpaddr_d[54+:54] = csr_wdata[53:0];
				12'h3b2:
					if (!pmpcfg_q[23] && !(pmpcfg_q[31] && (pmpcfg_q[28-:2] == 2'b01)))
						pmpaddr_d[108+:54] = csr_wdata[53:0];
				12'h3b3:
					if (!pmpcfg_q[31] && !(pmpcfg_q[39] && (pmpcfg_q[36-:2] == 2'b01)))
						pmpaddr_d[162+:54] = csr_wdata[53:0];
				12'h3b4:
					if (!pmpcfg_q[39] && !(pmpcfg_q[47] && (pmpcfg_q[44-:2] == 2'b01)))
						pmpaddr_d[216+:54] = csr_wdata[53:0];
				12'h3b5:
					if (!pmpcfg_q[47] && !(pmpcfg_q[55] && (pmpcfg_q[52-:2] == 2'b01)))
						pmpaddr_d[270+:54] = csr_wdata[53:0];
				12'h3b6:
					if (!pmpcfg_q[55] && !(pmpcfg_q[63] && (pmpcfg_q[60-:2] == 2'b01)))
						pmpaddr_d[324+:54] = csr_wdata[53:0];
				12'h3b7:
					if (!pmpcfg_q[63] && !(pmpcfg_q[71] && (pmpcfg_q[68-:2] == 2'b01)))
						pmpaddr_d[378+:54] = csr_wdata[53:0];
				12'h3b8:
					if (!pmpcfg_q[71] && !(pmpcfg_q[79] && (pmpcfg_q[76-:2] == 2'b01)))
						pmpaddr_d[432+:54] = csr_wdata[53:0];
				12'h3b9:
					if (!pmpcfg_q[79] && !(pmpcfg_q[87] && (pmpcfg_q[84-:2] == 2'b01)))
						pmpaddr_d[486+:54] = csr_wdata[53:0];
				12'h3ba:
					if (!pmpcfg_q[87] && !(pmpcfg_q[95] && (pmpcfg_q[92-:2] == 2'b01)))
						pmpaddr_d[540+:54] = csr_wdata[53:0];
				12'h3bb:
					if (!pmpcfg_q[95] && !(pmpcfg_q[103] && (pmpcfg_q[100-:2] == 2'b01)))
						pmpaddr_d[594+:54] = csr_wdata[53:0];
				12'h3bc:
					if (!pmpcfg_q[103] && !(pmpcfg_q[111] && (pmpcfg_q[108-:2] == 2'b01)))
						pmpaddr_d[648+:54] = csr_wdata[53:0];
				12'h3bd:
					if (!pmpcfg_q[111] && !(pmpcfg_q[119] && (pmpcfg_q[116-:2] == 2'b01)))
						pmpaddr_d[702+:54] = csr_wdata[53:0];
				12'h3be:
					if (!pmpcfg_q[119] && !(pmpcfg_q[127] && (pmpcfg_q[124-:2] == 2'b01)))
						pmpaddr_d[756+:54] = csr_wdata[53:0];
				12'h3bf:
					if (!pmpcfg_q[127])
						pmpaddr_d[810+:54] = csr_wdata[53:0];
				default: update_access_exception = 1'b1;
			endcase
		mstatus_d[35-:2] = 2'b10;
		mstatus_d[33-:2] = 2'b10;
		if (ariane_pkg_FP_PRESENT && (dirty_fp_state_csr || dirty_fp_state_i))
			mstatus_d[14-:2] = 2'b11;
		mstatus_d[63] = (mstatus_q[16-:2] == 2'b11) | (mstatus_q[14-:2] == 2'b11);
		if (csr_write_fflags_i)
			fcsr_d[4-:5] = csr_wdata_i[4:0] | fcsr_q[4-:5];
		mip_d[riscv_IRQ_M_EXT] = irq_i[0];
		mip_d[riscv_IRQ_M_SOFT] = ipi_i;
		mip_d[riscv_IRQ_M_TIMER] = time_irq_i;
		trap_to_priv_lvl = 2'b11;
		if ((!debug_mode_q && (ex_i[128-:64] != riscv_DEBUG_REQUEST)) && ex_i[0]) begin
			flush_o = 1'b0;
			if ((ex_i[128] && mideleg_q[ex_i[70:65]]) || (~ex_i[128] && medeleg_q[ex_i[70:65]]))
				trap_to_priv_lvl = (priv_lvl_o == 2'b11 ? 2'b11 : 2'b01);
			if (trap_to_priv_lvl == 2'b01) begin
				mstatus_d[1] = 1'b0;
				mstatus_d[5] = mstatus_q[1];
				mstatus_d[8] = priv_lvl_q[0];
				scause_d = ex_i[128-:64];
				sepc_d = {pc_i};
				stval_d = (1'b0 && (|{ex_i[128-:64] == 64'd2, ex_i[128-:64] == 64'd3, ex_i[128-:64] == 64'd8, ex_i[128-:64] == 64'd9, ex_i[128-:64] == 64'd11} || ex_i[128]) ? {64 {1'sb0}} : ex_i[64-:64]);
			end
			else begin
				mstatus_d[3] = 1'b0;
				mstatus_d[7] = mstatus_q[3];
				mstatus_d[12-:2] = priv_lvl_q;
				mcause_d = ex_i[128-:64];
				mepc_d = {pc_i};
				mtval_d = (1'b0 && (|{ex_i[128-:64] == 64'd2, ex_i[128-:64] == 64'd3, ex_i[128-:64] == 64'd8, ex_i[128-:64] == 64'd9, ex_i[128-:64] == 64'd11} || ex_i[128]) ? {64 {1'sb0}} : ex_i[64-:64]);
			end
			priv_lvl_d = trap_to_priv_lvl;
		end
		if (!debug_mode_q) begin
			dcsr_d[1-:2] = priv_lvl_o;
			if (ex_i[0] && (ex_i[128-:64] == riscv_BREAKPOINT)) begin
				dcsr_d[1-:2] = priv_lvl_o;
				case (priv_lvl_o)
					2'b11: begin
						debug_mode_d = dcsr_q[15];
						set_debug_pc_o = dcsr_q[15];
					end
					2'b01: begin
						debug_mode_d = dcsr_q[13];
						set_debug_pc_o = dcsr_q[13];
					end
					2'b00: begin
						debug_mode_d = dcsr_q[12];
						set_debug_pc_o = dcsr_q[12];
					end
					default:
						;
				endcase
				dpc_d = {pc_i};
				dcsr_d[8-:3] = dm_CauseBreakpoint;
			end
			if (ex_i[0] && (ex_i[128-:64] == riscv_DEBUG_REQUEST)) begin
				dcsr_d[1-:2] = priv_lvl_o;
				dpc_d = {pc_i};
				debug_mode_d = 1'b1;
				set_debug_pc_o = 1'b1;
				dcsr_d[8-:3] = dm_CauseRequest;
			end
			if (dcsr_q[2] && commit_ack_i[0]) begin
				dcsr_d[1-:2] = priv_lvl_o;
				if (commit_instr_i[293-:4] == 4'd4)
					dpc_d = {commit_instr_i[64-:riscv_VLEN]};
				else if (ex_i[0])
					dpc_d = {trap_vector_base_o};
				else if (eret_o)
					dpc_d = {epc_o};
				else
					dpc_d = {commit_instr_i[360-:64] + (commit_instr_i[0] ? 'h2 : 'h4)};
				debug_mode_d = 1'b1;
				set_debug_pc_o = 1'b1;
				dcsr_d[8-:3] = dm_CauseSingleStep;
			end
		end
		if ((debug_mode_q && ex_i[0]) && (ex_i[128-:64] == riscv_BREAKPOINT))
			set_debug_pc_o = 1'b1;
		if ((mprv && (sv2v_cast_4(satp_q[63-:4]) == riscv_MODE_SV)) && (mstatus_q[12-:2] != 2'b11))
			en_ld_st_translation_d = 1'b1;
		else
			en_ld_st_translation_d = en_translation_o;
		ld_st_priv_lvl_o = (mprv ? mstatus_q[12-:2] : priv_lvl_o);
		en_ld_st_translation_o = en_ld_st_translation_q;
		if (mret) begin
			eret_o = 1'b1;
			mstatus_d[3] = mstatus_q[7];
			priv_lvl_d = mstatus_q[12-:2];
			mstatus_d[12-:2] = 2'b00;
			mstatus_d[7] = 1'b1;
		end
		if (sret) begin
			eret_o = 1'b1;
			mstatus_d[1] = mstatus_q[5];
			priv_lvl_d = sv2v_cast_2({1'b0, mstatus_q[8]});
			mstatus_d[8] = 1'b0;
			mstatus_d[5] = 1'b1;
		end
		if (dret) begin
			eret_o = 1'b1;
			priv_lvl_d = sv2v_cast_2(dcsr_q[1-:2]);
			debug_mode_d = 1'b0;
		end
	end
	always @(*) begin : csr_op_logic
		csr_wdata = csr_wdata_i;
		csr_we = 1'b1;
		csr_read = 1'b1;
		mret = 1'b0;
		sret = 1'b0;
		dret = 1'b0;
		case (csr_op_i)
			7'd31: csr_wdata = csr_wdata_i;
			7'd33: csr_wdata = csr_wdata_i | csr_rdata;
			7'd34: csr_wdata = ~csr_wdata_i & csr_rdata;
			7'd32: csr_we = 1'b0;
			7'd24: begin
				csr_we = 1'b0;
				csr_read = 1'b0;
				sret = 1'b1;
			end
			7'd23: begin
				csr_we = 1'b0;
				csr_read = 1'b0;
				mret = 1'b1;
			end
			7'd25: begin
				csr_we = 1'b0;
				csr_read = 1'b0;
				dret = 1'b1;
			end
			default: begin
				csr_we = 1'b0;
				csr_read = 1'b0;
			end
		endcase
		if (privilege_violation) begin
			csr_we = 1'b0;
			csr_read = 1'b0;
		end
	end
	assign irq_ctrl_o[193-:64] = mie_q;
	assign irq_ctrl_o[129-:64] = mip_q;
	assign irq_ctrl_o[1] = mstatus_q[1];
	assign irq_ctrl_o[65-:64] = mideleg_q;
	assign irq_ctrl_o[0] = (~debug_mode_q & (~dcsr_q[2] | dcsr_q[11])) & ((mstatus_q[3] & (priv_lvl_o == 2'b11)) | (priv_lvl_o != 2'b11));
	always @(*) begin : privilege_check
		privilege_violation = 1'b0;
		if (|{csr_op_i == 7'd31, csr_op_i == 7'd33, csr_op_i == 7'd34, csr_op_i == 7'd32}) begin
			if (sv2v_cast_2(priv_lvl_o & csr_addr[9-:2]) != csr_addr[9-:2])
				privilege_violation = 1'b1;
			if ((csr_addr_i[11:4] == 8'h7b) && !debug_mode_q)
				privilege_violation = 1'b1;
			if ((12'hc00 <= csr_addr_i) && (12'hc1f >= csr_addr_i))
				case (csr_addr[9-:2])
					2'b11: privilege_violation = 1'b0;
					2'b01: privilege_violation = ~mcounteren_q[csr_addr_i[4:0]];
					2'b00: privilege_violation = ~mcounteren_q[csr_addr_i[4:0]] & ~scounteren_q[csr_addr_i[4:0]];
				endcase
		end
	end
	always @(*) begin : exception_ctrl
		csr_exception_o = 3'b000;
		if (update_access_exception || read_access_exception) begin
			csr_exception_o[128-:64] = riscv_ILLEGAL_INSTR;
			csr_exception_o[0] = 1'b1;
		end
		if (privilege_violation) begin
			csr_exception_o[128-:64] = riscv_ILLEGAL_INSTR;
			csr_exception_o[0] = 1'b1;
		end
	end
	always @(*) begin : wfi_ctrl
		wfi_d = wfi_q;
		if ((|mip_q || debug_req_i) || irq_i[1])
			wfi_d = 1'b0;
		else if ((!debug_mode_q && (csr_op_i == 7'd27)) && !ex_i[0])
			wfi_d = 1'b1;
	end
	localparam [63:0] dm_HaltAddress = 64'h0000000000000800;
	localparam [63:0] dm_ExceptionAddress = 2056;
	always @(*) begin : priv_output
		trap_vector_base_o = {mtvec_q[63:2], 2'b00};
		if (trap_to_priv_lvl == 2'b01)
			trap_vector_base_o = {stvec_q[63:2], 2'b00};
		if (debug_mode_q)
			trap_vector_base_o = DmBaseAddress[63:0] + dm_ExceptionAddress[63:0];
		if ((mtvec_q[0] || stvec_q[0]) && ex_i[128])
			trap_vector_base_o[7:2] = ex_i[70:65];
		epc_o = mepc_q[63:0];
		if (sret)
			epc_o = sepc_q[63:0];
		if (dret)
			epc_o = dpc_q[63:0];
	end
	always @(*) begin
		csr_rdata_o = csr_rdata;
		case (csr_addr[11-:12])
			12'h344: csr_rdata_o = csr_rdata | (irq_i[1] << riscv_IRQ_S_EXT);
			12'h144: csr_rdata_o = csr_rdata | ((irq_i[1] & mideleg_q[riscv_IRQ_S_EXT]) << riscv_IRQ_S_EXT);
			default:
				;
		endcase
	end
	assign priv_lvl_o = (debug_mode_q ? 2'b11 : priv_lvl_q);
	assign fflags_o = fcsr_q[4-:5];
	assign frm_o = fcsr_q[7-:3];
	assign fprec_o = fcsr_q[14-:7];
	assign satp_ppn_o = satp_q[43-:riscv_PPNW];
	assign asid_o = satp_q[43 + AsidWidth:44];
	assign sum_o = mstatus_q[18];
	assign en_translation_o = ((sv2v_cast_4(satp_q[63-:4]) == riscv_MODE_SV) && (priv_lvl_o != 2'b11) ? 1'b1 : 1'b0);
	assign mxr_o = mstatus_q[19];
	assign tvm_o = mstatus_q[20];
	assign tw_o = mstatus_q[21];
	assign tsr_o = mstatus_q[22];
	assign halt_csr_o = wfi_q;
	assign icache_en_o = icache_q[0] & ~debug_mode_q;
	assign dcache_en_o = dcache_q[0];
	assign mprv = (debug_mode_q && !dcsr_q[4] ? 1'b0 : mstatus_q[17]);
	assign debug_mode_o = debug_mode_q;
	assign single_step_o = dcsr_q[2];
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			priv_lvl_q <= 2'b11;
			fcsr_q <= 1'sb0;
			debug_mode_q <= 1'b0;
			dcsr_q <= 1'sb0;
			dcsr_q[1-:2] <= 2'b11;
			dpc_q <= 1'sb0;
			dscratch0_q <= {riscv_XLEN {1'b0}};
			dscratch1_q <= {riscv_XLEN {1'b0}};
			mstatus_q <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
			mtvec_rst_load_q <= 1'b1;
			mtvec_q <= 1'sb0;
			medeleg_q <= {riscv_XLEN {1'b0}};
			mideleg_q <= {riscv_XLEN {1'b0}};
			mip_q <= {riscv_XLEN {1'b0}};
			mie_q <= {riscv_XLEN {1'b0}};
			mepc_q <= {riscv_XLEN {1'b0}};
			mcause_q <= {riscv_XLEN {1'b0}};
			mcounteren_q <= {riscv_XLEN {1'b0}};
			mscratch_q <= {riscv_XLEN {1'b0}};
			mtval_q <= {riscv_XLEN {1'b0}};
			dcache_q <= {{63 {1'b0}}, 1'b1};
			icache_q <= {{63 {1'b0}}, 1'b1};
			sepc_q <= {riscv_XLEN {1'b0}};
			scause_q <= {riscv_XLEN {1'b0}};
			stvec_q <= {riscv_XLEN {1'b0}};
			scounteren_q <= {riscv_XLEN {1'b0}};
			sscratch_q <= {riscv_XLEN {1'b0}};
			stval_q <= {riscv_XLEN {1'b0}};
			satp_q <= {riscv_XLEN {1'b0}};
			cycle_q <= {riscv_XLEN {1'b0}};
			instret_q <= {riscv_XLEN {1'b0}};
			en_ld_st_translation_q <= 1'b0;
			wfi_q <= 1'b0;
			pmpcfg_q <= 1'sb0;
			pmpaddr_q <= 1'sb0;
		end
		else begin
			priv_lvl_q <= priv_lvl_d;
			fcsr_q <= fcsr_d;
			debug_mode_q <= debug_mode_d;
			dcsr_q <= dcsr_d;
			dpc_q <= dpc_d;
			dscratch0_q <= dscratch0_d;
			dscratch1_q <= dscratch1_d;
			mstatus_q <= mstatus_d;
			mtvec_rst_load_q <= 1'b0;
			mtvec_q <= mtvec_d;
			medeleg_q <= medeleg_d;
			mideleg_q <= mideleg_d;
			mip_q <= mip_d;
			mie_q <= mie_d;
			mepc_q <= mepc_d;
			mcause_q <= mcause_d;
			mcounteren_q <= mcounteren_d;
			mscratch_q <= mscratch_d;
			mtval_q <= mtval_d;
			dcache_q <= dcache_d;
			icache_q <= icache_d;
			sepc_q <= sepc_d;
			scause_q <= scause_d;
			stvec_q <= stvec_d;
			scounteren_q <= scounteren_d;
			sscratch_q <= sscratch_d;
			stval_q <= stval_d;
			satp_q <= satp_d;
			cycle_q <= cycle_d;
			instret_q <= instret_d;
			en_ld_st_translation_q <= en_ld_st_translation_d;
			wfi_q <= wfi_d;
			begin : sv2v_autoblock_4
				reg signed [31:0] i;
				for (i = 0; i < 16; i = i + 1)
					if (i < NrPMPEntries) begin
						pmpcfg_q[i * 8+:8] <= pmpcfg_d[i * 8+:8];
						pmpaddr_q[i * 54+:54] <= pmpaddr_d[i * 54+:54];
					end
					else begin
						pmpcfg_q[i * 8+:8] <= 1'sb0;
						pmpaddr_q[i * 54+:54] <= 1'sb0;
					end
			end
		end
endmodule
module decoder (
	debug_req_i,
	pc_i,
	is_compressed_i,
	compressed_instr_i,
	is_illegal_i,
	instruction_i,
	branch_predict_i,
	ex_i,
	irq_i,
	irq_ctrl_i,
	priv_lvl_i,
	debug_mode_i,
	fs_i,
	frm_i,
	tvm_i,
	tw_i,
	tsr_i,
	instruction_o,
	is_control_flow_instr_o
);
	input wire debug_req_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] pc_i;
	input wire is_compressed_i;
	input wire [15:0] compressed_instr_i;
	input wire is_illegal_i;
	input wire [31:0] instruction_i;
	input wire [66:0] branch_predict_i;
	input wire [128:0] ex_i;
	input wire [1:0] irq_i;
	input wire [193:0] irq_ctrl_i;
	input wire [1:0] priv_lvl_i;
	input wire debug_mode_i;
	input wire [1:0] fs_i;
	input wire [2:0] frm_i;
	input wire tvm_i;
	input wire tw_i;
	input wire tsr_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	output reg [360:0] instruction_o;
	output reg is_control_flow_instr_o;
	reg illegal_instr;
	reg ecall;
	reg ebreak;
	reg check_fprm;
	wire [31:0] instr;
	assign instr = instruction_i;
	reg [3:0] imm_select;
	reg [63:0] imm_i_type;
	reg [63:0] imm_s_type;
	reg [63:0] imm_sb_type;
	reg [63:0] imm_u_type;
	reg [63:0] imm_uj_type;
	reg [63:0] imm_bi_type;
	localparam [0:0] ariane_pkg_ENABLE_WFI = 1'b1;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	localparam [0:0] ariane_pkg_RVA = 1'b1;
	localparam ariane_pkg_FLEN = (ariane_pkg_RVD ? 64 : (ariane_pkg_RVF ? 32 : (ariane_pkg_XF16 ? 16 : (ariane_pkg_XF16ALT ? 16 : (ariane_pkg_XF8 ? 8 : 1)))));
	localparam [0:0] ariane_pkg_XFVEC = 1'b0;
	localparam [0:0] ariane_pkg_RVFVEC = (ariane_pkg_RVF & ariane_pkg_XFVEC) & (ariane_pkg_FLEN > 32);
	localparam [0:0] ariane_pkg_XF16ALTVEC = (ariane_pkg_XF16ALT & ariane_pkg_XFVEC) & (ariane_pkg_FLEN > 16);
	localparam [0:0] ariane_pkg_XF16VEC = (ariane_pkg_XF16 & ariane_pkg_XFVEC) & (ariane_pkg_FLEN > 16);
	localparam [0:0] ariane_pkg_XF8VEC = (ariane_pkg_XF8 & ariane_pkg_XFVEC) & (ariane_pkg_FLEN > 8);
	localparam riscv_OpcodeAmo = 7'b0101111;
	localparam riscv_OpcodeAuipc = 7'b0010111;
	localparam riscv_OpcodeBranch = 7'b1100011;
	localparam riscv_OpcodeJal = 7'b1101111;
	localparam riscv_OpcodeJalr = 7'b1100111;
	localparam riscv_OpcodeLoad = 7'b0000011;
	localparam riscv_OpcodeLoadFp = 7'b0000111;
	localparam riscv_OpcodeLui = 7'b0110111;
	localparam riscv_OpcodeMadd = 7'b1000011;
	localparam riscv_OpcodeMiscMem = 7'b0001111;
	localparam riscv_OpcodeMsub = 7'b1000111;
	localparam riscv_OpcodeNmadd = 7'b1001111;
	localparam riscv_OpcodeNmsub = 7'b1001011;
	localparam riscv_OpcodeOp = 7'b0110011;
	localparam riscv_OpcodeOp32 = 7'b0111011;
	localparam riscv_OpcodeOpFp = 7'b1010011;
	localparam riscv_OpcodeOpImm = 7'b0010011;
	localparam riscv_OpcodeOpImm32 = 7'b0011011;
	localparam riscv_OpcodeStore = 7'b0100011;
	localparam riscv_OpcodeStoreFp = 7'b0100111;
	localparam riscv_OpcodeSystem = 7'b1110011;
	always @(*) begin : decoder
		imm_select = 4'd0;
		is_control_flow_instr_o = 1'b0;
		illegal_instr = 1'b0;
		instruction_o[360-:64] = pc_i;
		instruction_o[296-:3] = 5'b00000;
		instruction_o[293-:4] = 4'd0;
		instruction_o[289-:7] = 7'd0;
		instruction_o[282-:6] = 1'sb0;
		instruction_o[276-:6] = 1'sb0;
		instruction_o[270-:6] = 1'sb0;
		instruction_o[197] = 1'b0;
		instruction_o[296-:3] = 1'sb0;
		instruction_o[0] = is_compressed_i;
		instruction_o[198] = 1'b0;
		instruction_o[67-:67] = branch_predict_i;
		ecall = 1'b0;
		ebreak = 1'b0;
		check_fprm = 1'b0;
		if (~ex_i[0])
			case (instr[6-:7])
				riscv_OpcodeSystem: begin
					instruction_o[293-:4] = 4'd6;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[275:271] = instr[24-:5];
					instruction_o[269:265] = instr[11-:5];
					case (instr[14-:3])
						3'b000: begin
							if ((instr[19-:5] != {5 {1'sb0}}) || (instr[11-:5] != {5 {1'sb0}}))
								illegal_instr = 1'b1;
							case (instr[31-:12])
								12'b000000000000: ecall = 1'b1;
								12'b000000000001: ebreak = 1'b1;
								12'b000100000010: begin
									instruction_o[289-:7] = 7'd24;
									if (priv_lvl_i == 2'b00) begin
										illegal_instr = 1'b1;
										instruction_o[289-:7] = 7'd0;
									end
									if ((priv_lvl_i == 2'b01) && tsr_i) begin
										illegal_instr = 1'b1;
										instruction_o[289-:7] = 7'd0;
									end
								end
								12'b001100000010: begin
									instruction_o[289-:7] = 7'd23;
									if (|{priv_lvl_i == 2'b00, priv_lvl_i == 2'b01})
										illegal_instr = 1'b1;
								end
								12'b011110110010: begin
									instruction_o[289-:7] = 7'd25;
									illegal_instr = (!debug_mode_i ? 1'b1 : 1'b0);
								end
								12'b000100000101: begin
									if (ariane_pkg_ENABLE_WFI)
										instruction_o[289-:7] = 7'd27;
									if ((priv_lvl_i == 2'b01) && tw_i) begin
										illegal_instr = 1'b1;
										instruction_o[289-:7] = 7'd0;
									end
									if (priv_lvl_i == 2'b00) begin
										illegal_instr = 1'b1;
										instruction_o[289-:7] = 7'd0;
									end
								end
								default:
									if (instr[31:25] == 7'b0001001) begin
										illegal_instr = (|{priv_lvl_i == 2'b11, priv_lvl_i == 2'b01} ? 1'b0 : 1'b1);
										instruction_o[289-:7] = 7'd30;
										if ((priv_lvl_i == 2'b01) && tvm_i)
											illegal_instr = 1'b1;
									end
							endcase
						end
						3'b001: begin
							imm_select = 4'd1;
							instruction_o[289-:7] = 7'd31;
						end
						3'b010: begin
							imm_select = 4'd1;
							if (instr[19-:5] == 5'b00000)
								instruction_o[289-:7] = 7'd32;
							else
								instruction_o[289-:7] = 7'd33;
						end
						3'b011: begin
							imm_select = 4'd1;
							if (instr[19-:5] == 5'b00000)
								instruction_o[289-:7] = 7'd32;
							else
								instruction_o[289-:7] = 7'd34;
						end
						3'b101: begin
							instruction_o[281:277] = instr[19-:5];
							imm_select = 4'd1;
							instruction_o[198] = 1'b1;
							instruction_o[289-:7] = 7'd31;
						end
						3'b110: begin
							instruction_o[281:277] = instr[19-:5];
							imm_select = 4'd1;
							instruction_o[198] = 1'b1;
							if (instr[19-:5] == 5'b00000)
								instruction_o[289-:7] = 7'd32;
							else
								instruction_o[289-:7] = 7'd33;
						end
						3'b111: begin
							instruction_o[281:277] = instr[19-:5];
							imm_select = 4'd1;
							instruction_o[198] = 1'b1;
							if (instr[19-:5] == 5'b00000)
								instruction_o[289-:7] = 7'd32;
							else
								instruction_o[289-:7] = 7'd34;
						end
						default: illegal_instr = 1'b1;
					endcase
				end
				riscv_OpcodeMiscMem: begin
					instruction_o[293-:4] = 4'd6;
					instruction_o[282-:6] = 1'sb0;
					instruction_o[276-:6] = 1'sb0;
					instruction_o[270-:6] = 1'sb0;
					case (instr[14-:3])
						3'b000: instruction_o[289-:7] = 7'd28;
						3'b001: begin
							if (instr[31:20] != {12 {1'sb0}})
								illegal_instr = 1'b1;
							instruction_o[289-:7] = 7'd29;
						end
						default: illegal_instr = 1'b1;
					endcase
					if (((instr[19-:5] != {5 {1'sb0}}) || (instr[11-:5] != {5 {1'sb0}})) || (instr[31:28] != {4 {1'sb0}}))
						illegal_instr = 1'b1;
				end
				riscv_OpcodeOp:
					if (instr[31-:2] == 2'b10) begin
						if ((ariane_pkg_FP_PRESENT && ariane_pkg_XFVEC) && (fs_i != 2'b00)) begin : sv2v_autoblock_1
							reg allow_replication;
							instruction_o[293-:4] = 4'd8;
							instruction_o[281:277] = instr[19-:5];
							instruction_o[275:271] = instr[24-:5];
							instruction_o[269:265] = instr[11-:5];
							check_fprm = 1'b1;
							allow_replication = 1'b1;
							case (instr[29-:5])
								5'b00001: begin
									instruction_o[289-:7] = 7'd89;
									instruction_o[282-:6] = 1'sb0;
									instruction_o[276-:6] = instr[19-:5];
									imm_select = 4'd1;
								end
								5'b00010: begin
									instruction_o[289-:7] = 7'd90;
									instruction_o[282-:6] = 1'sb0;
									instruction_o[276-:6] = instr[19-:5];
									imm_select = 4'd1;
								end
								5'b00011: instruction_o[289-:7] = 7'd91;
								5'b00100: instruction_o[289-:7] = 7'd92;
								5'b00101: begin
									instruction_o[289-:7] = 7'd107;
									check_fprm = 1'b0;
								end
								5'b00110: begin
									instruction_o[289-:7] = 7'd108;
									check_fprm = 1'b0;
								end
								5'b00111: begin
									instruction_o[289-:7] = 7'd94;
									allow_replication = 1'b0;
									if (instr[24-:5] != 5'b00000)
										illegal_instr = 1'b1;
								end
								5'b01000: begin
									instruction_o[289-:7] = 7'd95;
									imm_select = 4'd2;
								end
								5'b01001: begin
									instruction_o[289-:7] = 7'd96;
									imm_select = 4'd2;
								end
								5'b01100:
									if (instr[24-:5] == 5'b00000) begin
										instruction_o[276-:6] = instr[19-:5];
										if (instr[14])
											instruction_o[289-:7] = 7'd104;
										else
											instruction_o[289-:7] = 7'd103;
										check_fprm = 1'b0;
									end
									else if (instr[24-:5] == 5'b00001) begin
										instruction_o[289-:7] = 7'd106;
										check_fprm = 1'b0;
										allow_replication = 1'b0;
									end
									else if (instr[24-:5] == 5'b00010)
										instruction_o[289-:7] = 7'd99;
									else if (instr[24-:5] == 5'b00011)
										instruction_o[289-:7] = 7'd100;
									else if ((instr[24-:5] | 5'b00011) == 5'b00111) begin
										instruction_o[289-:7] = 7'd101;
										instruction_o[276-:6] = instr[11-:5];
										imm_select = 4'd1;
										case (instr[21:20])
											2'b00:
												if (~ariane_pkg_RVFVEC)
													illegal_instr = 1'b1;
											2'b01:
												if (~ariane_pkg_XF16ALTVEC)
													illegal_instr = 1'b1;
											2'b10:
												if (~ariane_pkg_XF16VEC)
													illegal_instr = 1'b1;
											2'b11:
												if (~ariane_pkg_XF8VEC)
													illegal_instr = 1'b1;
											default: illegal_instr = 1'b1;
										endcase
									end
									else
										illegal_instr = 1'b1;
								5'b01101: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd109;
								end
								5'b01110: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd110;
								end
								5'b01111: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd111;
								end
								5'b10000: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd112;
								end
								5'b10001: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd113;
								end
								5'b10010: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd114;
								end
								5'b10011: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd115;
								end
								5'b10100: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd116;
								end
								5'b10101: begin
									check_fprm = 1'b0;
									instruction_o[289-:7] = 7'd117;
								end
								5'b11000: begin
									instruction_o[289-:7] = 7'd118;
									imm_select = 4'd2;
									if (~ariane_pkg_RVF)
										illegal_instr = 1'b1;
									case (instr[13-:2])
										2'b00: begin
											if (~ariane_pkg_RVFVEC)
												illegal_instr = 1'b1;
											if (instr[14])
												illegal_instr = 1'b1;
										end
										2'b01:
											if (~ariane_pkg_XF16ALTVEC)
												illegal_instr = 1'b1;
										2'b10:
											if (~ariane_pkg_XF16VEC)
												illegal_instr = 1'b1;
										2'b11:
											if (~ariane_pkg_XF8VEC)
												illegal_instr = 1'b1;
										default: illegal_instr = 1'b1;
									endcase
								end
								5'b11001: begin
									instruction_o[289-:7] = 7'd119;
									imm_select = 4'd2;
									if (~ariane_pkg_RVF)
										illegal_instr = 1'b1;
									case (instr[13-:2])
										2'b00: illegal_instr = 1'b1;
										2'b01: illegal_instr = 1'b1;
										2'b10: illegal_instr = 1'b1;
										2'b11:
											if (~ariane_pkg_XF8VEC)
												illegal_instr = 1'b1;
										default: illegal_instr = 1'b1;
									endcase
								end
								5'b11010: begin
									instruction_o[289-:7] = 7'd120;
									imm_select = 4'd2;
									if (~ariane_pkg_RVD)
										illegal_instr = 1'b1;
									case (instr[13-:2])
										2'b00: begin
											if (~ariane_pkg_RVFVEC)
												illegal_instr = 1'b1;
											if (instr[14])
												illegal_instr = 1'b1;
										end
										2'b01:
											if (~ariane_pkg_XF16ALTVEC)
												illegal_instr = 1'b1;
										2'b10:
											if (~ariane_pkg_XF16VEC)
												illegal_instr = 1'b1;
										2'b11:
											if (~ariane_pkg_XF8VEC)
												illegal_instr = 1'b1;
										default: illegal_instr = 1'b1;
									endcase
								end
								5'b11011: begin
									instruction_o[289-:7] = 7'd121;
									imm_select = 4'd2;
									if (~ariane_pkg_RVD)
										illegal_instr = 1'b1;
									case (instr[13-:2])
										2'b00: illegal_instr = 1'b1;
										2'b01: illegal_instr = 1'b1;
										2'b10: illegal_instr = 1'b1;
										2'b11:
											if (~ariane_pkg_XF8VEC)
												illegal_instr = 1'b1;
										default: illegal_instr = 1'b1;
									endcase
								end
								default: illegal_instr = 1'b1;
							endcase
							case (instr[13-:2])
								2'b00:
									if (~ariane_pkg_RVFVEC)
										illegal_instr = 1'b1;
								2'b01:
									if (~ariane_pkg_XF16ALTVEC)
										illegal_instr = 1'b1;
								2'b10:
									if (~ariane_pkg_XF16VEC)
										illegal_instr = 1'b1;
								2'b11:
									if (~ariane_pkg_XF8VEC)
										illegal_instr = 1'b1;
								default: illegal_instr = 1'b1;
							endcase
							if (~allow_replication & instr[14])
								illegal_instr = 1'b1;
							if (check_fprm) begin
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									;
								else
									illegal_instr = 1'b1;
							end
						end
						else
							illegal_instr = 1'b1;
					end
					else begin
						instruction_o[293-:4] = (instr[31-:7] == 7'b0000001 ? 4'd5 : 4'd3);
						instruction_o[282-:6] = instr[19-:5];
						instruction_o[276-:6] = instr[24-:5];
						instruction_o[270-:6] = instr[11-:5];
						case ({instr[31-:7], instr[14-:3]})
							10'b0000000000: instruction_o[289-:7] = 7'd0;
							10'b0100000000: instruction_o[289-:7] = 7'd1;
							10'b0000000010: instruction_o[289-:7] = 7'd21;
							10'b0000000011: instruction_o[289-:7] = 7'd22;
							10'b0000000100: instruction_o[289-:7] = 7'd4;
							10'b0000000110: instruction_o[289-:7] = 7'd5;
							10'b0000000111: instruction_o[289-:7] = 7'd6;
							10'b0000000001: instruction_o[289-:7] = 7'd9;
							10'b0000000101: instruction_o[289-:7] = 7'd8;
							10'b0100000101: instruction_o[289-:7] = 7'd7;
							10'b0000001000: instruction_o[289-:7] = 7'd68;
							10'b0000001001: instruction_o[289-:7] = 7'd69;
							10'b0000001010: instruction_o[289-:7] = 7'd71;
							10'b0000001011: instruction_o[289-:7] = 7'd70;
							10'b0000001100: instruction_o[289-:7] = 7'd73;
							10'b0000001101: instruction_o[289-:7] = 7'd74;
							10'b0000001110: instruction_o[289-:7] = 7'd77;
							10'b0000001111: instruction_o[289-:7] = 7'd78;
							default: illegal_instr = 1'b1;
						endcase
					end
				riscv_OpcodeOp32: begin
					instruction_o[293-:4] = (instr[31-:7] == 7'b0000001 ? 4'd5 : 4'd3);
					instruction_o[281:277] = instr[19-:5];
					instruction_o[275:271] = instr[24-:5];
					instruction_o[269:265] = instr[11-:5];
					if (riscv_IS_XLEN64)
						case ({instr[31-:7], instr[14-:3]})
							10'b0000000000: instruction_o[289-:7] = 7'd2;
							10'b0100000000: instruction_o[289-:7] = 7'd3;
							10'b0000000001: instruction_o[289-:7] = 7'd11;
							10'b0000000101: instruction_o[289-:7] = 7'd10;
							10'b0100000101: instruction_o[289-:7] = 7'd12;
							10'b0000001000: instruction_o[289-:7] = 7'd72;
							10'b0000001100: instruction_o[289-:7] = 7'd75;
							10'b0000001101: instruction_o[289-:7] = 7'd76;
							10'b0000001110: instruction_o[289-:7] = 7'd79;
							10'b0000001111: instruction_o[289-:7] = 7'd80;
							default: illegal_instr = 1'b1;
						endcase
					else
						illegal_instr = 1'b1;
				end
				riscv_OpcodeOpImm: begin
					instruction_o[293-:4] = 4'd3;
					imm_select = 4'd1;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[269:265] = instr[11-:5];
					case (instr[14-:3])
						3'b000: instruction_o[289-:7] = 7'd0;
						3'b010: instruction_o[289-:7] = 7'd21;
						3'b011: instruction_o[289-:7] = 7'd22;
						3'b100: instruction_o[289-:7] = 7'd4;
						3'b110: instruction_o[289-:7] = 7'd5;
						3'b111: instruction_o[289-:7] = 7'd6;
						3'b001: begin
							instruction_o[289-:7] = 7'd9;
							if (instr[31:26] != 6'b000000)
								illegal_instr = 1'b1;
							if ((instr[25] != 1'b0) && 1'd0)
								illegal_instr = 1'b1;
						end
						3'b101: begin
							if (instr[31:26] == 6'b000000)
								instruction_o[289-:7] = 7'd8;
							else if (instr[31:26] == 6'b010000)
								instruction_o[289-:7] = 7'd7;
							else
								illegal_instr = 1'b1;
							if ((instr[25] != 1'b0) && 1'd0)
								illegal_instr = 1'b1;
						end
					endcase
				end
				riscv_OpcodeOpImm32: begin
					instruction_o[293-:4] = 4'd3;
					imm_select = 4'd1;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[269:265] = instr[11-:5];
					if (riscv_IS_XLEN64)
						case (instr[14-:3])
							3'b000: instruction_o[289-:7] = 7'd2;
							3'b001: begin
								instruction_o[289-:7] = 7'd11;
								if (instr[31:25] != 7'b0000000)
									illegal_instr = 1'b1;
							end
							3'b101:
								if (instr[31:25] == 7'b0000000)
									instruction_o[289-:7] = 7'd10;
								else if (instr[31:25] == 7'b0100000)
									instruction_o[289-:7] = 7'd12;
								else
									illegal_instr = 1'b1;
							default: illegal_instr = 1'b1;
						endcase
					else
						illegal_instr = 1'b1;
				end
				riscv_OpcodeStore: begin
					instruction_o[293-:4] = 4'd2;
					imm_select = 4'd2;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[275:271] = instr[24-:5];
					case (instr[14-:3])
						3'b000: instruction_o[289-:7] = 7'd44;
						3'b001: instruction_o[289-:7] = 7'd42;
						3'b010: instruction_o[289-:7] = 7'd39;
						3'b011: instruction_o[289-:7] = 7'd36;
						default: illegal_instr = 1'b1;
					endcase
				end
				riscv_OpcodeLoad: begin
					instruction_o[293-:4] = 4'd1;
					imm_select = 4'd1;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[269:265] = instr[11-:5];
					case (instr[14-:3])
						3'b000: instruction_o[289-:7] = 7'd43;
						3'b001: instruction_o[289-:7] = 7'd40;
						3'b010: instruction_o[289-:7] = 7'd37;
						3'b100: instruction_o[289-:7] = 7'd45;
						3'b101: instruction_o[289-:7] = 7'd41;
						3'b110: instruction_o[289-:7] = 7'd38;
						3'b011: instruction_o[289-:7] = 7'd35;
						default: illegal_instr = 1'b1;
					endcase
				end
				riscv_OpcodeStoreFp:
					if (ariane_pkg_FP_PRESENT && (fs_i != 2'b00)) begin
						instruction_o[293-:4] = 4'd2;
						imm_select = 4'd2;
						instruction_o[282-:6] = instr[19-:5];
						instruction_o[276-:6] = instr[24-:5];
						case (instr[14-:3])
							3'b000:
								if (ariane_pkg_XF8)
									instruction_o[289-:7] = 7'd88;
								else
									illegal_instr = 1'b1;
							3'b001:
								if (ariane_pkg_XF16 | ariane_pkg_XF16ALT)
									instruction_o[289-:7] = 7'd87;
								else
									illegal_instr = 1'b1;
							3'b010:
								if (ariane_pkg_RVF)
									instruction_o[289-:7] = 7'd86;
								else
									illegal_instr = 1'b1;
							3'b011:
								if (ariane_pkg_RVD)
									instruction_o[289-:7] = 7'd85;
								else
									illegal_instr = 1'b1;
							default: illegal_instr = 1'b1;
						endcase
					end
					else
						illegal_instr = 1'b1;
				riscv_OpcodeLoadFp:
					if (ariane_pkg_FP_PRESENT && (fs_i != 2'b00)) begin
						instruction_o[293-:4] = 4'd1;
						imm_select = 4'd1;
						instruction_o[282-:6] = instr[19-:5];
						instruction_o[270-:6] = instr[11-:5];
						case (instr[14-:3])
							3'b000:
								if (ariane_pkg_XF8)
									instruction_o[289-:7] = 7'd84;
								else
									illegal_instr = 1'b1;
							3'b001:
								if (ariane_pkg_XF16 | ariane_pkg_XF16ALT)
									instruction_o[289-:7] = 7'd83;
								else
									illegal_instr = 1'b1;
							3'b010:
								if (ariane_pkg_RVF)
									instruction_o[289-:7] = 7'd82;
								else
									illegal_instr = 1'b1;
							3'b011:
								if (ariane_pkg_RVD)
									instruction_o[289-:7] = 7'd81;
								else
									illegal_instr = 1'b1;
							default: illegal_instr = 1'b1;
						endcase
					end
					else
						illegal_instr = 1'b1;
				riscv_OpcodeMadd, riscv_OpcodeMsub, riscv_OpcodeNmsub, riscv_OpcodeNmadd:
					if (ariane_pkg_FP_PRESENT && (fs_i != 2'b00)) begin
						instruction_o[293-:4] = 4'd7;
						instruction_o[282-:6] = instr[19-:5];
						instruction_o[276-:6] = instr[24-:5];
						instruction_o[270-:6] = instr[11-:5];
						imm_select = 4'd6;
						check_fprm = 1'b1;
						case (instr[6-:7])
							default: instruction_o[289-:7] = 7'd95;
							riscv_OpcodeMsub: instruction_o[289-:7] = 7'd96;
							riscv_OpcodeNmsub: instruction_o[289-:7] = 7'd97;
							riscv_OpcodeNmadd: instruction_o[289-:7] = 7'd98;
						endcase
						case (instr[26-:2])
							2'b00:
								if (~ariane_pkg_RVF)
									illegal_instr = 1'b1;
							2'b01:
								if (~ariane_pkg_RVD)
									illegal_instr = 1'b1;
							2'b10:
								if (~ariane_pkg_XF16 & ~ariane_pkg_XF16ALT)
									illegal_instr = 1'b1;
							2'b11:
								if (~ariane_pkg_XF8)
									illegal_instr = 1'b1;
							default: illegal_instr = 1'b1;
						endcase
						if (check_fprm) begin
							if ((3'b000 <= instr[14-:3]) && (3'b100 >= instr[14-:3]))
								;
							else if (instr[14-:3] == 3'b101) begin
								if (~ariane_pkg_XF16ALT || (instr[26-:2] != 2'b10))
									illegal_instr = 1'b1;
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									;
								else
									illegal_instr = 1'b1;
							end
							else if (instr[14-:3] == 3'b111) begin
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									;
								else
									illegal_instr = 1'b1;
							end
							else
								illegal_instr = 1'b1;
						end
					end
					else
						illegal_instr = 1'b1;
				riscv_OpcodeOpFp:
					if (ariane_pkg_FP_PRESENT && (fs_i != 2'b00)) begin
						instruction_o[293-:4] = 4'd7;
						instruction_o[282-:6] = instr[19-:5];
						instruction_o[276-:6] = instr[24-:5];
						instruction_o[270-:6] = instr[11-:5];
						check_fprm = 1'b1;
						case (instr[31-:5])
							5'b00000: begin
								instruction_o[289-:7] = 7'd89;
								instruction_o[282-:6] = 1'sb0;
								instruction_o[276-:6] = instr[19-:5];
								imm_select = 4'd1;
							end
							5'b00001: begin
								instruction_o[289-:7] = 7'd90;
								instruction_o[282-:6] = 1'sb0;
								instruction_o[276-:6] = instr[19-:5];
								imm_select = 4'd1;
							end
							5'b00010: instruction_o[289-:7] = 7'd91;
							5'b00011: instruction_o[289-:7] = 7'd92;
							5'b01011: begin
								instruction_o[289-:7] = 7'd94;
								if (instr[24-:5] != 5'b00000)
									illegal_instr = 1'b1;
							end
							5'b00100: begin
								instruction_o[289-:7] = 7'd102;
								check_fprm = 1'b0;
								if (ariane_pkg_XF16ALT) begin
									if (!(|{(3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b110 >= instr[14-:3])}))
										illegal_instr = 1'b1;
								end
								else if (!((3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3])))
									illegal_instr = 1'b1;
							end
							5'b00101: begin
								instruction_o[289-:7] = 7'd93;
								check_fprm = 1'b0;
								if (ariane_pkg_XF16ALT) begin
									if (!(|{(3'b000 <= instr[14-:3]) && (3'b001 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b101 >= instr[14-:3])}))
										illegal_instr = 1'b1;
								end
								else if (!((3'b000 <= instr[14-:3]) && (3'b001 >= instr[14-:3])))
									illegal_instr = 1'b1;
							end
							5'b01000: begin
								instruction_o[289-:7] = 7'd101;
								instruction_o[276-:6] = instr[19-:5];
								imm_select = 4'd1;
								if (instr[24:23])
									illegal_instr = 1'b1;
								case (instr[22:20])
									3'b000:
										if (~ariane_pkg_RVF)
											illegal_instr = 1'b1;
									3'b001:
										if (~ariane_pkg_RVD)
											illegal_instr = 1'b1;
									3'b010:
										if (~ariane_pkg_XF16)
											illegal_instr = 1'b1;
									3'b110:
										if (~ariane_pkg_XF16ALT)
											illegal_instr = 1'b1;
									3'b011:
										if (~ariane_pkg_XF8)
											illegal_instr = 1'b1;
									default: illegal_instr = 1'b1;
								endcase
							end
							5'b10100: begin
								instruction_o[289-:7] = 7'd105;
								check_fprm = 1'b0;
								if (ariane_pkg_XF16ALT) begin
									if (!(|{(3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3]), (3'b100 <= instr[14-:3]) && (3'b110 >= instr[14-:3])}))
										illegal_instr = 1'b1;
								end
								else if (!((3'b000 <= instr[14-:3]) && (3'b010 >= instr[14-:3])))
									illegal_instr = 1'b1;
							end
							5'b11000: begin
								instruction_o[289-:7] = 7'd99;
								imm_select = 4'd1;
								if (instr[24:22])
									illegal_instr = 1'b1;
							end
							5'b11010: begin
								instruction_o[289-:7] = 7'd100;
								imm_select = 4'd1;
								if (instr[24:22])
									illegal_instr = 1'b1;
							end
							5'b11100: begin
								instruction_o[276-:6] = instr[19-:5];
								check_fprm = 1'b0;
								if ((instr[14-:3] == 3'b000) || (ariane_pkg_XF16ALT && (instr[14-:3] == 3'b100)))
									instruction_o[289-:7] = 7'd103;
								else if ((instr[14-:3] == 3'b001) || (ariane_pkg_XF16ALT && (instr[14-:3] == 3'b101)))
									instruction_o[289-:7] = 7'd106;
								else
									illegal_instr = 1'b1;
								if (instr[24-:5] != 5'b00000)
									illegal_instr = 1'b1;
							end
							5'b11110: begin
								instruction_o[289-:7] = 7'd104;
								instruction_o[276-:6] = instr[19-:5];
								check_fprm = 1'b0;
								if (!((instr[14-:3] == 3'b000) || (ariane_pkg_XF16ALT && (instr[14-:3] == 3'b100))))
									illegal_instr = 1'b1;
								if (instr[24-:5] != 5'b00000)
									illegal_instr = 1'b1;
							end
							default: illegal_instr = 1'b1;
						endcase
						case (instr[26-:2])
							2'b00:
								if (~ariane_pkg_RVF)
									illegal_instr = 1'b1;
							2'b01:
								if (~ariane_pkg_RVD)
									illegal_instr = 1'b1;
							2'b10:
								if (~ariane_pkg_XF16 & ~ariane_pkg_XF16ALT)
									illegal_instr = 1'b1;
							2'b11:
								if (~ariane_pkg_XF8)
									illegal_instr = 1'b1;
							default: illegal_instr = 1'b1;
						endcase
						if (check_fprm) begin
							if ((3'b000 <= instr[14-:3]) && (3'b100 >= instr[14-:3]))
								;
							else if (instr[14-:3] == 3'b101) begin
								if (~ariane_pkg_XF16ALT || (instr[26-:2] != 2'b10))
									illegal_instr = 1'b1;
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									;
								else
									illegal_instr = 1'b1;
							end
							else if (instr[14-:3] == 3'b111) begin
								if ((3'b000 <= frm_i) && (3'b100 >= frm_i))
									;
								else
									illegal_instr = 1'b1;
							end
							else
								illegal_instr = 1'b1;
						end
					end
					else
						illegal_instr = 1'b1;
				riscv_OpcodeAmo: begin
					instruction_o[293-:4] = 4'd2;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[275:271] = instr[24-:5];
					instruction_o[269:265] = instr[11-:5];
					if (ariane_pkg_RVA && (instr[14-:3] == 3'h2))
						case (instr[31:27])
							5'h00: instruction_o[289-:7] = 7'd51;
							5'h01: instruction_o[289-:7] = 7'd50;
							5'h02: begin
								instruction_o[289-:7] = 7'd46;
								if (instr[24-:5] != 0)
									illegal_instr = 1'b1;
							end
							5'h03: instruction_o[289-:7] = 7'd48;
							5'h04: instruction_o[289-:7] = 7'd54;
							5'h08: instruction_o[289-:7] = 7'd53;
							5'h0c: instruction_o[289-:7] = 7'd52;
							5'h10: instruction_o[289-:7] = 7'd57;
							5'h14: instruction_o[289-:7] = 7'd55;
							5'h18: instruction_o[289-:7] = 7'd58;
							5'h1c: instruction_o[289-:7] = 7'd56;
							default: illegal_instr = 1'b1;
						endcase
					else if (ariane_pkg_RVA && (instr[14-:3] == 3'h3))
						case (instr[31:27])
							5'h00: instruction_o[289-:7] = 7'd60;
							5'h01: instruction_o[289-:7] = 7'd59;
							5'h02: begin
								instruction_o[289-:7] = 7'd47;
								if (instr[24-:5] != 0)
									illegal_instr = 1'b1;
							end
							5'h03: instruction_o[289-:7] = 7'd49;
							5'h04: instruction_o[289-:7] = 7'd63;
							5'h08: instruction_o[289-:7] = 7'd62;
							5'h0c: instruction_o[289-:7] = 7'd61;
							5'h10: instruction_o[289-:7] = 7'd66;
							5'h14: instruction_o[289-:7] = 7'd64;
							5'h18: instruction_o[289-:7] = 7'd67;
							5'h1c: instruction_o[289-:7] = 7'd65;
							default: illegal_instr = 1'b1;
						endcase
					else
						illegal_instr = 1'b1;
				end
				riscv_OpcodeBranch: begin
					imm_select = 4'd3;
					instruction_o[293-:4] = 4'd4;
					instruction_o[281:277] = instr[19-:5];
					instruction_o[275:271] = instr[24-:5];
					is_control_flow_instr_o = 1'b1;
					case (instr[14-:3])
						3'b000: instruction_o[289-:7] = 7'd17;
						3'b001: instruction_o[289-:7] = 7'd18;
						3'b100: instruction_o[289-:7] = 7'd13;
						3'b101: instruction_o[289-:7] = 7'd15;
						3'b110: instruction_o[289-:7] = 7'd14;
						3'b111: instruction_o[289-:7] = 7'd16;
						default: begin
							is_control_flow_instr_o = 1'b0;
							illegal_instr = 1'b1;
						end
					endcase
				end
				riscv_OpcodeJalr: begin
					instruction_o[293-:4] = 4'd4;
					instruction_o[289-:7] = 7'd19;
					instruction_o[281:277] = instr[19-:5];
					imm_select = 4'd1;
					instruction_o[269:265] = instr[11-:5];
					is_control_flow_instr_o = 1'b1;
					if (instr[14-:3] != 3'b000)
						illegal_instr = 1'b1;
				end
				riscv_OpcodeJal: begin
					instruction_o[293-:4] = 4'd4;
					imm_select = 4'd5;
					instruction_o[269:265] = instr[11-:5];
					is_control_flow_instr_o = 1'b1;
				end
				riscv_OpcodeAuipc: begin
					instruction_o[293-:4] = 4'd3;
					imm_select = 4'd4;
					instruction_o[197] = 1'b1;
					instruction_o[269:265] = instr[11-:5];
				end
				riscv_OpcodeLui: begin
					imm_select = 4'd4;
					instruction_o[293-:4] = 4'd3;
					instruction_o[269:265] = instr[11-:5];
				end
				default: illegal_instr = 1'b1;
			endcase
	end
	always @(*) begin : sign_extend
		imm_i_type = {{52 {instruction_i[31]}}, instruction_i[31:20]};
		imm_s_type = {{52 {instruction_i[31]}}, instruction_i[31:25], instruction_i[11:7]};
		imm_sb_type = {{51 {instruction_i[31]}}, instruction_i[31], instruction_i[7], instruction_i[30:25], instruction_i[11:8], 1'b0};
		imm_u_type = {{32 {instruction_i[31]}}, instruction_i[31:12], 12'b000000000000};
		imm_uj_type = {{44 {instruction_i[31]}}, instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0};
		imm_bi_type = {{59 {instruction_i[24]}}, instruction_i[24:20]};
		case (imm_select)
			4'd1: begin
				instruction_o[264-:64] = imm_i_type;
				instruction_o[199] = 1'b1;
			end
			4'd2: begin
				instruction_o[264-:64] = imm_s_type;
				instruction_o[199] = 1'b1;
			end
			4'd3: begin
				instruction_o[264-:64] = imm_sb_type;
				instruction_o[199] = 1'b1;
			end
			4'd4: begin
				instruction_o[264-:64] = imm_u_type;
				instruction_o[199] = 1'b1;
			end
			4'd5: begin
				instruction_o[264-:64] = imm_uj_type;
				instruction_o[199] = 1'b1;
			end
			4'd6: begin
				instruction_o[264-:64] = {{59 {1'b0}}, instr[31-:5]};
				instruction_o[199] = 1'b0;
			end
			default: begin
				instruction_o[264-:64] = {riscv_XLEN {1'b0}};
				instruction_o[199] = 1'b0;
			end
		endcase
	end
	reg [63:0] interrupt_cause;
	wire [1:1] sv2v_tmp_DF233;
	assign sv2v_tmp_DF233 = instruction_o[68];
	always @(*) instruction_o[200] = sv2v_tmp_DF233;
	localparam ariane_pkg_SupervisorIrq = 1;
	localparam [63:0] riscv_BREAKPOINT = 3;
	localparam [63:0] riscv_DEBUG_REQUEST = 24;
	localparam [63:0] riscv_ENV_CALL_MMODE = 11;
	localparam [63:0] riscv_ENV_CALL_SMODE = 9;
	localparam [63:0] riscv_ENV_CALL_UMODE = 8;
	localparam [63:0] riscv_ILLEGAL_INSTR = 2;
	localparam [31:0] riscv_IRQ_M_EXT = 11;
	localparam [63:0] riscv_M_EXT_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_M_EXT;
	localparam [31:0] riscv_IRQ_M_SOFT = 3;
	localparam [63:0] riscv_M_SW_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_M_SOFT;
	localparam [31:0] riscv_IRQ_M_TIMER = 7;
	localparam [63:0] riscv_M_TIMER_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_M_TIMER;
	localparam [31:0] riscv_IRQ_S_EXT = 9;
	localparam [63:0] riscv_S_EXT_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_S_EXT;
	localparam [31:0] riscv_IRQ_S_SOFT = 1;
	localparam [63:0] riscv_S_SW_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_S_SOFT;
	localparam [31:0] riscv_IRQ_S_TIMER = 5;
	localparam [63:0] riscv_S_TIMER_INTERRUPT = 65'sd9223372036854775808 | riscv_IRQ_S_TIMER;
	always @(*) begin : exception_handling
		interrupt_cause = 1'sb0;
		instruction_o[196-:129] = ex_i;
		if (~ex_i[0]) begin
			instruction_o[132-:64] = (is_compressed_i ? {{48 {1'b0}}, compressed_instr_i} : {{32 {1'b0}}, instruction_i});
			if (illegal_instr || is_illegal_i) begin
				instruction_o[68] = 1'b1;
				instruction_o[196-:64] = riscv_ILLEGAL_INSTR;
			end
			else if (ecall) begin
				instruction_o[68] = 1'b1;
				case (priv_lvl_i)
					2'b11: instruction_o[196-:64] = riscv_ENV_CALL_MMODE;
					2'b01: instruction_o[196-:64] = riscv_ENV_CALL_SMODE;
					2'b00: instruction_o[196-:64] = riscv_ENV_CALL_UMODE;
					default:
						;
				endcase
			end
			else if (ebreak) begin
				instruction_o[68] = 1'b1;
				instruction_o[196-:64] = riscv_BREAKPOINT;
			end
			if (irq_ctrl_i[130 + riscv_S_TIMER_INTERRUPT[5:0]] && irq_ctrl_i[66 + riscv_S_TIMER_INTERRUPT[5:0]])
				interrupt_cause = riscv_S_TIMER_INTERRUPT;
			if (irq_ctrl_i[130 + riscv_S_SW_INTERRUPT[5:0]] && irq_ctrl_i[66 + riscv_S_SW_INTERRUPT[5:0]])
				interrupt_cause = riscv_S_SW_INTERRUPT;
			if (irq_ctrl_i[130 + riscv_S_EXT_INTERRUPT[5:0]] && (irq_ctrl_i[66 + riscv_S_EXT_INTERRUPT[5:0]] | irq_i[ariane_pkg_SupervisorIrq]))
				interrupt_cause = riscv_S_EXT_INTERRUPT;
			if (irq_ctrl_i[66 + riscv_M_TIMER_INTERRUPT[5:0]] && irq_ctrl_i[130 + riscv_M_TIMER_INTERRUPT[5:0]])
				interrupt_cause = riscv_M_TIMER_INTERRUPT;
			if (irq_ctrl_i[66 + riscv_M_SW_INTERRUPT[5:0]] && irq_ctrl_i[130 + riscv_M_SW_INTERRUPT[5:0]])
				interrupt_cause = riscv_M_SW_INTERRUPT;
			if (irq_ctrl_i[66 + riscv_M_EXT_INTERRUPT[5:0]] && irq_ctrl_i[130 + riscv_M_EXT_INTERRUPT[5:0]])
				interrupt_cause = riscv_M_EXT_INTERRUPT;
			if (interrupt_cause[63] && irq_ctrl_i[0]) begin
				if (irq_ctrl_i[2 + interrupt_cause[5:0]]) begin
					if ((irq_ctrl_i[1] && (priv_lvl_i == 2'b01)) || (priv_lvl_i == 2'b00)) begin
						instruction_o[68] = 1'b1;
						instruction_o[196-:64] = interrupt_cause;
					end
				end
				else begin
					instruction_o[68] = 1'b1;
					instruction_o[196-:64] = interrupt_cause;
				end
			end
		end
		if (debug_req_i && !debug_mode_i) begin
			instruction_o[68] = 1'b1;
			instruction_o[196-:64] = riscv_DEBUG_REQUEST;
		end
	end
endmodule
module dromajo_ram (
	Clk_CI,
	Rst_RBI,
	CSel_SI,
	WrEn_SI,
	BEn_SI,
	WrData_DI,
	Addr_DI,
	RdData_DO
);
	parameter ADDR_WIDTH = 10;
	parameter DATA_DEPTH = 1024;
	parameter OUT_REGS = 0;
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire CSel_SI;
	input wire WrEn_SI;
	input wire [7:0] BEn_SI;
	input wire [63:0] WrData_DI;
	input wire [ADDR_WIDTH - 1:0] Addr_DI;
	output wire [63:0] RdData_DO;
	localparam DATA_BYTES = 8;
	reg [63:0] RdData_DN;
	reg [63:0] RdData_DP;
	reg [63:0] Mem_DP [DATA_DEPTH - 1:0];
	// initial begin : sv2v_autoblock_1
	// 	integer hex_file;
	// 	integer num_bytes;
	// 	reg signed [63:0] address;
	// 	reg signed [63:0] value;
	// 	string f_name;
	// 	begin : sv2v_autoblock_2
	// 		reg signed [31:0] k;
	// 		for (k = 0; k < DATA_DEPTH; k = k + 1)
	// 			Mem_DP[k] = 0;
	// 	end
	// 	if ($value$plusargs("checkpoint=%s", f_name)) begin
	// 		hex_file = $fopen({f_name, ".mainram.hex"}, "r");
	// 		while (!$feof(hex_file)) begin
	// 			num_bytes = $fscanf(hex_file, "%d %h\n", address, value);
	// 			Mem_DP[address] = value;
	// 		end
	// 		$display("Done syncing RAM with dromajo...\n");
	// 	end
	// 	else
	// 		$display("Failed syncing RAM: provide path to a checkpoint.\n");
	// end
	always @(posedge Clk_CI)
		if (CSel_SI) begin
			if (WrEn_SI) begin
				if (BEn_SI[0])
					Mem_DP[Addr_DI][7:0] <= WrData_DI[7:0];
				if (BEn_SI[1])
					Mem_DP[Addr_DI][15:8] <= WrData_DI[15:8];
				if (BEn_SI[2])
					Mem_DP[Addr_DI][23:16] <= WrData_DI[23:16];
				if (BEn_SI[3])
					Mem_DP[Addr_DI][31:24] <= WrData_DI[31:24];
				if (BEn_SI[4])
					Mem_DP[Addr_DI][39:32] <= WrData_DI[39:32];
				if (BEn_SI[5])
					Mem_DP[Addr_DI][47:40] <= WrData_DI[47:40];
				if (BEn_SI[6])
					Mem_DP[Addr_DI][55:48] <= WrData_DI[55:48];
				if (BEn_SI[7])
					Mem_DP[Addr_DI][63:56] <= WrData_DI[63:56];
			end
			RdData_DN <= Mem_DP[Addr_DI];
		end
	generate
		if (OUT_REGS > 0) begin : g_outreg
			always @(posedge Clk_CI or negedge Rst_RBI)
				if (Rst_RBI == 1'b0)
					RdData_DP <= 0;
				else
					RdData_DP <= RdData_DN;
		end
		if (OUT_REGS == 0) begin : g_oureg_byp
			wire [64:1] sv2v_tmp_7FD8C;
			assign sv2v_tmp_7FD8C = RdData_DN;
			always @(*) RdData_DP = sv2v_tmp_7FD8C;
		end
	endgenerate
	assign RdData_DO = RdData_DP;
endmodule
module ex_stage (
	clk_i,
	rst_ni,
	flush_i,
	debug_mode_i,
	rs1_forwarding_i,
	rs2_forwarding_i,
	fu_data_i,
	pc_i,
	is_compressed_instr_i,
	flu_result_o,
	flu_trans_id_o,
	flu_exception_o,
	flu_ready_o,
	flu_valid_o,
	alu_valid_i,
	branch_valid_i,
	branch_predict_i,
	resolved_branch_o,
	resolve_branch_o,
	csr_valid_i,
	csr_addr_o,
	csr_commit_i,
	mult_valid_i,
	lsu_ready_o,
	lsu_valid_i,
	load_valid_o,
	load_result_o,
	load_trans_id_o,
	load_exception_o,
	store_valid_o,
	store_result_o,
	store_trans_id_o,
	store_exception_o,
	lsu_commit_i,
	lsu_commit_ready_o,
	commit_tran_id_i,
	no_st_pending_o,
	amo_valid_commit_i,
	fpu_ready_o,
	fpu_valid_i,
	fpu_fmt_i,
	fpu_rm_i,
	fpu_frm_i,
	fpu_prec_i,
	fpu_trans_id_o,
	fpu_result_o,
	fpu_valid_o,
	fpu_exception_o,
	enable_translation_i,
	en_ld_st_translation_i,
	flush_tlb_i,
	priv_lvl_i,
	ld_st_priv_lvl_i,
	sum_i,
	mxr_i,
	satp_ppn_i,
	asid_i,
	icache_areq_i,
	icache_areq_o,
	dcache_req_ports_i,
	dcache_req_ports_o,
	dcache_wbuffer_empty_i,
	dcache_wbuffer_not_ni_i,
	amo_req_o,
	amo_resp_i,
	itlb_miss_o,
	dtlb_miss_o,
	pmpcfg_i,
	pmpaddr_i
);
	parameter [31:0] ASID_WIDTH = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire debug_mode_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] rs1_forwarding_i;
	input wire [63:0] rs2_forwarding_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	input wire [205:0] fu_data_i;
	input wire [63:0] pc_i;
	input wire is_compressed_instr_i;
	output reg [63:0] flu_result_o;
	output reg [2:0] flu_trans_id_o;
	output wire [128:0] flu_exception_o;
	output reg flu_ready_o;
	output wire flu_valid_o;
	input wire alu_valid_i;
	input wire branch_valid_i;
	input wire [66:0] branch_predict_i;
	output wire [133:0] resolved_branch_o;
	output wire resolve_branch_o;
	input wire csr_valid_i;
	output wire [11:0] csr_addr_o;
	input wire csr_commit_i;
	input wire mult_valid_i;
	output wire lsu_ready_o;
	input wire lsu_valid_i;
	output wire load_valid_o;
	output wire [63:0] load_result_o;
	output wire [2:0] load_trans_id_o;
	output wire [128:0] load_exception_o;
	output wire store_valid_o;
	output wire [63:0] store_result_o;
	output wire [2:0] store_trans_id_o;
	output wire [128:0] store_exception_o;
	input wire lsu_commit_i;
	output wire lsu_commit_ready_o;
	input wire [2:0] commit_tran_id_i;
	output wire no_st_pending_o;
	input wire amo_valid_commit_i;
	output wire fpu_ready_o;
	input wire fpu_valid_i;
	input wire [1:0] fpu_fmt_i;
	input wire [2:0] fpu_rm_i;
	input wire [2:0] fpu_frm_i;
	input wire [6:0] fpu_prec_i;
	output wire [2:0] fpu_trans_id_o;
	output wire [63:0] fpu_result_o;
	output wire fpu_valid_o;
	output wire [128:0] fpu_exception_o;
	input wire enable_translation_i;
	input wire en_ld_st_translation_i;
	input wire flush_tlb_i;
	input wire [1:0] priv_lvl_i;
	input wire [1:0] ld_st_priv_lvl_i;
	input wire sum_i;
	input wire mxr_i;
	localparam riscv_PPNW = 44;
	input wire [43:0] satp_ppn_i;
	input wire [ASID_WIDTH - 1:0] asid_i;
	input wire [64:0] icache_areq_i;
	localparam riscv_PLEN = 56;
	output wire [185:0] icache_areq_o;
	input wire [197:0] dcache_req_ports_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (3 * ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78)) - 1 : (3 * (1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 76)):(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)] dcache_req_ports_o;
	input wire dcache_wbuffer_empty_i;
	input wire dcache_wbuffer_not_ni_i;
	output wire [134:0] amo_req_o;
	input wire [64:0] amo_resp_i;
	output wire itlb_miss_o;
	output wire dtlb_miss_o;
	input wire [127:0] pmpcfg_i;
	input wire [863:0] pmpaddr_i;
	reg current_instruction_is_sfence_vma;
	reg [ASID_WIDTH - 1:0] asid_to_be_flushed;
	reg [63:0] vaddr_to_be_flushed;
	wire alu_branch_res;
	wire [63:0] alu_result;
	wire [63:0] csr_result;
	wire [63:0] mult_result;
	wire [63:0] branch_result;
	wire csr_ready;
	wire mult_ready;
	wire [2:0] mult_trans_id;
	wire mult_valid;
	wire [205:0] alu_data;
	assign alu_data = (alu_valid_i | branch_valid_i ? fu_data_i : {206 {1'sb0}});
	alu alu_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.fu_data_i(alu_data),
		.result_o(alu_result),
		.alu_branch_res_o(alu_branch_res)
	);
	branch_unit branch_unit_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.debug_mode_i(debug_mode_i),
		.fu_data_i(fu_data_i),
		.pc_i(pc_i),
		.is_compressed_instr_i(is_compressed_instr_i),
		.fu_valid_i((((alu_valid_i || lsu_valid_i) || csr_valid_i) || mult_valid_i) || fpu_valid_i),
		.branch_valid_i(branch_valid_i),
		.branch_comp_res_i(alu_branch_res),
		.branch_result_o(branch_result),
		.branch_predict_i(branch_predict_i),
		.resolved_branch_o(resolved_branch_o),
		.resolve_branch_o(resolve_branch_o),
		.branch_exception_o(flu_exception_o)
	);
	csr_buffer csr_buffer_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.fu_data_i(fu_data_i),
		.csr_valid_i(csr_valid_i),
		.csr_ready_o(csr_ready),
		.csr_result_o(csr_result),
		.csr_commit_i(csr_commit_i),
		.csr_addr_o(csr_addr_o)
	);
	assign flu_valid_o = ((alu_valid_i | branch_valid_i) | csr_valid_i) | mult_valid;
	always @(*) begin
		flu_result_o = {branch_result};
		flu_trans_id_o = fu_data_i[2-:ariane_pkg_TRANS_ID_BITS];
		if (alu_valid_i)
			flu_result_o = alu_result;
		else if (csr_valid_i)
			flu_result_o = csr_result;
		else if (mult_valid) begin
			flu_result_o = mult_result;
			flu_trans_id_o = mult_trans_id;
		end
	end
	always @(*) flu_ready_o = csr_ready & mult_ready;
	wire [205:0] mult_data;
	assign mult_data = (mult_valid_i ? fu_data_i : {206 {1'sb0}});
	mult i_mult(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.mult_valid_i(mult_valid_i),
		.fu_data_i(mult_data),
		.result_o(mult_result),
		.mult_valid_o(mult_valid),
		.mult_ready_o(mult_ready),
		.mult_trans_id_o(mult_trans_id)
	);
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	generate
		if (ariane_pkg_FP_PRESENT) begin : fpu_gen
			wire [205:0] fpu_data;
			assign fpu_data = (fpu_valid_i ? fu_data_i : {206 {1'sb0}});
			fpu_wrap fpu_i(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.fpu_valid_i(fpu_valid_i),
				.fpu_ready_o(fpu_ready_o),
				.fu_data_i(fpu_data),
				.fpu_fmt_i(fpu_fmt_i),
				.fpu_rm_i(fpu_rm_i),
				.fpu_frm_i(fpu_frm_i),
				.fpu_prec_i(fpu_prec_i),
				.fpu_trans_id_o(fpu_trans_id_o),
				.result_o(fpu_result_o),
				.fpu_valid_o(fpu_valid_o),
				.fpu_exception_o(fpu_exception_o)
			);
		end
		else begin : no_fpu_gen
			assign fpu_ready_o = 1'sb0;
			assign fpu_trans_id_o = 1'sb0;
			assign fpu_result_o = 1'sb0;
			assign fpu_valid_o = 1'sb0;
			assign fpu_exception_o = 1'sb0;
		end
	endgenerate
	wire [205:0] lsu_data;
	assign lsu_data = (lsu_valid_i ? fu_data_i : {206 {1'sb0}});
	load_store_unit #(
		.ASID_WIDTH(ASID_WIDTH),
		.ArianeCfg(ArianeCfg)
	) lsu_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.no_st_pending_o(no_st_pending_o),
		.fu_data_i(lsu_data),
		.lsu_ready_o(lsu_ready_o),
		.lsu_valid_i(lsu_valid_i),
		.load_trans_id_o(load_trans_id_o),
		.load_result_o(load_result_o),
		.load_valid_o(load_valid_o),
		.load_exception_o(load_exception_o),
		.store_trans_id_o(store_trans_id_o),
		.store_result_o(store_result_o),
		.store_valid_o(store_valid_o),
		.store_exception_o(store_exception_o),
		.commit_i(lsu_commit_i),
		.commit_ready_o(lsu_commit_ready_o),
		.commit_tran_id_i(commit_tran_id_i),
		.enable_translation_i(enable_translation_i),
		.en_ld_st_translation_i(en_ld_st_translation_i),
		.icache_areq_i(icache_areq_i),
		.icache_areq_o(icache_areq_o),
		.priv_lvl_i(priv_lvl_i),
		.ld_st_priv_lvl_i(ld_st_priv_lvl_i),
		.sum_i(sum_i),
		.mxr_i(mxr_i),
		.satp_ppn_i(satp_ppn_i),
		.asid_i(asid_i),
		.asid_to_be_flushed_i(asid_to_be_flushed),
		.vaddr_to_be_flushed_i(vaddr_to_be_flushed),
		.flush_tlb_i(flush_tlb_i),
		.itlb_miss_o(itlb_miss_o),
		.dtlb_miss_o(dtlb_miss_o),
		.dcache_req_ports_i(dcache_req_ports_i),
		.dcache_req_ports_o(dcache_req_ports_o),
		.dcache_wbuffer_empty_i(dcache_wbuffer_empty_i),
		.dcache_wbuffer_not_ni_i(dcache_wbuffer_not_ni_i),
		.amo_valid_commit_i(amo_valid_commit_i),
		.amo_req_o(amo_req_o),
		.amo_resp_i(amo_resp_i),
		.pmpcfg_i(pmpcfg_i),
		.pmpaddr_i(pmpaddr_i)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			current_instruction_is_sfence_vma <= 1'b0;
		else if (flush_i)
			current_instruction_is_sfence_vma <= 1'b0;
		else if ((fu_data_i[201-:7] == 7'd30) && csr_valid_i)
			current_instruction_is_sfence_vma <= 1'b1;
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			asid_to_be_flushed <= 1'sb0;
			vaddr_to_be_flushed <= 1'sb0;
		end
		else if (~current_instruction_is_sfence_vma && ~((fu_data_i[201-:7] == 7'd30) && csr_valid_i)) begin
			vaddr_to_be_flushed <= rs1_forwarding_i;
			asid_to_be_flushed <= rs2_forwarding_i[ASID_WIDTH - 1:0];
		end
endmodule
module fpu_wrap (
	clk_i,
	rst_ni,
	flush_i,
	fpu_valid_i,
	fpu_ready_o,
	fu_data_i,
	fpu_fmt_i,
	fpu_rm_i,
	fpu_frm_i,
	fpu_prec_i,
	fpu_trans_id_o,
	result_o,
	fpu_valid_o,
	fpu_exception_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire fpu_valid_i;
	output reg fpu_ready_o;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	input wire [1:0] fpu_fmt_i;
	input wire [2:0] fpu_rm_i;
	input wire [2:0] fpu_frm_i;
	input wire [6:0] fpu_prec_i;
	output wire [2:0] fpu_trans_id_o;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam ariane_pkg_FLEN = (ariane_pkg_RVD ? 64 : (ariane_pkg_RVF ? 32 : (ariane_pkg_XF16 ? 16 : (ariane_pkg_XF16ALT ? 16 : (ariane_pkg_XF8 ? 8 : 1)))));
	output wire [ariane_pkg_FLEN - 1:0] result_o;
	output wire fpu_valid_o;
	output wire [128:0] fpu_exception_o;
	reg state_q;
	reg state_d;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	localparam [31:0] ariane_pkg_LAT_COMP_FP16 = 'd1;
	localparam [31:0] ariane_pkg_LAT_COMP_FP16ALT = 'd1;
	localparam [31:0] ariane_pkg_LAT_COMP_FP32 = 'd2;
	localparam [31:0] ariane_pkg_LAT_COMP_FP64 = 'd3;
	localparam [31:0] ariane_pkg_LAT_COMP_FP8 = 'd1;
	localparam [31:0] ariane_pkg_LAT_CONV = 'd2;
	localparam [31:0] ariane_pkg_LAT_DIVSQRT = 'd2;
	localparam [31:0] ariane_pkg_LAT_NONCOMP = 'd1;
	localparam [0:0] ariane_pkg_XFVEC = 1'b0;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_5;
		input reg [4:0] inp;
		sv2v_cast_5 = inp;
	endfunction
	function automatic [3:0] sv2v_cast_4;
		input reg [3:0] inp;
		sv2v_cast_4 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	generate
		if (ariane_pkg_FP_PRESENT) begin : fpu_gen
			wire [ariane_pkg_FLEN - 1:0] operand_a_i;
			wire [ariane_pkg_FLEN - 1:0] operand_b_i;
			wire [ariane_pkg_FLEN - 1:0] operand_c_i;
			assign operand_a_i = fu_data_i[130 + ariane_pkg_FLEN:131];
			assign operand_b_i = fu_data_i[66 + ariane_pkg_FLEN:67];
			assign operand_c_i = fu_data_i[2 + ariane_pkg_FLEN:3];
			localparam OPBITS = fpnew_pkg_OP_BITS;
			localparam FMTBITS = 3;
			localparam IFMTBITS = 2;
			localparam [42:0] FPU_FEATURES = {32'd64, ariane_pkg_XFVEC, 1'b1, sv2v_cast_5({ariane_pkg_RVF, ariane_pkg_RVD, ariane_pkg_XF16, ariane_pkg_XF8, ariane_pkg_XF16ALT}), sv2v_cast_4({ariane_pkg_XFVEC && ariane_pkg_XF8, ariane_pkg_XFVEC && (ariane_pkg_XF16 || ariane_pkg_XF16ALT), 2'b11})};
			localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] FPU_IMPLEMENTATION = {sv2v_cast_CDC93({ariane_pkg_LAT_COMP_FP32, ariane_pkg_LAT_COMP_FP64, ariane_pkg_LAT_COMP_FP16, ariane_pkg_LAT_COMP_FP8, ariane_pkg_LAT_COMP_FP16ALT, {fpnew_pkg_NUM_FP_FORMATS {ariane_pkg_LAT_DIVSQRT}}, {fpnew_pkg_NUM_FP_FORMATS {ariane_pkg_LAT_NONCOMP}}, {fpnew_pkg_NUM_FP_FORMATS {ariane_pkg_LAT_CONV}}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd3};
			reg [ariane_pkg_FLEN - 1:0] operand_a_d;
			reg [ariane_pkg_FLEN - 1:0] operand_a_q;
			wire [ariane_pkg_FLEN - 1:0] operand_a;
			reg [ariane_pkg_FLEN - 1:0] operand_b_d;
			reg [ariane_pkg_FLEN - 1:0] operand_b_q;
			wire [ariane_pkg_FLEN - 1:0] operand_b;
			reg [ariane_pkg_FLEN - 1:0] operand_c_d;
			reg [ariane_pkg_FLEN - 1:0] operand_c_q;
			wire [ariane_pkg_FLEN - 1:0] operand_c;
			reg [3:0] fpu_op_d;
			reg [3:0] fpu_op_q;
			wire [3:0] fpu_op;
			reg fpu_op_mod_d;
			reg fpu_op_mod_q;
			wire fpu_op_mod;
			reg [2:0] fpu_srcfmt_d;
			reg [2:0] fpu_srcfmt_q;
			wire [2:0] fpu_srcfmt;
			reg [2:0] fpu_dstfmt_d;
			reg [2:0] fpu_dstfmt_q;
			wire [2:0] fpu_dstfmt;
			reg [1:0] fpu_ifmt_d;
			reg [1:0] fpu_ifmt_q;
			wire [1:0] fpu_ifmt;
			reg [2:0] fpu_rm_d;
			reg [2:0] fpu_rm_q;
			wire [2:0] fpu_rm;
			reg fpu_vec_op_d;
			reg fpu_vec_op_q;
			wire fpu_vec_op;
			reg [2:0] fpu_tag_d;
			reg [2:0] fpu_tag_q;
			wire [2:0] fpu_tag;
			wire fpu_in_ready;
			reg fpu_in_valid;
			wire fpu_out_ready;
			wire fpu_out_valid;
			wire [4:0] fpu_status;
			reg hold_inputs;
			reg use_hold;
			always @(*) begin : input_translation
				reg vec_replication;
				reg replicate_c;
				reg check_ah;
				operand_a_d = operand_a_i;
				operand_b_d = operand_b_i;
				operand_c_d = operand_c_i;
				fpu_op_d = sv2v_cast_A53F3(6);
				fpu_op_mod_d = 1'b0;
				fpu_dstfmt_d = sv2v_cast_0BC43('d0);
				fpu_ifmt_d = sv2v_cast_87CC5(2);
				fpu_rm_d = fpu_rm_i;
				fpu_vec_op_d = fu_data_i[205-:4] == 4'd8;
				fpu_tag_d = fu_data_i[2-:ariane_pkg_TRANS_ID_BITS];
				vec_replication = fpu_rm_i[0];
				replicate_c = 1'b0;
				check_ah = 1'b0;
				if (!((3'b000 <= fpu_rm_i) && (3'b100 >= fpu_rm_i)))
					fpu_rm_d = fpu_frm_i;
				if (fpu_vec_op_d)
					fpu_rm_d = fpu_frm_i;
				case (fpu_fmt_i)
					2'b00: fpu_dstfmt_d = sv2v_cast_0BC43('d0);
					2'b01: fpu_dstfmt_d = (fpu_vec_op_d ? sv2v_cast_0BC43('d4) : sv2v_cast_0BC43('d1));
					2'b10:
						if (!fpu_vec_op_d && (fpu_rm_i == 3'b101))
							fpu_dstfmt_d = sv2v_cast_0BC43('d4);
						else
							fpu_dstfmt_d = sv2v_cast_0BC43('d2);
					default: fpu_dstfmt_d = sv2v_cast_0BC43('d3);
				endcase
				fpu_srcfmt_d = fpu_dstfmt_d;
				case (fu_data_i[201-:7])
					7'd89: begin
						fpu_op_d = sv2v_cast_A53F3(2);
						replicate_c = 1'b1;
					end
					7'd90: begin
						fpu_op_d = sv2v_cast_A53F3(2);
						fpu_op_mod_d = 1'b1;
						replicate_c = 1'b1;
					end
					7'd91: fpu_op_d = sv2v_cast_A53F3(3);
					7'd92: fpu_op_d = sv2v_cast_A53F3(4);
					7'd93: begin
						fpu_op_d = sv2v_cast_A53F3(7);
						fpu_rm_d = {1'b0, fpu_rm_i[1:0]};
						check_ah = 1'b1;
					end
					7'd94: fpu_op_d = sv2v_cast_A53F3(5);
					7'd95: fpu_op_d = sv2v_cast_A53F3(0);
					7'd96: begin
						fpu_op_d = sv2v_cast_A53F3(0);
						fpu_op_mod_d = 1'b1;
					end
					7'd97: fpu_op_d = sv2v_cast_A53F3(1);
					7'd98: begin
						fpu_op_d = sv2v_cast_A53F3(1);
						fpu_op_mod_d = 1'b1;
					end
					7'd99: begin
						fpu_op_d = sv2v_cast_A53F3(11);
						if (fpu_vec_op_d) begin
							fpu_op_mod_d = fpu_rm_i[0];
							vec_replication = 1'b0;
							case (fpu_fmt_i)
								2'b00: fpu_ifmt_d = sv2v_cast_87CC5(2);
								2'b01, 2'b10: fpu_ifmt_d = sv2v_cast_87CC5(1);
								2'b11: fpu_ifmt_d = sv2v_cast_87CC5(0);
							endcase
						end
						else begin
							fpu_op_mod_d = operand_c_i[0];
							if (operand_c_i[1])
								fpu_ifmt_d = sv2v_cast_87CC5(3);
							else
								fpu_ifmt_d = sv2v_cast_87CC5(2);
						end
					end
					7'd100: begin
						fpu_op_d = sv2v_cast_A53F3(12);
						if (fpu_vec_op_d) begin
							fpu_op_mod_d = fpu_rm_i[0];
							vec_replication = 1'b0;
							case (fpu_fmt_i)
								2'b00: fpu_ifmt_d = sv2v_cast_87CC5(2);
								2'b01, 2'b10: fpu_ifmt_d = sv2v_cast_87CC5(1);
								2'b11: fpu_ifmt_d = sv2v_cast_87CC5(0);
							endcase
						end
						else begin
							fpu_op_mod_d = operand_c_i[0];
							if (operand_c_i[1])
								fpu_ifmt_d = sv2v_cast_87CC5(3);
							else
								fpu_ifmt_d = sv2v_cast_87CC5(2);
						end
					end
					7'd101: begin
						fpu_op_d = sv2v_cast_A53F3(10);
						if (fpu_vec_op_d) begin
							vec_replication = 1'b0;
							case (operand_c_i[1:0])
								2'b00: fpu_srcfmt_d = sv2v_cast_0BC43('d0);
								2'b01: fpu_srcfmt_d = sv2v_cast_0BC43('d4);
								2'b10: fpu_srcfmt_d = sv2v_cast_0BC43('d2);
								2'b11: fpu_srcfmt_d = sv2v_cast_0BC43('d3);
							endcase
						end
						else
							case (operand_c_i[2:0])
								3'b000: fpu_srcfmt_d = sv2v_cast_0BC43('d0);
								3'b001: fpu_srcfmt_d = sv2v_cast_0BC43('d1);
								3'b010: fpu_srcfmt_d = sv2v_cast_0BC43('d2);
								3'b110: fpu_srcfmt_d = sv2v_cast_0BC43('d4);
								3'b011: fpu_srcfmt_d = sv2v_cast_0BC43('d3);
							endcase
					end
					7'd102: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = {1'b0, fpu_rm_i[1:0]};
						check_ah = 1'b1;
					end
					7'd103: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = 3'b011;
						fpu_op_mod_d = 1'b1;
						check_ah = 1'b1;
						vec_replication = 1'b0;
					end
					7'd104: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = 3'b011;
						check_ah = 1'b1;
						vec_replication = 1'b0;
					end
					7'd105: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_rm_d = {1'b0, fpu_rm_i[1:0]};
						check_ah = 1'b1;
					end
					7'd106: begin
						fpu_op_d = sv2v_cast_A53F3(9);
						fpu_rm_d = {1'b0, fpu_rm_i[1:0]};
						check_ah = 1'b1;
					end
					7'd107: begin
						fpu_op_d = sv2v_cast_A53F3(7);
						fpu_rm_d = 3'b000;
					end
					7'd108: begin
						fpu_op_d = sv2v_cast_A53F3(7);
						fpu_rm_d = 3'b001;
					end
					7'd109: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = 3'b000;
					end
					7'd110: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = 3'b001;
					end
					7'd111: begin
						fpu_op_d = sv2v_cast_A53F3(6);
						fpu_rm_d = 3'b010;
					end
					7'd112: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_rm_d = 3'b010;
					end
					7'd113: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_op_mod_d = 1'b1;
						fpu_rm_d = 3'b010;
					end
					7'd114: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_rm_d = 3'b001;
					end
					7'd115: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_op_mod_d = 1'b1;
						fpu_rm_d = 3'b001;
					end
					7'd116: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_rm_d = 3'b000;
					end
					7'd117: begin
						fpu_op_d = sv2v_cast_A53F3(8);
						fpu_op_mod_d = 1'b1;
						fpu_rm_d = 3'b000;
					end
					7'd118: begin
						fpu_op_d = sv2v_cast_A53F3(13);
						fpu_op_mod_d = fpu_rm_i[0];
						vec_replication = 1'b0;
						fpu_srcfmt_d = sv2v_cast_0BC43('d0);
					end
					7'd119: begin
						fpu_op_d = sv2v_cast_A53F3(14);
						fpu_op_mod_d = fpu_rm_i[0];
						vec_replication = 1'b0;
						fpu_srcfmt_d = sv2v_cast_0BC43('d0);
					end
					7'd120: begin
						fpu_op_d = sv2v_cast_A53F3(13);
						fpu_op_mod_d = fpu_rm_i[0];
						vec_replication = 1'b0;
						fpu_srcfmt_d = sv2v_cast_0BC43('d1);
					end
					7'd121: begin
						fpu_op_d = sv2v_cast_A53F3(14);
						fpu_op_mod_d = fpu_rm_i[0];
						vec_replication = 1'b0;
						fpu_srcfmt_d = sv2v_cast_0BC43('d1);
					end
					default:
						;
				endcase
				if (!fpu_vec_op_d && check_ah) begin
					if (fpu_rm_i[2])
						fpu_dstfmt_d = sv2v_cast_0BC43('d4);
				end
				if (fpu_vec_op_d && vec_replication) begin
					if (replicate_c)
						case (fpu_dstfmt_d)
							sv2v_cast_0BC43('d0): operand_c_d = (ariane_pkg_RVD ? {2 {operand_c_i[31:0]}} : operand_c_i);
							sv2v_cast_0BC43('d2), sv2v_cast_0BC43('d4): operand_c_d = (ariane_pkg_RVD ? {4 {operand_c_i[15:0]}} : {2 {operand_c_i[15:0]}});
							sv2v_cast_0BC43('d3): operand_c_d = (ariane_pkg_RVD ? {8 {operand_c_i[7:0]}} : {4 {operand_c_i[7:0]}});
						endcase
					else
						case (fpu_dstfmt_d)
							sv2v_cast_0BC43('d0): operand_b_d = (ariane_pkg_RVD ? {2 {operand_b_i[31:0]}} : operand_b_i);
							sv2v_cast_0BC43('d2), sv2v_cast_0BC43('d4): operand_b_d = (ariane_pkg_RVD ? {4 {operand_b_i[15:0]}} : {2 {operand_b_i[15:0]}});
							sv2v_cast_0BC43('d3): operand_b_d = (ariane_pkg_RVD ? {8 {operand_b_i[7:0]}} : {4 {operand_b_i[7:0]}});
						endcase
				end
			end
			always @(*) begin : p_inputFSM
				fpu_ready_o = 1'b0;
				fpu_in_valid = 1'b0;
				hold_inputs = 1'b0;
				use_hold = 1'b0;
				state_d = state_q;
				case (state_q)
					1'd0: begin
						fpu_ready_o = 1'b1;
						fpu_in_valid = fpu_valid_i;
						if (fpu_valid_i & ~fpu_in_ready) begin
							fpu_ready_o = 1'b0;
							hold_inputs = 1'b1;
							state_d = 1'd1;
						end
					end
					1'd1: begin
						fpu_in_valid = 1'b1;
						use_hold = 1'b1;
						if (fpu_in_ready) begin
							fpu_ready_o = 1'b1;
							state_d = 1'd0;
						end
					end
					default:
						;
				endcase
				if (flush_i)
					state_d = 1'd0;
			end
			always @(posedge clk_i or negedge rst_ni) begin : fp_hold_reg
				if (~rst_ni) begin
					state_q <= 1'd0;
					operand_a_q <= 1'sb0;
					operand_b_q <= 1'sb0;
					operand_c_q <= 1'sb0;
					fpu_op_q <= 1'sb0;
					fpu_op_mod_q <= 1'sb0;
					fpu_srcfmt_q <= 1'sb0;
					fpu_dstfmt_q <= 1'sb0;
					fpu_ifmt_q <= 1'sb0;
					fpu_rm_q <= 1'sb0;
					fpu_vec_op_q <= 1'sb0;
					fpu_tag_q <= 1'sb0;
				end
				else begin
					state_q <= state_d;
					if (hold_inputs) begin
						operand_a_q <= operand_a_d;
						operand_b_q <= operand_b_d;
						operand_c_q <= operand_c_d;
						fpu_op_q <= fpu_op_d;
						fpu_op_mod_q <= fpu_op_mod_d;
						fpu_srcfmt_q <= fpu_srcfmt_d;
						fpu_dstfmt_q <= fpu_dstfmt_d;
						fpu_ifmt_q <= fpu_ifmt_d;
						fpu_rm_q <= fpu_rm_d;
						fpu_vec_op_q <= fpu_vec_op_d;
						fpu_tag_q <= fpu_tag_d;
					end
				end
			end
			assign operand_a = (use_hold ? operand_a_q : operand_a_d);
			assign operand_b = (use_hold ? operand_b_q : operand_b_d);
			assign operand_c = (use_hold ? operand_c_q : operand_c_d);
			assign fpu_op = (use_hold ? fpu_op_q : fpu_op_d);
			assign fpu_op_mod = (use_hold ? fpu_op_mod_q : fpu_op_mod_d);
			assign fpu_srcfmt = (use_hold ? fpu_srcfmt_q : fpu_srcfmt_d);
			assign fpu_dstfmt = (use_hold ? fpu_dstfmt_q : fpu_dstfmt_d);
			assign fpu_ifmt = (use_hold ? fpu_ifmt_q : fpu_ifmt_d);
			assign fpu_rm = (use_hold ? fpu_rm_q : fpu_rm_d);
			assign fpu_vec_op = (use_hold ? fpu_vec_op_q : fpu_vec_op_d);
			assign fpu_tag = (use_hold ? fpu_tag_q : fpu_tag_d);
			wire [(3 * ariane_pkg_FLEN) - 1:0] fpu_operands;
			assign fpu_operands[0+:ariane_pkg_FLEN] = operand_a;
			assign fpu_operands[ariane_pkg_FLEN+:ariane_pkg_FLEN] = operand_b;
			assign fpu_operands[2 * ariane_pkg_FLEN+:ariane_pkg_FLEN] = operand_c;
			fpnew_top_60D59 #(
				.Features(FPU_FEATURES),
				.Implementation(FPU_IMPLEMENTATION)
			) i_fpnew_bulk(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(fpu_operands),
				.rnd_mode_i(fpu_rm),
				.op_i(sv2v_cast_A53F3(fpu_op)),
				.op_mod_i(fpu_op_mod),
				.src_fmt_i(sv2v_cast_0BC43(fpu_srcfmt)),
				.dst_fmt_i(sv2v_cast_0BC43(fpu_dstfmt)),
				.int_fmt_i(sv2v_cast_87CC5(fpu_ifmt)),
				.vectorial_op_i(fpu_vec_op),
				.tag_i(fpu_tag),
				.in_valid_i(fpu_in_valid),
				.in_ready_o(fpu_in_ready),
				.flush_i(flush_i),
				.result_o(result_o),
				.status_o(fpu_status),
				.tag_o(fpu_trans_id_o),
				.out_valid_o(fpu_out_valid),
				.out_ready_i(fpu_out_ready),
				.busy_o()
			);
			assign fpu_exception_o[128-:64] = {59'h000000000000000, fpu_status};
			assign fpu_exception_o[0] = 1'b0;
			assign fpu_out_ready = 1'b1;
			assign fpu_valid_o = fpu_out_valid;
		end
	endgenerate
endmodule
module id_stage (
	clk_i,
	rst_ni,
	flush_i,
	debug_req_i,
	fetch_entry_i,
	fetch_entry_valid_i,
	fetch_entry_ready_o,
	issue_entry_o,
	issue_entry_valid_o,
	is_ctrl_flow_o,
	issue_instr_ack_i,
	priv_lvl_i,
	fs_i,
	frm_i,
	irq_i,
	irq_ctrl_i,
	debug_mode_i,
	tvm_i,
	tw_i,
	tsr_i
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire debug_req_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [291:0] fetch_entry_i;
	input wire fetch_entry_valid_i;
	output reg fetch_entry_ready_o;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	output wire [360:0] issue_entry_o;
	output wire issue_entry_valid_o;
	output wire is_ctrl_flow_o;
	input wire issue_instr_ack_i;
	input wire [1:0] priv_lvl_i;
	input wire [1:0] fs_i;
	input wire [2:0] frm_i;
	input wire [1:0] irq_i;
	input wire [193:0] irq_ctrl_i;
	input wire debug_mode_i;
	input wire tvm_i;
	input wire tw_i;
	input wire tsr_i;
	reg [362:0] issue_n;
	reg [362:0] issue_q;
	wire is_control_flow_instr;
	wire [360:0] decoded_instruction;
	wire is_illegal;
	wire [31:0] instruction;
	wire is_compressed;
	compressed_decoder compressed_decoder_i(
		.instr_i(fetch_entry_i[227-:32]),
		.instr_o(instruction),
		.illegal_instr_o(is_illegal),
		.is_compressed_o(is_compressed)
	);
	decoder decoder_i(
		.debug_req_i(debug_req_i),
		.irq_ctrl_i(irq_ctrl_i),
		.irq_i(irq_i),
		.pc_i(fetch_entry_i[291-:64]),
		.is_compressed_i(is_compressed),
		.is_illegal_i(is_illegal),
		.instruction_i(instruction),
		.compressed_instr_i(fetch_entry_i[211:196]),
		.branch_predict_i(fetch_entry_i[195-:67]),
		.ex_i(fetch_entry_i[128-:129]),
		.priv_lvl_i(priv_lvl_i),
		.debug_mode_i(debug_mode_i),
		.fs_i(fs_i),
		.frm_i(frm_i),
		.tvm_i(tvm_i),
		.tw_i(tw_i),
		.tsr_i(tsr_i),
		.instruction_o(decoded_instruction),
		.is_control_flow_instr_o(is_control_flow_instr)
	);
	assign issue_entry_o = issue_q[361-:361];
	assign issue_entry_valid_o = issue_q[362];
	assign is_ctrl_flow_o = issue_q[0];
	always @(*) begin
		issue_n = issue_q;
		fetch_entry_ready_o = 1'b0;
		if (issue_instr_ack_i)
			issue_n[362] = 1'b0;
		if ((!issue_q[362] || issue_instr_ack_i) && fetch_entry_valid_i) begin
			fetch_entry_ready_o = 1'b1;
			issue_n = {1'b1, decoded_instruction, is_control_flow_instr};
		end
		if (flush_i)
			issue_n[362] = 1'b0;
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			issue_q <= 1'sb0;
		else
			issue_q <= issue_n;
endmodule
module instr_realign (
	clk_i,
	rst_ni,
	flush_i,
	valid_i,
	serving_unaligned_o,
	address_i,
	data_i,
	valid_o,
	addr_o,
	instr_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire valid_i;
	output wire serving_unaligned_o;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] address_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	input wire [31:0] data_i;
	localparam [31:0] ariane_pkg_INSTR_PER_FETCH = 2;
	output reg [1:0] valid_o;
	output reg [127:0] addr_o;
	output reg [63:0] instr_o;
	wire [3:0] instr_is_compressed;
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : genblk1
			assign instr_is_compressed[i] = ~&data_i[i * 16+:2];
		end
	endgenerate
	reg [15:0] unaligned_instr_d;
	reg [15:0] unaligned_instr_q;
	reg unaligned_d;
	reg unaligned_q;
	reg [63:0] unaligned_address_d;
	reg [63:0] unaligned_address_q;
	assign serving_unaligned_o = unaligned_q;
	generate
		if (1) begin : realign_bp_32
			always @(*) begin : re_align
				unaligned_d = unaligned_q;
				unaligned_address_d = {address_i[63:2], 2'b10};
				unaligned_instr_d = data_i[31:16];
				valid_o[0] = valid_i;
				instr_o[0+:32] = (unaligned_q ? {data_i[15:0], unaligned_instr_q} : data_i[31:0]);
				addr_o[0+:64] = (unaligned_q ? unaligned_address_q : address_i);
				valid_o[1] = 1'b0;
				instr_o[32+:32] = 1'sb0;
				addr_o[64+:64] = {address_i[63:2], 2'b10};
				if (instr_is_compressed[0] || unaligned_q) begin
					if (instr_is_compressed[1]) begin
						unaligned_d = 1'b0;
						valid_o[1] = valid_i;
						instr_o[32+:32] = {16'b0000000000000000, data_i[31:16]};
					end
					else begin
						unaligned_d = 1'b1;
						unaligned_instr_d = data_i[31:16];
						unaligned_address_d = {address_i[63:2], 2'b10};
					end
				end
				if (valid_i && address_i[1]) begin
					if (!instr_is_compressed[0]) begin
						valid_o = 1'sb0;
						unaligned_d = 1'b1;
						unaligned_address_d = {address_i[63:2], 2'b10};
						unaligned_instr_d = data_i[15:0];
					end
					else
						valid_o = 1'b1;
				end
			end
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			unaligned_q <= 1'b0;
			unaligned_address_q <= 1'sb0;
			unaligned_instr_q <= 1'sb0;
		end
		else begin
			if (valid_i) begin
				unaligned_address_q <= unaligned_address_d;
				unaligned_instr_q <= unaligned_instr_d;
			end
			if (flush_i)
				unaligned_q <= 1'b0;
			else if (valid_i)
				unaligned_q <= unaligned_d;
		end
endmodule
module issue_read_operands (
	clk_i,
	rst_ni,
	flush_i,
	issue_instr_i,
	issue_instr_valid_i,
	issue_ack_o,
	rs1_o,
	rs1_i,
	rs1_valid_i,
	rs2_o,
	rs2_i,
	rs2_valid_i,
	rs3_o,
	rs3_i,
	rs3_valid_i,
	rd_clobber_gpr_i,
	rd_clobber_fpr_i,
	fu_data_o,
	rs1_forwarding_o,
	rs2_forwarding_o,
	pc_o,
	is_compressed_instr_o,
	flu_ready_i,
	alu_valid_o,
	branch_valid_o,
	branch_predict_o,
	lsu_ready_i,
	lsu_valid_o,
	mult_valid_o,
	fpu_ready_i,
	fpu_valid_o,
	fpu_fmt_o,
	fpu_rm_o,
	csr_valid_o,
	waddr_i,
	wdata_i,
	we_gpr_i,
	we_fpr_i
);
	parameter [31:0] NR_COMMIT_PORTS = 2;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [360:0] issue_instr_i;
	input wire issue_instr_valid_i;
	output reg issue_ack_o;
	output reg [5:0] rs1_o;
	input wire [63:0] rs1_i;
	input wire rs1_valid_i;
	output reg [5:0] rs2_o;
	input wire [63:0] rs2_i;
	input wire rs2_valid_i;
	output reg [5:0] rs3_o;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam ariane_pkg_FLEN = (ariane_pkg_RVD ? 64 : (ariane_pkg_RVF ? 32 : (ariane_pkg_XF16 ? 16 : (ariane_pkg_XF16ALT ? 16 : (ariane_pkg_XF8 ? 8 : 1)))));
	input wire [ariane_pkg_FLEN - 1:0] rs3_i;
	input wire rs3_valid_i;
	input wire [255:0] rd_clobber_gpr_i;
	input wire [255:0] rd_clobber_fpr_i;
	output wire [205:0] fu_data_o;
	output wire [63:0] rs1_forwarding_o;
	output wire [63:0] rs2_forwarding_o;
	output reg [63:0] pc_o;
	output reg is_compressed_instr_o;
	input wire flu_ready_i;
	output wire alu_valid_o;
	output wire branch_valid_o;
	output reg [66:0] branch_predict_o;
	input wire lsu_ready_i;
	output wire lsu_valid_o;
	output wire mult_valid_o;
	input wire fpu_ready_i;
	output wire fpu_valid_o;
	output wire [1:0] fpu_fmt_o;
	output wire [2:0] fpu_rm_o;
	output wire csr_valid_o;
	input wire [(NR_COMMIT_PORTS * 5) - 1:0] waddr_i;
	input wire [(NR_COMMIT_PORTS * 64) - 1:0] wdata_i;
	input wire [NR_COMMIT_PORTS - 1:0] we_gpr_i;
	input wire [NR_COMMIT_PORTS - 1:0] we_fpr_i;
	reg stall;
	reg fu_busy;
	wire [63:0] operand_a_regfile;
	wire [63:0] operand_b_regfile;
	wire [ariane_pkg_FLEN - 1:0] operand_c_regfile;
	reg [63:0] operand_a_n;
	reg [63:0] operand_a_q;
	reg [63:0] operand_b_n;
	reg [63:0] operand_b_q;
	reg [63:0] imm_n;
	reg [63:0] imm_q;
	reg alu_valid_q;
	reg mult_valid_q;
	reg fpu_valid_q;
	reg [1:0] fpu_fmt_q;
	reg [2:0] fpu_rm_q;
	reg lsu_valid_q;
	reg csr_valid_q;
	reg branch_valid_q;
	reg [2:0] trans_id_n;
	reg [2:0] trans_id_q;
	reg [6:0] operator_n;
	reg [6:0] operator_q;
	reg [3:0] fu_n;
	reg [3:0] fu_q;
	reg forward_rs1;
	reg forward_rs2;
	reg forward_rs3;
	wire [31:0] orig_instr;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	assign orig_instr = sv2v_cast_32(issue_instr_i[100:69]);
	assign rs1_forwarding_o = operand_a_n[63:0];
	assign rs2_forwarding_o = operand_b_n[63:0];
	assign fu_data_o[194-:64] = operand_a_q;
	assign fu_data_o[130-:64] = operand_b_q;
	assign fu_data_o[205-:4] = fu_q;
	assign fu_data_o[201-:7] = operator_q;
	assign fu_data_o[2-:ariane_pkg_TRANS_ID_BITS] = trans_id_q;
	assign fu_data_o[66-:64] = imm_q;
	assign alu_valid_o = alu_valid_q;
	assign branch_valid_o = branch_valid_q;
	assign lsu_valid_o = lsu_valid_q;
	assign csr_valid_o = csr_valid_q;
	assign mult_valid_o = mult_valid_q;
	assign fpu_valid_o = fpu_valid_q;
	assign fpu_fmt_o = fpu_fmt_q;
	assign fpu_rm_o = fpu_rm_q;
	always @(*) begin : unit_busy
		case (issue_instr_i[293-:4])
			4'd0: fu_busy = 1'b0;
			4'd3, 4'd4, 4'd6, 4'd5: fu_busy = ~flu_ready_i;
			4'd7, 4'd8: fu_busy = ~fpu_ready_i;
			4'd1, 4'd2: fu_busy = ~lsu_ready_i;
			default: fu_busy = 1'b0;
		endcase
	end
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	function automatic ariane_pkg_is_imm_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd89 <= op) && (7'd90 >= op), (7'd95 <= op) && (7'd98 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_imm_fpr = 1'b1;
			else
				ariane_pkg_is_imm_fpr = 1'b0;
		end
		else
			ariane_pkg_is_imm_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs1_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd91 <= op) && (7'd98 >= op), op == 7'd99, op == 7'd101, op == 7'd102, op == 7'd103, op == 7'd105, op == 7'd106, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs1_fpr = 1'b1;
			else
				ariane_pkg_is_rs1_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs1_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs2_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd85 <= op) && (7'd88 >= op), (7'd89 <= op) && (7'd93 >= op), (7'd95 <= op) && (7'd98 >= op), op == 7'd101, (7'd102 <= op) && (7'd103 >= op), op == 7'd105, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs2_fpr = 1'b1;
			else
				ariane_pkg_is_rs2_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs2_fpr = 1'b0;
	endfunction
	always @(*) begin : operands_available
		stall = 1'b0;
		forward_rs1 = 1'b0;
		forward_rs2 = 1'b0;
		forward_rs3 = 1'b0;
		rs1_o = issue_instr_i[282-:6];
		rs2_o = issue_instr_i[276-:6];
		rs3_o = issue_instr_i[206:201];
		if (!issue_instr_i[198] && (ariane_pkg_is_rs1_fpr(issue_instr_i[289-:7]) ? rd_clobber_fpr_i[issue_instr_i[282-:6] * 4+:4] != 4'd0 : rd_clobber_gpr_i[issue_instr_i[282-:6] * 4+:4] != 4'd0)) begin
			if (rs1_valid_i && (ariane_pkg_is_rs1_fpr(issue_instr_i[289-:7]) ? 1'b1 : (rd_clobber_gpr_i[issue_instr_i[282-:6] * 4+:4] != 4'd6) || (issue_instr_i[289-:7] == 7'd30)))
				forward_rs1 = 1'b1;
			else
				stall = 1'b1;
		end
		if ((ariane_pkg_is_rs2_fpr(issue_instr_i[289-:7]) ? rd_clobber_fpr_i[issue_instr_i[276-:6] * 4+:4] != 4'd0 : rd_clobber_gpr_i[issue_instr_i[276-:6] * 4+:4] != 4'd0)) begin
			if (rs2_valid_i && (ariane_pkg_is_rs2_fpr(issue_instr_i[289-:7]) ? 1'b1 : (rd_clobber_gpr_i[issue_instr_i[276-:6] * 4+:4] != 4'd6) || (issue_instr_i[289-:7] == 7'd30)))
				forward_rs2 = 1'b1;
			else
				stall = 1'b1;
		end
		if (ariane_pkg_is_imm_fpr(issue_instr_i[289-:7]) && (rd_clobber_fpr_i[issue_instr_i[206:201] * 4+:4] != 4'd0)) begin
			if (rs3_valid_i)
				forward_rs3 = 1'b1;
			else
				stall = 1'b1;
		end
	end
	always @(*) begin : forwarding_operand_select
		operand_a_n = operand_a_regfile;
		operand_b_n = operand_b_regfile;
		imm_n = (ariane_pkg_is_imm_fpr(issue_instr_i[289-:7]) ? {{riscv_XLEN - ariane_pkg_FLEN {1'b0}}, operand_c_regfile} : issue_instr_i[264-:64]);
		trans_id_n = issue_instr_i[296-:3];
		fu_n = issue_instr_i[293-:4];
		operator_n = issue_instr_i[289-:7];
		if (forward_rs1)
			operand_a_n = rs1_i;
		if (forward_rs2)
			operand_b_n = rs2_i;
		if (forward_rs3)
			imm_n = {{riscv_XLEN - ariane_pkg_FLEN {1'b0}}, rs3_i};
		if (issue_instr_i[197])
			operand_a_n = {issue_instr_i[360-:64]};
		if (issue_instr_i[198])
			operand_a_n = {{59 {1'b0}}, issue_instr_i[281:277]};
		if (((issue_instr_i[199] && (issue_instr_i[293-:4] != 4'd2)) && (issue_instr_i[293-:4] != 4'd4)) && !ariane_pkg_is_rs2_fpr(issue_instr_i[289-:7]))
			operand_b_n = issue_instr_i[264-:64];
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			alu_valid_q <= 1'b0;
			lsu_valid_q <= 1'b0;
			mult_valid_q <= 1'b0;
			fpu_valid_q <= 1'b0;
			fpu_fmt_q <= 2'b00;
			fpu_rm_q <= 3'b000;
			csr_valid_q <= 1'b0;
			branch_valid_q <= 1'b0;
		end
		else begin
			alu_valid_q <= 1'b0;
			lsu_valid_q <= 1'b0;
			mult_valid_q <= 1'b0;
			fpu_valid_q <= 1'b0;
			fpu_fmt_q <= 2'b00;
			fpu_rm_q <= 3'b000;
			csr_valid_q <= 1'b0;
			branch_valid_q <= 1'b0;
			if ((!issue_instr_i[68] && issue_instr_valid_i) && issue_ack_o)
				case (issue_instr_i[293-:4])
					4'd3: alu_valid_q <= 1'b1;
					4'd4: branch_valid_q <= 1'b1;
					4'd5: mult_valid_q <= 1'b1;
					4'd7: begin
						fpu_valid_q <= 1'b1;
						fpu_fmt_q <= orig_instr[26-:2];
						fpu_rm_q <= orig_instr[14-:3];
					end
					4'd8: begin
						fpu_valid_q <= 1'b1;
						fpu_fmt_q <= orig_instr[13-:2];
						fpu_rm_q <= {2'b00, orig_instr[14]};
					end
					4'd1, 4'd2: lsu_valid_q <= 1'b1;
					4'd6: csr_valid_q <= 1'b1;
					default:
						;
				endcase
			if (flush_i) begin
				alu_valid_q <= 1'b0;
				lsu_valid_q <= 1'b0;
				mult_valid_q <= 1'b0;
				fpu_valid_q <= 1'b0;
				csr_valid_q <= 1'b0;
				branch_valid_q <= 1'b0;
			end
		end
	function automatic ariane_pkg_is_rd_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd81 <= op) && (7'd84 >= op), (7'd89 <= op) && (7'd98 >= op), op == 7'd100, op == 7'd101, op == 7'd102, op == 7'd104, (7'd107 <= op) && (7'd111 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rd_fpr = 1'b1;
			else
				ariane_pkg_is_rd_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rd_fpr = 1'b0;
	endfunction
	always @(*) begin : issue_scoreboard
		issue_ack_o = 1'b0;
		if (issue_instr_valid_i) begin
			if (!stall && !fu_busy) begin
				if ((ariane_pkg_is_rd_fpr(issue_instr_i[289-:7]) ? rd_clobber_fpr_i[issue_instr_i[270-:6] * 4+:4] == 4'd0 : rd_clobber_gpr_i[issue_instr_i[270-:6] * 4+:4] == 4'd0))
					issue_ack_o = 1'b1;
				begin : sv2v_autoblock_1
					reg [31:0] i;
					for (i = 0; i < NR_COMMIT_PORTS; i = i + 1)
						if ((ariane_pkg_is_rd_fpr(issue_instr_i[289-:7]) ? we_fpr_i[i] && (waddr_i[i * 5+:5] == issue_instr_i[270-:6]) : we_gpr_i[i] && (waddr_i[i * 5+:5] == issue_instr_i[270-:6])))
							issue_ack_o = 1'b1;
				end
			end
			if (issue_instr_i[68])
				issue_ack_o = 1'b1;
			if (issue_instr_i[293-:4] == 4'd0)
				issue_ack_o = 1'b1;
		end
		if (mult_valid_q && (issue_instr_i[293-:4] != 4'd5))
			issue_ack_o = 1'b0;
	end
	wire [127:0] rdata;
	wire [9:0] raddr_pack;
	wire [(NR_COMMIT_PORTS * 5) - 1:0] waddr_pack;
	wire [(NR_COMMIT_PORTS * 64) - 1:0] wdata_pack;
	wire [NR_COMMIT_PORTS - 1:0] we_pack;
	assign raddr_pack = {issue_instr_i[275:271], issue_instr_i[281:277]};
	genvar i;
	generate
		for (i = 0; i < NR_COMMIT_PORTS; i = i + 1) begin : gen_write_back_port
			assign waddr_pack[i * 5+:5] = waddr_i[i * 5+:5];
			assign wdata_pack[i * 64+:64] = wdata_i[i * 64+:64];
			assign we_pack[i] = we_gpr_i[i];
		end
	endgenerate
	ariane_regfile #(
		.DATA_WIDTH(riscv_XLEN),
		.NR_READ_PORTS(2),
		.NR_WRITE_PORTS(NR_COMMIT_PORTS),
		.ZERO_REG_ZERO(1)
	) i_ariane_regfile(
		.test_en_i(1'b0),
		.raddr_i(raddr_pack),
		.rdata_o(rdata),
		.waddr_i(waddr_pack),
		.wdata_i(wdata_pack),
		.we_i(we_pack),
		.clk_i(clk_i),
		.rst_ni(rst_ni)
	);
	wire [(3 * ariane_pkg_FLEN) - 1:0] fprdata;
	wire [14:0] fp_raddr_pack;
	wire [(NR_COMMIT_PORTS * 64) - 1:0] fp_wdata_pack;
	function automatic [ariane_pkg_FLEN - 1:0] sv2v_cast_83D81;
		input reg [ariane_pkg_FLEN - 1:0] inp;
		sv2v_cast_83D81 = inp;
	endfunction
	generate
		if (ariane_pkg_FP_PRESENT) begin : float_regfile_gen
			assign fp_raddr_pack = {issue_instr_i[205:201], issue_instr_i[275:271], issue_instr_i[281:277]};
			genvar i;
			for (i = 0; i < NR_COMMIT_PORTS; i = i + 1) begin : gen_fp_wdata_pack
				assign fp_wdata_pack[i * 64+:64] = {wdata_i[(i * 64) + (ariane_pkg_FLEN - 1)-:ariane_pkg_FLEN]};
			end
			ariane_regfile #(
				.DATA_WIDTH(ariane_pkg_FLEN),
				.NR_READ_PORTS(3),
				.NR_WRITE_PORTS(NR_COMMIT_PORTS),
				.ZERO_REG_ZERO(0)
			) i_ariane_fp_regfile(
				.test_en_i(1'b0),
				.raddr_i(fp_raddr_pack),
				.rdata_o(fprdata),
				.waddr_i(waddr_pack),
				.wdata_i(wdata_pack),
				.we_i(we_fpr_i),
				.clk_i(clk_i),
				.rst_ni(rst_ni)
			);
		end
		else begin : no_fpr_gen
			assign fprdata = {3 {sv2v_cast_83D81(1'sb0)}};
		end
	endgenerate
	assign operand_a_regfile = (ariane_pkg_is_rs1_fpr(issue_instr_i[289-:7]) ? {{riscv_XLEN - ariane_pkg_FLEN {1'b0}}, fprdata[0+:ariane_pkg_FLEN]} : rdata[0+:64]);
	assign operand_b_regfile = (ariane_pkg_is_rs2_fpr(issue_instr_i[289-:7]) ? {{riscv_XLEN - ariane_pkg_FLEN {1'b0}}, fprdata[ariane_pkg_FLEN+:ariane_pkg_FLEN]} : rdata[64+:64]);
	assign operand_c_regfile = fprdata[2 * ariane_pkg_FLEN+:ariane_pkg_FLEN];
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			operand_a_q <= {riscv_XLEN {1'd0}};
			operand_b_q <= {riscv_XLEN {1'd0}};
			imm_q <= 1'sb0;
			fu_q <= 4'd0;
			operator_q <= 7'd0;
			trans_id_q <= 1'sb0;
			pc_o <= 1'sb0;
			is_compressed_instr_o <= 1'b0;
			branch_predict_o <= {3'd0, {riscv_VLEN {1'b0}}};
		end
		else begin
			operand_a_q <= operand_a_n;
			operand_b_q <= operand_b_n;
			imm_q <= imm_n;
			fu_q <= fu_n;
			operator_q <= operator_n;
			trans_id_q <= trans_id_n;
			pc_o <= issue_instr_i[360-:64];
			is_compressed_instr_o <= issue_instr_i[0];
			branch_predict_o <= issue_instr_i[67-:67];
		end
endmodule
module issue_stage (
	clk_i,
	rst_ni,
	sb_full_o,
	flush_unissued_instr_i,
	flush_i,
	decoded_instr_i,
	decoded_instr_valid_i,
	is_ctrl_flow_i,
	decoded_instr_ack_o,
	rs1_forwarding_o,
	rs2_forwarding_o,
	fu_data_o,
	pc_o,
	is_compressed_instr_o,
	flu_ready_i,
	alu_valid_o,
	resolve_branch_i,
	lsu_ready_i,
	lsu_valid_o,
	branch_valid_o,
	branch_predict_o,
	mult_valid_o,
	fpu_ready_i,
	fpu_valid_o,
	fpu_fmt_o,
	fpu_rm_o,
	csr_valid_o,
	trans_id_i,
	resolved_branch_i,
	wbdata_i,
	ex_ex_i,
	wt_valid_i,
	waddr_i,
	wdata_i,
	we_gpr_i,
	we_fpr_i,
	commit_instr_o,
	commit_ack_i
);
	parameter [31:0] NR_ENTRIES = 8;
	parameter [31:0] NR_WB_PORTS = 4;
	parameter [31:0] NR_COMMIT_PORTS = 2;
	input wire clk_i;
	input wire rst_ni;
	output wire sb_full_o;
	input wire flush_unissued_instr_i;
	input wire flush_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [360:0] decoded_instr_i;
	input wire decoded_instr_valid_i;
	input wire is_ctrl_flow_i;
	output wire decoded_instr_ack_o;
	output wire [63:0] rs1_forwarding_o;
	output wire [63:0] rs2_forwarding_o;
	output wire [205:0] fu_data_o;
	output wire [63:0] pc_o;
	output wire is_compressed_instr_o;
	input wire flu_ready_i;
	output wire alu_valid_o;
	input wire resolve_branch_i;
	input wire lsu_ready_i;
	output wire lsu_valid_o;
	output wire branch_valid_o;
	output wire [66:0] branch_predict_o;
	output wire mult_valid_o;
	input wire fpu_ready_i;
	output wire fpu_valid_o;
	output wire [1:0] fpu_fmt_o;
	output wire [2:0] fpu_rm_o;
	output wire csr_valid_o;
	input wire [(NR_WB_PORTS * 3) - 1:0] trans_id_i;
	input wire [133:0] resolved_branch_i;
	input wire [(NR_WB_PORTS * 64) - 1:0] wbdata_i;
	input wire [(NR_WB_PORTS * 129) - 1:0] ex_ex_i;
	input wire [NR_WB_PORTS - 1:0] wt_valid_i;
	input wire [(NR_COMMIT_PORTS * 5) - 1:0] waddr_i;
	input wire [(NR_COMMIT_PORTS * 64) - 1:0] wdata_i;
	input wire [NR_COMMIT_PORTS - 1:0] we_gpr_i;
	input wire [NR_COMMIT_PORTS - 1:0] we_fpr_i;
	output wire [(NR_COMMIT_PORTS * 361) - 1:0] commit_instr_o;
	input wire [NR_COMMIT_PORTS - 1:0] commit_ack_i;
	wire [255:0] rd_clobber_gpr_sb_iro;
	wire [255:0] rd_clobber_fpr_sb_iro;
	wire [5:0] rs1_iro_sb;
	wire [63:0] rs1_sb_iro;
	wire rs1_valid_sb_iro;
	wire [5:0] rs2_iro_sb;
	wire [63:0] rs2_sb_iro;
	wire rs2_valid_iro_sb;
	wire [5:0] rs3_iro_sb;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam ariane_pkg_FLEN = (ariane_pkg_RVD ? 64 : (ariane_pkg_RVF ? 32 : (ariane_pkg_XF16 ? 16 : (ariane_pkg_XF16ALT ? 16 : (ariane_pkg_XF8 ? 8 : 1)))));
	wire [ariane_pkg_FLEN - 1:0] rs3_sb_iro;
	wire rs3_valid_iro_sb;
	wire [360:0] issue_instr_rename_sb;
	wire issue_instr_valid_rename_sb;
	wire issue_ack_sb_rename;
	wire [360:0] issue_instr_sb_iro;
	wire issue_instr_valid_sb_iro;
	wire issue_ack_iro_sb;
	re_name i_re_name(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.flush_unissied_instr_i(flush_unissued_instr_i),
		.issue_instr_i(decoded_instr_i),
		.issue_instr_valid_i(decoded_instr_valid_i),
		.issue_ack_o(decoded_instr_ack_o),
		.issue_instr_o(issue_instr_rename_sb),
		.issue_instr_valid_o(issue_instr_valid_rename_sb),
		.issue_ack_i(issue_ack_sb_rename)
	);
	scoreboard #(
		.NR_ENTRIES(NR_ENTRIES),
		.NR_WB_PORTS(NR_WB_PORTS),
		.NR_COMMIT_PORTS(NR_COMMIT_PORTS)
	) i_scoreboard(
		.sb_full_o(sb_full_o),
		.unresolved_branch_i(1'b0),
		.rd_clobber_gpr_o(rd_clobber_gpr_sb_iro),
		.rd_clobber_fpr_o(rd_clobber_fpr_sb_iro),
		.rs1_i(rs1_iro_sb),
		.rs1_o(rs1_sb_iro),
		.rs1_valid_o(rs1_valid_sb_iro),
		.rs2_i(rs2_iro_sb),
		.rs2_o(rs2_sb_iro),
		.rs2_valid_o(rs2_valid_iro_sb),
		.rs3_i(rs3_iro_sb),
		.rs3_o(rs3_sb_iro),
		.rs3_valid_o(rs3_valid_iro_sb),
		.decoded_instr_i(issue_instr_rename_sb),
		.decoded_instr_valid_i(issue_instr_valid_rename_sb),
		.decoded_instr_ack_o(issue_ack_sb_rename),
		.issue_instr_o(issue_instr_sb_iro),
		.issue_instr_valid_o(issue_instr_valid_sb_iro),
		.issue_ack_i(issue_ack_iro_sb),
		.resolved_branch_i(resolved_branch_i),
		.trans_id_i(trans_id_i),
		.wbdata_i(wbdata_i),
		.ex_i(ex_ex_i),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_unissued_instr_i(flush_unissued_instr_i),
		.flush_i(flush_i),
		.commit_instr_o(commit_instr_o),
		.commit_ack_i(commit_ack_i),
		.wt_valid_i(wt_valid_i)
	);
	issue_read_operands #(.NR_COMMIT_PORTS(NR_COMMIT_PORTS)) i_issue_read_operands(
		.flush_i(flush_unissued_instr_i),
		.issue_instr_i(issue_instr_sb_iro),
		.issue_instr_valid_i(issue_instr_valid_sb_iro),
		.issue_ack_o(issue_ack_iro_sb),
		.fu_data_o(fu_data_o),
		.flu_ready_i(flu_ready_i),
		.rs1_o(rs1_iro_sb),
		.rs1_i(rs1_sb_iro),
		.rs1_valid_i(rs1_valid_sb_iro),
		.rs2_o(rs2_iro_sb),
		.rs2_i(rs2_sb_iro),
		.rs2_valid_i(rs2_valid_iro_sb),
		.rs3_o(rs3_iro_sb),
		.rs3_i(rs3_sb_iro),
		.rs3_valid_i(rs3_valid_iro_sb),
		.rd_clobber_gpr_i(rd_clobber_gpr_sb_iro),
		.rd_clobber_fpr_i(rd_clobber_fpr_sb_iro),
		.alu_valid_o(alu_valid_o),
		.branch_valid_o(branch_valid_o),
		.csr_valid_o(csr_valid_o),
		.mult_valid_o(mult_valid_o),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rs1_forwarding_o(rs1_forwarding_o),
		.rs2_forwarding_o(rs2_forwarding_o),
		.pc_o(pc_o),
		.is_compressed_instr_o(is_compressed_instr_o),
		.branch_predict_o(branch_predict_o),
		.lsu_ready_i(lsu_ready_i),
		.lsu_valid_o(lsu_valid_o),
		.fpu_ready_i(fpu_ready_i),
		.fpu_valid_o(fpu_valid_o),
		.fpu_fmt_o(fpu_fmt_o),
		.fpu_rm_o(fpu_rm_o),
		.waddr_i(waddr_i),
		.wdata_i(wdata_i),
		.we_gpr_i(we_gpr_i),
		.we_fpr_i(we_fpr_i)
	);
endmodule
module load_store_unit (
	clk_i,
	rst_ni,
	flush_i,
	no_st_pending_o,
	amo_valid_commit_i,
	fu_data_i,
	lsu_ready_o,
	lsu_valid_i,
	load_trans_id_o,
	load_result_o,
	load_valid_o,
	load_exception_o,
	store_trans_id_o,
	store_result_o,
	store_valid_o,
	store_exception_o,
	commit_i,
	commit_ready_o,
	commit_tran_id_i,
	enable_translation_i,
	en_ld_st_translation_i,
	icache_areq_i,
	icache_areq_o,
	priv_lvl_i,
	ld_st_priv_lvl_i,
	sum_i,
	mxr_i,
	satp_ppn_i,
	asid_i,
	asid_to_be_flushed_i,
	vaddr_to_be_flushed_i,
	flush_tlb_i,
	itlb_miss_o,
	dtlb_miss_o,
	dcache_req_ports_i,
	dcache_req_ports_o,
	dcache_wbuffer_empty_i,
	dcache_wbuffer_not_ni_i,
	amo_req_o,
	amo_resp_i,
	pmpcfg_i,
	pmpaddr_i
);
	parameter [31:0] ASID_WIDTH = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	output wire no_st_pending_o;
	input wire amo_valid_commit_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	output wire lsu_ready_o;
	input wire lsu_valid_i;
	output wire [2:0] load_trans_id_o;
	output wire [63:0] load_result_o;
	output wire load_valid_o;
	output wire [128:0] load_exception_o;
	output wire [2:0] store_trans_id_o;
	output wire [63:0] store_result_o;
	output wire store_valid_o;
	output wire [128:0] store_exception_o;
	input wire commit_i;
	output wire commit_ready_o;
	input wire [2:0] commit_tran_id_i;
	input wire enable_translation_i;
	input wire en_ld_st_translation_i;
	localparam riscv_VLEN = 64;
	input wire [64:0] icache_areq_i;
	localparam riscv_PLEN = 56;
	output wire [185:0] icache_areq_o;
	input wire [1:0] priv_lvl_i;
	input wire [1:0] ld_st_priv_lvl_i;
	input wire sum_i;
	input wire mxr_i;
	localparam riscv_PPNW = 44;
	input wire [43:0] satp_ppn_i;
	input wire [ASID_WIDTH - 1:0] asid_i;
	input wire [ASID_WIDTH - 1:0] asid_to_be_flushed_i;
	input wire [63:0] vaddr_to_be_flushed_i;
	input wire flush_tlb_i;
	output wire itlb_miss_o;
	output wire dtlb_miss_o;
	input wire [197:0] dcache_req_ports_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (3 * ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78)) - 1 : (3 * (1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 76)):(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)] dcache_req_ports_o;
	input wire dcache_wbuffer_empty_i;
	input wire dcache_wbuffer_not_ni_i;
	output wire [134:0] amo_req_o;
	input wire [64:0] amo_resp_i;
	input wire [127:0] pmpcfg_i;
	input wire [863:0] pmpaddr_i;
	reg data_misaligned;
	wire [151:0] lsu_ctrl;
	wire pop_st;
	wire pop_ld;
	wire [63:0] vaddr_i;
	wire [63:0] vaddr_xlen;
	wire overflow;
	wire [7:0] be_i;
	assign vaddr_xlen = $unsigned($signed(fu_data_i[66-:64]) + $signed(fu_data_i[194-:64]));
	assign vaddr_i = vaddr_xlen[63:0];
	localparam [3:0] riscv_MODE_SV = 4'd8;
	localparam riscv_SV = 39;
	assign overflow = !((&vaddr_xlen[63:38] == 1'b1) || (|vaddr_xlen[63:38] == 1'b0));
	reg st_valid_i;
	reg ld_valid_i;
	wire ld_translation_req;
	wire st_translation_req;
	wire [63:0] ld_vaddr;
	wire [63:0] st_vaddr;
	reg translation_req;
	wire translation_valid;
	reg [63:0] mmu_vaddr;
	wire [55:0] mmu_paddr;
	wire [128:0] mmu_exception;
	wire dtlb_hit;
	wire [43:0] dtlb_ppn;
	wire ld_valid;
	wire [2:0] ld_trans_id;
	wire [63:0] ld_result;
	wire st_valid;
	wire [2:0] st_trans_id;
	wire [63:0] st_result;
	wire [11:0] page_offset;
	wire page_offset_matches;
	reg [128:0] misaligned_exception;
	wire [128:0] ld_ex;
	wire [128:0] st_ex;
	mmu #(
		.INSTR_TLB_ENTRIES(16),
		.DATA_TLB_ENTRIES(16),
		.ASID_WIDTH(ASID_WIDTH),
		.ArianeCfg(ArianeCfg)
	) i_mmu(
		.misaligned_ex_i(misaligned_exception),
		.lsu_is_store_i(st_translation_req),
		.lsu_req_i(translation_req),
		.lsu_vaddr_i(mmu_vaddr),
		.lsu_valid_o(translation_valid),
		.lsu_paddr_o(mmu_paddr),
		.lsu_exception_o(mmu_exception),
		.lsu_dtlb_hit_o(dtlb_hit),
		.lsu_dtlb_ppn_o(dtlb_ppn),
		.req_port_i(dcache_req_ports_i[0+:66]),
		.req_port_o(dcache_req_ports_o[(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) + 0+:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))]),
		.icache_areq_i(icache_areq_i),
		.asid_to_be_flushed_i(asid_to_be_flushed_i),
		.vaddr_to_be_flushed_i(vaddr_to_be_flushed_i),
		.icache_areq_o(icache_areq_o),
		.pmpcfg_i(pmpcfg_i),
		.pmpaddr_i(pmpaddr_i),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.enable_translation_i(enable_translation_i),
		.en_ld_st_translation_i(en_ld_st_translation_i),
		.priv_lvl_i(priv_lvl_i),
		.ld_st_priv_lvl_i(ld_st_priv_lvl_i),
		.sum_i(sum_i),
		.mxr_i(mxr_i),
		.satp_ppn_i(satp_ppn_i),
		.asid_i(asid_i),
		.flush_tlb_i(flush_tlb_i),
		.itlb_miss_o(itlb_miss_o),
		.dtlb_miss_o(dtlb_miss_o)
	);
	wire store_buffer_empty;
	store_unit i_store_unit(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.no_st_pending_o(no_st_pending_o),
		.store_buffer_empty_o(store_buffer_empty),
		.valid_i(st_valid_i),
		.lsu_ctrl_i(lsu_ctrl),
		.pop_st_o(pop_st),
		.commit_i(commit_i),
		.commit_ready_o(commit_ready_o),
		.amo_valid_commit_i(amo_valid_commit_i),
		.valid_o(st_valid),
		.trans_id_o(st_trans_id),
		.result_o(st_result),
		.ex_o(st_ex),
		.translation_req_o(st_translation_req),
		.vaddr_o(st_vaddr),
		.paddr_i(mmu_paddr),
		.ex_i(mmu_exception),
		.dtlb_hit_i(dtlb_hit),
		.page_offset_i(page_offset),
		.page_offset_matches_o(page_offset_matches),
		.amo_req_o(amo_req_o),
		.amo_resp_i(amo_resp_i),
		.req_port_i(dcache_req_ports_i[132+:66]),
		.req_port_o(dcache_req_ports_o[(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) + (2 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)))+:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))])
	);
	load_unit #(.ArianeCfg(ArianeCfg)) i_load_unit(
		.valid_i(ld_valid_i),
		.lsu_ctrl_i(lsu_ctrl),
		.pop_ld_o(pop_ld),
		.valid_o(ld_valid),
		.trans_id_o(ld_trans_id),
		.result_o(ld_result),
		.ex_o(ld_ex),
		.translation_req_o(ld_translation_req),
		.vaddr_o(ld_vaddr),
		.paddr_i(mmu_paddr),
		.ex_i(mmu_exception),
		.dtlb_hit_i(dtlb_hit),
		.dtlb_ppn_i(dtlb_ppn),
		.page_offset_o(page_offset),
		.page_offset_matches_i(page_offset_matches),
		.store_buffer_empty_i(store_buffer_empty),
		.req_port_i(dcache_req_ports_i[66+:66]),
		.req_port_o(dcache_req_ports_o[(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) + (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))+:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))]),
		.dcache_wbuffer_not_ni_i(dcache_wbuffer_not_ni_i),
		.commit_tran_id_i(commit_tran_id_i),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i)
	);
	localparam [31:0] ariane_pkg_NR_LOAD_PIPE_REGS = 1;
	shift_reg_1F3E0_50B1B #(
		.dtype_riscv_XLEN(riscv_XLEN),
		.Depth(ariane_pkg_NR_LOAD_PIPE_REGS)
	) i_pipe_reg_load(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({ld_valid, ld_trans_id, ld_result, ld_ex}),
		.d_o({load_valid_o, load_trans_id_o, load_result_o, load_exception_o})
	);
	localparam [31:0] ariane_pkg_NR_STORE_PIPE_REGS = 0;
	shift_reg_1F3E0_50B1B #(
		.dtype_riscv_XLEN(riscv_XLEN),
		.Depth(ariane_pkg_NR_STORE_PIPE_REGS)
	) i_pipe_reg_store(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.d_i({st_valid, st_trans_id, st_result, st_ex}),
		.d_o({store_valid_o, store_trans_id_o, store_result_o, store_exception_o})
	);
	always @(*) begin : which_op
		ld_valid_i = 1'b0;
		st_valid_i = 1'b0;
		translation_req = 1'b0;
		mmu_vaddr = {riscv_VLEN {1'b0}};
		case (lsu_ctrl[13-:4])
			4'd1: begin
				ld_valid_i = lsu_ctrl[151];
				translation_req = ld_translation_req;
				mmu_vaddr = ld_vaddr;
			end
			4'd2: begin
				st_valid_i = lsu_ctrl[151];
				translation_req = st_translation_req;
				mmu_vaddr = st_vaddr;
			end
			default:
				;
		endcase
	end
	function automatic [7:0] ariane_pkg_be_gen;
		input reg [2:0] addr;
		input reg [1:0] size;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			case (size)
				2'b11: begin
					ariane_pkg_be_gen = 8'b11111111;
					_sv2v_jump = 2'b11;
				end
				2'b10:
					case (addr[2:0])
						3'b000: begin
							ariane_pkg_be_gen = 8'b00001111;
							_sv2v_jump = 2'b11;
						end
						3'b001: begin
							ariane_pkg_be_gen = 8'b00011110;
							_sv2v_jump = 2'b11;
						end
						3'b010: begin
							ariane_pkg_be_gen = 8'b00111100;
							_sv2v_jump = 2'b11;
						end
						3'b011: begin
							ariane_pkg_be_gen = 8'b01111000;
							_sv2v_jump = 2'b11;
						end
						3'b100: begin
							ariane_pkg_be_gen = 8'b11110000;
							_sv2v_jump = 2'b11;
						end
					endcase
				2'b01:
					case (addr[2:0])
						3'b000: begin
							ariane_pkg_be_gen = 8'b00000011;
							_sv2v_jump = 2'b11;
						end
						3'b001: begin
							ariane_pkg_be_gen = 8'b00000110;
							_sv2v_jump = 2'b11;
						end
						3'b010: begin
							ariane_pkg_be_gen = 8'b00001100;
							_sv2v_jump = 2'b11;
						end
						3'b011: begin
							ariane_pkg_be_gen = 8'b00011000;
							_sv2v_jump = 2'b11;
						end
						3'b100: begin
							ariane_pkg_be_gen = 8'b00110000;
							_sv2v_jump = 2'b11;
						end
						3'b101: begin
							ariane_pkg_be_gen = 8'b01100000;
							_sv2v_jump = 2'b11;
						end
						3'b110: begin
							ariane_pkg_be_gen = 8'b11000000;
							_sv2v_jump = 2'b11;
						end
					endcase
				2'b00:
					case (addr[2:0])
						3'b000: begin
							ariane_pkg_be_gen = 8'b00000001;
							_sv2v_jump = 2'b11;
						end
						3'b001: begin
							ariane_pkg_be_gen = 8'b00000010;
							_sv2v_jump = 2'b11;
						end
						3'b010: begin
							ariane_pkg_be_gen = 8'b00000100;
							_sv2v_jump = 2'b11;
						end
						3'b011: begin
							ariane_pkg_be_gen = 8'b00001000;
							_sv2v_jump = 2'b11;
						end
						3'b100: begin
							ariane_pkg_be_gen = 8'b00010000;
							_sv2v_jump = 2'b11;
						end
						3'b101: begin
							ariane_pkg_be_gen = 8'b00100000;
							_sv2v_jump = 2'b11;
						end
						3'b110: begin
							ariane_pkg_be_gen = 8'b01000000;
							_sv2v_jump = 2'b11;
						end
						3'b111: begin
							ariane_pkg_be_gen = 8'b10000000;
							_sv2v_jump = 2'b11;
						end
					endcase
			endcase
			if (_sv2v_jump == 2'b00) begin
				ariane_pkg_be_gen = 8'b00000000;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [1:0] ariane_pkg_extract_transfer_size;
		input reg [6:0] op;
		case (op)
			7'd35, 7'd36, 7'd81, 7'd85, 7'd47, 7'd49, 7'd59, 7'd60, 7'd61, 7'd62, 7'd63, 7'd64, 7'd65, 7'd66, 7'd67: ariane_pkg_extract_transfer_size = 2'b11;
			7'd37, 7'd38, 7'd39, 7'd82, 7'd86, 7'd46, 7'd48, 7'd50, 7'd51, 7'd52, 7'd53, 7'd54, 7'd55, 7'd56, 7'd57, 7'd58: ariane_pkg_extract_transfer_size = 2'b10;
			7'd40, 7'd41, 7'd42, 7'd83, 7'd87: ariane_pkg_extract_transfer_size = 2'b01;
			7'd43, 7'd45, 7'd44, 7'd84, 7'd88: ariane_pkg_extract_transfer_size = 2'b00;
			default: ariane_pkg_extract_transfer_size = 2'b11;
		endcase
	endfunction
	assign be_i = ariane_pkg_be_gen(vaddr_i[2:0], ariane_pkg_extract_transfer_size(fu_data_i[201-:7]));
	localparam [63:0] riscv_LD_ACCESS_FAULT = 5;
	localparam [63:0] riscv_LD_ADDR_MISALIGNED = 4;
	localparam [63:0] riscv_ST_ACCESS_FAULT = 7;
	localparam [63:0] riscv_ST_ADDR_MISALIGNED = 6;
	always @(*) begin : data_misaligned_detection
		misaligned_exception = {{riscv_XLEN {1'b0}}, {riscv_XLEN {1'b0}}, 1'b0};
		data_misaligned = 1'b0;
		if (lsu_ctrl[151])
			case (lsu_ctrl[9-:7])
				7'd35, 7'd36, 7'd81, 7'd85, 7'd47, 7'd49, 7'd59, 7'd60, 7'd61, 7'd62, 7'd63, 7'd64, 7'd65, 7'd66, 7'd67:
					if (lsu_ctrl[89:87] != 3'b000)
						data_misaligned = 1'b1;
				7'd37, 7'd38, 7'd39, 7'd82, 7'd86, 7'd46, 7'd48, 7'd50, 7'd51, 7'd52, 7'd53, 7'd54, 7'd55, 7'd56, 7'd57, 7'd58:
					if (lsu_ctrl[88:87] != 2'b00)
						data_misaligned = 1'b1;
				7'd40, 7'd41, 7'd42, 7'd83, 7'd87:
					if (lsu_ctrl[87] != 1'b0)
						data_misaligned = 1'b1;
				default:
					;
			endcase
		if (data_misaligned) begin
			if (lsu_ctrl[13-:4] == 4'd1)
				misaligned_exception = {riscv_LD_ADDR_MISALIGNED, lsu_ctrl[150-:64], 1'b1};
			else if (lsu_ctrl[13-:4] == 4'd2)
				misaligned_exception = {riscv_ST_ADDR_MISALIGNED, lsu_ctrl[150-:64], 1'b1};
		end
		if (en_ld_st_translation_i && lsu_ctrl[86]) begin
			if (lsu_ctrl[13-:4] == 4'd1)
				misaligned_exception = {riscv_LD_ACCESS_FAULT, lsu_ctrl[150-:64], 1'b1};
			else if (lsu_ctrl[13-:4] == 4'd2)
				misaligned_exception = {riscv_ST_ACCESS_FAULT, lsu_ctrl[150-:64], 1'b1};
		end
	end
	wire [151:0] lsu_req_i;
	assign lsu_req_i = {lsu_valid_i, vaddr_i, overflow, fu_data_i[130-:64], be_i, fu_data_i[205-:4], fu_data_i[201-:7], fu_data_i[2-:ariane_pkg_TRANS_ID_BITS]};
	lsu_bypass lsu_bypass_i(
		.lsu_req_i(lsu_req_i),
		.lus_req_valid_i(lsu_valid_i),
		.pop_ld_i(pop_ld),
		.pop_st_i(pop_st),
		.lsu_ctrl_o(lsu_ctrl),
		.ready_o(lsu_ready_o),
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i)
	);
endmodule
module lsu_bypass (
	clk_i,
	rst_ni,
	flush_i,
	lsu_req_i,
	lus_req_valid_i,
	pop_ld_i,
	pop_st_i,
	lsu_ctrl_o,
	ready_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [151:0] lsu_req_i;
	input wire lus_req_valid_i;
	input wire pop_ld_i;
	input wire pop_st_i;
	output reg [151:0] lsu_ctrl_o;
	output wire ready_o;
	reg [303:0] mem_n;
	reg [303:0] mem_q;
	reg read_pointer_n;
	reg read_pointer_q;
	reg write_pointer_n;
	reg write_pointer_q;
	reg [1:0] status_cnt_n;
	reg [1:0] status_cnt_q;
	wire empty;
	assign empty = status_cnt_q == 0;
	assign ready_o = empty;
	always @(*) begin : sv2v_autoblock_1
		reg [1:0] status_cnt;
		reg write_pointer;
		reg read_pointer;
		status_cnt = status_cnt_q;
		write_pointer = write_pointer_q;
		read_pointer = read_pointer_q;
		mem_n = mem_q;
		if (lus_req_valid_i) begin
			mem_n[write_pointer_q * 152+:152] = lsu_req_i;
			write_pointer = write_pointer + 1;
			status_cnt = status_cnt + 1;
		end
		if (pop_ld_i) begin
			mem_n[(read_pointer_q * 152) + 151] = 1'b0;
			read_pointer = read_pointer + 1;
			status_cnt = status_cnt - 1;
		end
		if (pop_st_i) begin
			mem_n[(read_pointer_q * 152) + 151] = 1'b0;
			read_pointer = read_pointer + 1;
			status_cnt = status_cnt - 1;
		end
		if (pop_st_i && pop_ld_i)
			mem_n = 1'sb0;
		if (flush_i) begin
			status_cnt = 1'sb0;
			write_pointer = 1'sb0;
			read_pointer = 1'sb0;
			mem_n = 1'sb0;
		end
		read_pointer_n = read_pointer;
		write_pointer_n = write_pointer;
		status_cnt_n = status_cnt;
	end
	always @(*) begin : output_assignments
		if (empty)
			lsu_ctrl_o = lsu_req_i;
		else
			lsu_ctrl_o = mem_q[read_pointer_q * 152+:152];
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			mem_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			read_pointer_q <= 1'sb0;
		end
		else begin
			mem_q <= mem_n;
			status_cnt_q <= status_cnt_n;
			write_pointer_q <= write_pointer_n;
			read_pointer_q <= read_pointer_n;
		end
endmodule
module load_unit (
	clk_i,
	rst_ni,
	flush_i,
	valid_i,
	lsu_ctrl_i,
	pop_ld_o,
	valid_o,
	trans_id_o,
	result_o,
	ex_o,
	translation_req_o,
	vaddr_o,
	paddr_i,
	ex_i,
	dtlb_hit_i,
	dtlb_ppn_i,
	page_offset_o,
	page_offset_matches_i,
	store_buffer_empty_i,
	commit_tran_id_i,
	req_port_i,
	req_port_o,
	dcache_wbuffer_not_ni_i
);
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire valid_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [151:0] lsu_ctrl_i;
	output reg pop_ld_o;
	output reg valid_o;
	output reg [2:0] trans_id_o;
	output reg [63:0] result_o;
	output reg [128:0] ex_o;
	output reg translation_req_o;
	output wire [63:0] vaddr_o;
	localparam riscv_PLEN = 56;
	input wire [55:0] paddr_i;
	input wire [128:0] ex_i;
	input wire dtlb_hit_i;
	localparam riscv_PPNW = 44;
	input wire [43:0] dtlb_ppn_i;
	output wire [11:0] page_offset_o;
	input wire page_offset_matches_i;
	input wire store_buffer_empty_i;
	input wire [2:0] commit_tran_id_i;
	input wire [65:0] req_port_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output reg [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_o;
	input wire dcache_wbuffer_not_ni_i;
	reg [3:0] state_d;
	reg [3:0] state_q;
	reg [12:0] load_data_d;
	reg [12:0] load_data_q;
	wire [12:0] in_data;
	assign page_offset_o = lsu_ctrl_i[98:87];
	assign vaddr_o = lsu_ctrl_i[150-:64];
	wire [1:1] sv2v_tmp_3B099;
	assign sv2v_tmp_3B099 = 1'b0;
	always @(*) req_port_o[12] = sv2v_tmp_3B099;
	wire [64:1] sv2v_tmp_43C6F;
	assign sv2v_tmp_43C6F = 1'sb0;
	always @(*) req_port_o[77-:64] = sv2v_tmp_43C6F;
	assign in_data = {lsu_ctrl_i[2-:ariane_pkg_TRANS_ID_BITS], lsu_ctrl_i[89:87], lsu_ctrl_i[9-:7]};
	wire [12:1] sv2v_tmp_BD91C;
	assign sv2v_tmp_BD91C = lsu_ctrl_i[98:87];
	always @(*) req_port_o[133-:12] = sv2v_tmp_BD91C;
	wire [44:1] sv2v_tmp_49A7B;
	assign sv2v_tmp_49A7B = paddr_i[(ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_INDEX_WIDTH) - 1:ariane_pkg_DCACHE_INDEX_WIDTH];
	always @(*) req_port_o[121-:44] = sv2v_tmp_49A7B;
	wire [64:1] sv2v_tmp_C5B66;
	assign sv2v_tmp_C5B66 = ex_i[128-:64];
	always @(*) ex_o[128-:64] = sv2v_tmp_C5B66;
	wire [64:1] sv2v_tmp_39B40;
	assign sv2v_tmp_39B40 = ex_i[64-:64];
	always @(*) ex_o[64-:64] = sv2v_tmp_39B40;
	wire paddr_ni;
	wire not_commit_time;
	wire inflight_stores;
	wire stall_ni;
	function automatic ariane_pkg_range_check;
		input reg [63:0] base;
		input reg [63:0] len;
		input reg [63:0] address;
		ariane_pkg_range_check = (address >= base) && (address < (base + len));
	endfunction
	function automatic ariane_pkg_is_inside_nonidempotent_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_1
				reg [31:0] k;
				for (k = 0; k < Cfg[6337-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[5282 + (k * 64)+:64], Cfg[4258 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_nonidempotent_regions = |pass;
		end
	endfunction
	assign paddr_ni = ariane_pkg_is_inside_nonidempotent_regions(ArianeCfg, {dtlb_ppn_i, 12'd0});
	assign not_commit_time = commit_tran_id_i != lsu_ctrl_i[2-:ariane_pkg_TRANS_ID_BITS];
	assign inflight_stores = !dcache_wbuffer_not_ni_i || !store_buffer_empty_i;
	assign stall_ni = (inflight_stores || not_commit_time) && paddr_ni;
	function automatic [1:0] ariane_pkg_extract_transfer_size;
		input reg [6:0] op;
		case (op)
			7'd35, 7'd36, 7'd81, 7'd85, 7'd47, 7'd49, 7'd59, 7'd60, 7'd61, 7'd62, 7'd63, 7'd64, 7'd65, 7'd66, 7'd67: ariane_pkg_extract_transfer_size = 2'b11;
			7'd37, 7'd38, 7'd39, 7'd82, 7'd86, 7'd46, 7'd48, 7'd50, 7'd51, 7'd52, 7'd53, 7'd54, 7'd55, 7'd56, 7'd57, 7'd58: ariane_pkg_extract_transfer_size = 2'b10;
			7'd40, 7'd41, 7'd42, 7'd83, 7'd87: ariane_pkg_extract_transfer_size = 2'b01;
			7'd43, 7'd45, 7'd44, 7'd84, 7'd88: ariane_pkg_extract_transfer_size = 2'b00;
			default: ariane_pkg_extract_transfer_size = 2'b11;
		endcase
	endfunction
	always @(*) begin : load_control
		state_d = state_q;
		load_data_d = load_data_q;
		translation_req_o = 1'b0;
		req_port_o[13] = 1'b0;
		req_port_o[1] = 1'b0;
		req_port_o[0] = 1'b0;
		req_port_o[11-:8] = lsu_ctrl_i[21-:8];
		req_port_o[3-:2] = ariane_pkg_extract_transfer_size(lsu_ctrl_i[9-:7]);
		pop_ld_o = 1'b0;
		case (state_q)
			4'd0:
				if (valid_i) begin
					translation_req_o = 1'b1;
					if (!page_offset_matches_i) begin
						req_port_o[13] = 1'b1;
						if (!req_port_i[65])
							state_d = 4'd1;
						else if (dtlb_hit_i && !stall_ni) begin
							state_d = 4'd2;
							pop_ld_o = 1'b1;
						end
						else if (dtlb_hit_i && stall_ni)
							state_d = 4'd5;
						else
							state_d = 4'd4;
					end
					else
						state_d = 4'd3;
				end
			4'd3:
				if (!page_offset_matches_i)
					state_d = 4'd1;
			4'd4, 4'd5: begin
				req_port_o[1] = 1'b1;
				req_port_o[0] = 1'b1;
				state_d = (state_q == 4'd5 ? 4'd8 : 4'd6);
			end
			4'd8:
				if (dcache_wbuffer_not_ni_i)
					state_d = 4'd6;
			4'd6: begin
				translation_req_o = 1'b1;
				if (dtlb_hit_i)
					state_d = 4'd1;
			end
			4'd1: begin
				translation_req_o = 1'b1;
				req_port_o[13] = 1'b1;
				if (req_port_i[65]) begin
					if (dtlb_hit_i && !stall_ni) begin
						state_d = 4'd2;
						pop_ld_o = 1'b1;
					end
					else if (dtlb_hit_i && stall_ni)
						state_d = 4'd5;
					else
						state_d = 4'd4;
				end
			end
			4'd2: begin
				req_port_o[0] = 1'b1;
				state_d = 4'd0;
				if (valid_i) begin
					translation_req_o = 1'b1;
					if (!page_offset_matches_i) begin
						req_port_o[13] = 1'b1;
						if (!req_port_i[65])
							state_d = 4'd1;
						else if (dtlb_hit_i && !stall_ni) begin
							state_d = 4'd2;
							pop_ld_o = 1'b1;
						end
						else if (dtlb_hit_i && stall_ni)
							state_d = 4'd5;
						else
							state_d = 4'd4;
					end
					else
						state_d = 4'd3;
				end
				if (ex_i[0])
					req_port_o[1] = 1'b1;
			end
			4'd7: begin
				req_port_o[1] = 1'b1;
				req_port_o[0] = 1'b1;
				state_d = 4'd0;
			end
		endcase
		if (ex_i[0] && valid_i) begin
			state_d = 4'd0;
			if (!req_port_i[64])
				pop_ld_o = 1'b1;
		end
		if (pop_ld_o && !ex_i[0])
			load_data_d = in_data;
		if (flush_i)
			state_d = 4'd7;
	end
	always @(*) begin : rvalid_output
		valid_o = 1'b0;
		ex_o[0] = 1'b0;
		trans_id_o = load_data_q[12-:3];
		if (req_port_i[64] && (state_q != 4'd7)) begin
			if (!req_port_o[1])
				valid_o = 1'b1;
			if (ex_i[0] && (state_q == 4'd2)) begin
				valid_o = 1'b1;
				ex_o[0] = 1'b1;
			end
		end
		if ((valid_i && ex_i[0]) && !req_port_i[64]) begin
			valid_o = 1'b1;
			ex_o[0] = 1'b1;
			trans_id_o = lsu_ctrl_i[2-:ariane_pkg_TRANS_ID_BITS];
		end
		else if (state_q == 4'd6)
			valid_o = 1'b0;
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			state_q <= 4'd0;
			load_data_q <= 1'sb0;
		end
		else begin
			state_q <= state_d;
			load_data_q <= load_data_d;
		end
	wire [63:0] shifted_data;
	assign shifted_data = req_port_i[63-:64] >> {load_data_q[9-:3], 3'b000};
	wire [7:0] sign_bits;
	wire [2:0] idx_d;
	reg [2:0] idx_q;
	wire sign_bit;
	wire signed_d;
	reg signed_q;
	wire fp_sign_d;
	reg fp_sign_q;
	assign signed_d = |{load_data_d[6-:7] == 7'd37, load_data_d[6-:7] == 7'd40, load_data_d[6-:7] == 7'd43};
	assign fp_sign_d = |{load_data_d[6-:7] == 7'd82, load_data_d[6-:7] == 7'd83, load_data_d[6-:7] == 7'd84};
	assign idx_d = (|{load_data_d[6-:7] == 7'd37, load_data_d[6-:7] == 7'd82} ? load_data_d[9-:3] + 3 : (|{load_data_d[6-:7] == 7'd40, load_data_d[6-:7] == 7'd83} ? load_data_d[9-:3] + 1 : load_data_d[9-:3]));
	assign sign_bits = {req_port_i[63], req_port_i[55], req_port_i[47], req_port_i[39], req_port_i[31], req_port_i[23], req_port_i[15], req_port_i[7]};
	assign sign_bit = (signed_q & sign_bits[idx_q]) | fp_sign_q;
	always @(*)
		case (load_data_q[6-:7])
			7'd37, 7'd38, 7'd82: result_o = {{32 {sign_bit}}, shifted_data[31:0]};
			7'd40, 7'd41, 7'd83: result_o = {{48 {sign_bit}}, shifted_data[15:0]};
			7'd43, 7'd45, 7'd84: result_o = {{56 {sign_bit}}, shifted_data[7:0]};
			default: result_o = shifted_data[63:0];
		endcase
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (~rst_ni) begin
			idx_q <= 0;
			signed_q <= 0;
			fp_sign_q <= 0;
		end
		else begin
			idx_q <= idx_d;
			signed_q <= signed_d;
			fp_sign_q <= fp_sign_d;
		end
	end
endmodule
module mmu (
	clk_i,
	rst_ni,
	flush_i,
	enable_translation_i,
	en_ld_st_translation_i,
	icache_areq_i,
	icache_areq_o,
	misaligned_ex_i,
	lsu_req_i,
	lsu_vaddr_i,
	lsu_is_store_i,
	lsu_dtlb_hit_o,
	lsu_dtlb_ppn_o,
	lsu_valid_o,
	lsu_paddr_o,
	lsu_exception_o,
	priv_lvl_i,
	ld_st_priv_lvl_i,
	sum_i,
	mxr_i,
	satp_ppn_i,
	asid_i,
	asid_to_be_flushed_i,
	vaddr_to_be_flushed_i,
	flush_tlb_i,
	itlb_miss_o,
	dtlb_miss_o,
	req_port_i,
	req_port_o,
	pmpcfg_i,
	pmpaddr_i
);
	parameter [31:0] INSTR_TLB_ENTRIES = 4;
	parameter [31:0] DATA_TLB_ENTRIES = 4;
	parameter [31:0] ASID_WIDTH = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire enable_translation_i;
	input wire en_ld_st_translation_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [64:0] icache_areq_i;
	localparam riscv_PLEN = 56;
	output reg [185:0] icache_areq_o;
	input wire [128:0] misaligned_ex_i;
	input wire lsu_req_i;
	input wire [63:0] lsu_vaddr_i;
	input wire lsu_is_store_i;
	output wire lsu_dtlb_hit_o;
	localparam riscv_PPNW = 44;
	output reg [43:0] lsu_dtlb_ppn_o;
	output reg lsu_valid_o;
	output reg [55:0] lsu_paddr_o;
	output reg [128:0] lsu_exception_o;
	input wire [1:0] priv_lvl_i;
	input wire [1:0] ld_st_priv_lvl_i;
	input wire sum_i;
	input wire mxr_i;
	input wire [43:0] satp_ppn_i;
	input wire [ASID_WIDTH - 1:0] asid_i;
	input wire [ASID_WIDTH - 1:0] asid_to_be_flushed_i;
	input wire [63:0] vaddr_to_be_flushed_i;
	input wire flush_tlb_i;
	output wire itlb_miss_o;
	output wire dtlb_miss_o;
	input wire [65:0] req_port_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output wire [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_o;
	input wire [127:0] pmpcfg_i;
	input wire [863:0] pmpaddr_i;
	reg iaccess_err;
	reg daccess_err;
	wire ptw_active;
	wire walking_instr;
	wire ptw_error;
	wire ptw_access_exception;
	wire [55:0] ptw_bad_paddr;
	wire [63:0] update_vaddr;
	localparam ariane_pkg_ASID_WIDTH = 16;
	wire [109:0] update_ptw_itlb;
	wire [109:0] update_ptw_dtlb;
	wire itlb_lu_access;
	wire [63:0] itlb_content;
	wire itlb_is_2M;
	wire itlb_is_1G;
	wire itlb_lu_hit;
	wire dtlb_lu_access;
	wire [63:0] dtlb_content;
	wire dtlb_is_2M;
	wire dtlb_is_1G;
	wire dtlb_lu_hit;
	assign itlb_lu_access = icache_areq_i[64];
	assign dtlb_lu_access = lsu_req_i;
	tlb #(
		.TLB_ENTRIES(INSTR_TLB_ENTRIES),
		.ASID_WIDTH(ASID_WIDTH)
	) i_itlb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_tlb_i),
		.update_i(update_ptw_itlb),
		.lu_access_i(itlb_lu_access),
		.lu_asid_i(asid_i),
		.asid_to_be_flushed_i(asid_to_be_flushed_i),
		.vaddr_to_be_flushed_i(vaddr_to_be_flushed_i),
		.lu_vaddr_i(icache_areq_i[63-:riscv_VLEN]),
		.lu_content_o(itlb_content),
		.lu_is_2M_o(itlb_is_2M),
		.lu_is_1G_o(itlb_is_1G),
		.lu_hit_o(itlb_lu_hit)
	);
	tlb #(
		.TLB_ENTRIES(DATA_TLB_ENTRIES),
		.ASID_WIDTH(ASID_WIDTH)
	) i_dtlb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_tlb_i),
		.update_i(update_ptw_dtlb),
		.lu_access_i(dtlb_lu_access),
		.lu_asid_i(asid_i),
		.asid_to_be_flushed_i(asid_to_be_flushed_i),
		.vaddr_to_be_flushed_i(vaddr_to_be_flushed_i),
		.lu_vaddr_i(lsu_vaddr_i),
		.lu_content_o(dtlb_content),
		.lu_is_2M_o(dtlb_is_2M),
		.lu_is_1G_o(dtlb_is_1G),
		.lu_hit_o(dtlb_lu_hit)
	);
	ptw #(
		.ASID_WIDTH(ASID_WIDTH),
		.ArianeCfg(ArianeCfg)
	) i_ptw(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.ptw_active_o(ptw_active),
		.walking_instr_o(walking_instr),
		.ptw_error_o(ptw_error),
		.ptw_access_exception_o(ptw_access_exception),
		.enable_translation_i(enable_translation_i),
		.update_vaddr_o(update_vaddr),
		.itlb_update_o(update_ptw_itlb),
		.dtlb_update_o(update_ptw_dtlb),
		.itlb_access_i(itlb_lu_access),
		.itlb_hit_i(itlb_lu_hit),
		.itlb_vaddr_i(icache_areq_i[63-:riscv_VLEN]),
		.dtlb_access_i(dtlb_lu_access),
		.dtlb_hit_i(dtlb_lu_hit),
		.dtlb_vaddr_i(lsu_vaddr_i),
		.req_port_i(req_port_i),
		.req_port_o(req_port_o),
		.pmpcfg_i(pmpcfg_i),
		.pmpaddr_i(pmpaddr_i),
		.bad_paddr_o(ptw_bad_paddr),
		.flush_i(flush_i),
		.en_ld_st_translation_i(en_ld_st_translation_i),
		.lsu_is_store_i(lsu_is_store_i),
		.asid_i(asid_i),
		.satp_ppn_i(satp_ppn_i),
		.mxr_i(mxr_i),
		.itlb_miss_o(itlb_miss_o),
		.dtlb_miss_o(dtlb_miss_o)
	);
	wire match_any_execute_region;
	wire pmp_instr_allow;
	localparam [63:0] riscv_INSTR_ACCESS_FAULT = 1;
	localparam [63:0] riscv_INSTR_PAGE_FAULT = 12;
	localparam [3:0] riscv_MODE_SV = 4'd8;
	localparam riscv_SV = 39;
	always @(*) begin : instr_interface
		icache_areq_o[185] = icache_areq_i[64];
		icache_areq_o[184-:56] = icache_areq_i[55:0];
		icache_areq_o[128-:129] = 1'sb0;
		iaccess_err = icache_areq_i[64] && (((priv_lvl_i == 2'b00) && ~itlb_content[4]) || ((priv_lvl_i == 2'b01) && itlb_content[4]));
		if (enable_translation_i) begin
			if (icache_areq_i[64] && !((&icache_areq_i[63:38] == 1'b1) || (|icache_areq_i[63:38] == 1'b0)))
				icache_areq_o[128-:129] = {riscv_INSTR_ACCESS_FAULT, icache_areq_i[63-:riscv_VLEN], 1'b1};
			icache_areq_o[185] = 1'b0;
			icache_areq_o[184-:56] = {itlb_content[53-:44], icache_areq_i[11:0]};
			if (itlb_is_2M)
				icache_areq_o[149:141] = icache_areq_i[20:12];
			if (itlb_is_1G)
				icache_areq_o[158:141] = icache_areq_i[29:12];
			if (itlb_lu_hit) begin
				icache_areq_o[185] = icache_areq_i[64];
				if (iaccess_err)
					icache_areq_o[128-:129] = {riscv_INSTR_PAGE_FAULT, icache_areq_i[63-:riscv_VLEN], 1'b1};
				else if (!pmp_instr_allow)
					icache_areq_o[128-:129] = {riscv_INSTR_ACCESS_FAULT, {8 {1'b0}}, icache_areq_i[63-:riscv_VLEN], 1'b1};
			end
			else if (ptw_active && walking_instr) begin
				icache_areq_o[185] = ptw_error | ptw_access_exception;
				if (ptw_error)
					icache_areq_o[128-:129] = {riscv_INSTR_PAGE_FAULT, update_vaddr, 1'b1};
				else
					icache_areq_o[128-:129] = {riscv_INSTR_ACCESS_FAULT, ptw_bad_paddr, 1'b1};
			end
		end
		if (!match_any_execute_region || (!enable_translation_i && !pmp_instr_allow))
			icache_areq_o[128-:129] = {riscv_INSTR_ACCESS_FAULT, {8 {1'b0}}, icache_areq_o[184-:56], 1'b1};
	end
	function automatic ariane_pkg_range_check;
		input reg [63:0] base;
		input reg [63:0] len;
		input reg [63:0] address;
		ariane_pkg_range_check = (address >= base) && (address < (base + len));
	endfunction
	function automatic ariane_pkg_is_inside_execute_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_1
				reg [31:0] k;
				for (k = 0; k < Cfg[4257-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[3202 + (k * 64)+:64], Cfg[2178 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_execute_regions = |pass;
		end
	endfunction
	assign match_any_execute_region = ariane_pkg_is_inside_execute_regions(ArianeCfg, {{8 {1'b0}}, icache_areq_o[184-:56]});
	pmp #(
		.PLEN(riscv_PLEN),
		.PMP_LEN(54),
		.NR_ENTRIES(ArianeCfg[31-:32])
	) i_pmp_if(
		.addr_i(icache_areq_o[184-:56]),
		.priv_lvl_i(priv_lvl_i),
		.access_type_i(3'b100),
		.conf_addr_i(pmpaddr_i),
		.conf_i(pmpcfg_i),
		.allow_o(pmp_instr_allow)
	);
	reg [63:0] lsu_vaddr_n;
	reg [63:0] lsu_vaddr_q;
	reg [63:0] dtlb_pte_n;
	reg [63:0] dtlb_pte_q;
	reg [128:0] misaligned_ex_n;
	reg [128:0] misaligned_ex_q;
	reg lsu_req_n;
	reg lsu_req_q;
	reg lsu_is_store_n;
	reg lsu_is_store_q;
	reg dtlb_hit_n;
	reg dtlb_hit_q;
	reg dtlb_is_2M_n;
	reg dtlb_is_2M_q;
	reg dtlb_is_1G_n;
	reg dtlb_is_1G_q;
	assign lsu_dtlb_hit_o = (en_ld_st_translation_i ? dtlb_lu_hit : 1'b1);
	reg [2:0] pmp_access_type;
	wire pmp_data_allow;
	localparam PPNWMin = 29;
	localparam [63:0] riscv_LD_ACCESS_FAULT = 5;
	localparam [63:0] riscv_LOAD_PAGE_FAULT = 13;
	localparam [63:0] riscv_STORE_PAGE_FAULT = 15;
	localparam [63:0] riscv_ST_ACCESS_FAULT = 7;
	always @(*) begin : data_interface
		lsu_vaddr_n = lsu_vaddr_i;
		lsu_req_n = lsu_req_i;
		misaligned_ex_n = misaligned_ex_i;
		dtlb_pte_n = dtlb_content;
		dtlb_hit_n = dtlb_lu_hit;
		lsu_is_store_n = lsu_is_store_i;
		dtlb_is_2M_n = dtlb_is_2M;
		dtlb_is_1G_n = dtlb_is_1G;
		lsu_paddr_o = lsu_vaddr_q[55:0];
		lsu_dtlb_ppn_o = lsu_vaddr_n[55:12];
		lsu_valid_o = lsu_req_q;
		lsu_exception_o = misaligned_ex_q;
		pmp_access_type = (lsu_is_store_q ? 3'b010 : 3'b001);
		misaligned_ex_n[0] = misaligned_ex_i[0] & lsu_req_i;
		daccess_err = (((ld_st_priv_lvl_i == 2'b01) && !sum_i) && dtlb_pte_q[4]) || ((ld_st_priv_lvl_i == 2'b00) && !dtlb_pte_q[4]);
		if (en_ld_st_translation_i && !misaligned_ex_q[0]) begin
			lsu_valid_o = 1'b0;
			lsu_paddr_o = {dtlb_pte_q[53-:44], lsu_vaddr_q[11:0]};
			lsu_dtlb_ppn_o = dtlb_content[53-:44];
			if (dtlb_is_2M_q) begin
				lsu_paddr_o[20:12] = lsu_vaddr_q[20:12];
				lsu_dtlb_ppn_o[20:12] = lsu_vaddr_n[20:12];
			end
			if (dtlb_is_1G_q) begin
				lsu_paddr_o[PPNWMin:12] = lsu_vaddr_q[PPNWMin:12];
				lsu_dtlb_ppn_o[PPNWMin:12] = lsu_vaddr_n[PPNWMin:12];
			end
			if (dtlb_hit_q && lsu_req_q) begin
				lsu_valid_o = 1'b1;
				if (lsu_is_store_q) begin
					if ((!dtlb_pte_q[2] || daccess_err) || !dtlb_pte_q[7])
						lsu_exception_o = {riscv_STORE_PAGE_FAULT, lsu_vaddr_q, 1'b1};
					else if (!pmp_data_allow)
						lsu_exception_o = {riscv_ST_ACCESS_FAULT, {8 {1'b0}}, lsu_paddr_o, 1'b1};
				end
				else if (daccess_err)
					lsu_exception_o = {riscv_LOAD_PAGE_FAULT, lsu_vaddr_q, 1'b1};
				else if (!pmp_data_allow)
					lsu_exception_o = {riscv_LD_ACCESS_FAULT, {8 {1'b0}}, lsu_paddr_o, 1'b1};
			end
			else if (ptw_active && !walking_instr) begin
				if (ptw_error) begin
					lsu_valid_o = 1'b1;
					if (lsu_is_store_q)
						lsu_exception_o = {riscv_STORE_PAGE_FAULT, update_vaddr, 1'b1};
					else
						lsu_exception_o = {riscv_LOAD_PAGE_FAULT, update_vaddr, 1'b1};
				end
				if (ptw_access_exception) begin
					lsu_valid_o = 1'b1;
					lsu_exception_o = {riscv_LD_ACCESS_FAULT, {8 {1'b0}}, ptw_bad_paddr, 1'b1};
				end
			end
		end
		else if ((lsu_req_q && !misaligned_ex_q[0]) && !pmp_data_allow) begin
			if (lsu_is_store_q)
				lsu_exception_o = {riscv_ST_ACCESS_FAULT, {8 {1'b0}}, lsu_paddr_o, 1'b1};
			else
				lsu_exception_o = {riscv_LD_ACCESS_FAULT, {8 {1'b0}}, lsu_paddr_o, 1'b1};
		end
	end
	pmp #(
		.PLEN(riscv_PLEN),
		.PMP_LEN(54),
		.NR_ENTRIES(ArianeCfg[31-:32])
	) i_pmp_data(
		.addr_i(lsu_paddr_o),
		.priv_lvl_i(ld_st_priv_lvl_i),
		.access_type_i(pmp_access_type),
		.conf_addr_i(pmpaddr_i),
		.conf_i(pmpcfg_i),
		.allow_o(pmp_data_allow)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			lsu_vaddr_q <= 1'sb0;
			lsu_req_q <= 1'sb0;
			misaligned_ex_q <= 1'sb0;
			dtlb_pte_q <= 1'sb0;
			dtlb_hit_q <= 1'sb0;
			lsu_is_store_q <= 1'sb0;
			dtlb_is_2M_q <= 1'sb0;
			dtlb_is_1G_q <= 1'sb0;
		end
		else begin
			lsu_vaddr_q <= lsu_vaddr_n;
			lsu_req_q <= lsu_req_n;
			misaligned_ex_q <= misaligned_ex_n;
			dtlb_pte_q <= dtlb_pte_n;
			dtlb_hit_q <= dtlb_hit_n;
			lsu_is_store_q <= lsu_is_store_n;
			dtlb_is_2M_q <= dtlb_is_2M_n;
			dtlb_is_1G_q <= dtlb_is_1G_n;
		end
endmodule
module multiplier (
	clk_i,
	rst_ni,
	trans_id_i,
	mult_valid_i,
	operator_i,
	operand_a_i,
	operand_b_i,
	result_o,
	mult_valid_o,
	mult_ready_o,
	mult_trans_id_o
);
	input wire clk_i;
	input wire rst_ni;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	input wire [2:0] trans_id_i;
	input wire mult_valid_i;
	input wire [6:0] operator_i;
	localparam riscv_XLEN = 64;
	input wire [63:0] operand_a_i;
	input wire [63:0] operand_b_i;
	output reg [63:0] result_o;
	output wire mult_valid_o;
	output wire mult_ready_o;
	output wire [2:0] mult_trans_id_o;
	reg [2:0] trans_id_q;
	reg mult_valid_q;
	wire [6:0] operator_d;
	reg [6:0] operator_q;
	wire [127:0] mult_result_d;
	reg [127:0] mult_result_q;
	reg sign_a;
	reg sign_b;
	wire mult_valid;
	assign mult_valid_o = mult_valid_q;
	assign mult_trans_id_o = trans_id_q;
	assign mult_ready_o = 1'b1;
	assign mult_valid = mult_valid_i && |{operator_i == 7'd68, operator_i == 7'd69, operator_i == 7'd70, operator_i == 7'd71, operator_i == 7'd72};
	wire [127:0] mult_result;
	assign mult_result = $signed({operand_a_i[63] & sign_a, operand_a_i}) * $signed({operand_b_i[63] & sign_b, operand_b_i});
	always @(*) begin
		sign_a = 1'b0;
		sign_b = 1'b0;
		if (operator_i == 7'd69) begin
			sign_a = 1'b1;
			sign_b = 1'b1;
		end
		else if (operator_i == 7'd71)
			sign_a = 1'b1;
		else begin
			sign_a = 1'b0;
			sign_b = 1'b0;
		end
	end
	assign mult_result_d = $signed({operand_a_i[63] & sign_a, operand_a_i}) * $signed({operand_b_i[63] & sign_b, operand_b_i});
	assign operator_d = operator_i;
	function automatic [63:0] ariane_pkg_sext32;
		input reg [31:0] operand;
		ariane_pkg_sext32 = {{32 {operand[31]}}, operand[31:0]};
	endfunction
	always @(*) begin : p_selmux
		case (operator_q)
			7'd69, 7'd70, 7'd71: result_o = mult_result_q[127:riscv_XLEN];
			7'd72: result_o = ariane_pkg_sext32(mult_result_q[31:0]);
			default: result_o = mult_result_q[63:0];
		endcase
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			mult_valid_q <= 1'sb0;
			trans_id_q <= 1'sb0;
			operator_q <= 7'd68;
			mult_result_q <= 1'sb0;
		end
		else begin
			trans_id_q <= trans_id_i;
			mult_valid_q <= mult_valid;
			operator_q <= operator_d;
			mult_result_q <= mult_result_d;
		end
endmodule
module mult (
	clk_i,
	rst_ni,
	flush_i,
	fu_data_i,
	mult_valid_i,
	result_o,
	mult_valid_o,
	mult_ready_o,
	mult_trans_id_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	input wire [205:0] fu_data_i;
	input wire mult_valid_i;
	output wire [63:0] result_o;
	output wire mult_valid_o;
	output wire mult_ready_o;
	output wire [2:0] mult_trans_id_o;
	wire mul_valid;
	wire div_valid;
	wire div_ready_i;
	wire [2:0] mul_trans_id;
	wire [2:0] div_trans_id;
	wire [63:0] mul_result;
	wire [63:0] div_result;
	wire div_valid_op;
	wire mul_valid_op;
	assign mul_valid_op = (~flush_i && mult_valid_i) && |{fu_data_i[201-:7] == 7'd68, fu_data_i[201-:7] == 7'd69, fu_data_i[201-:7] == 7'd70, fu_data_i[201-:7] == 7'd71, fu_data_i[201-:7] == 7'd72};
	assign div_valid_op = (~flush_i && mult_valid_i) && |{fu_data_i[201-:7] == 7'd73, fu_data_i[201-:7] == 7'd74, fu_data_i[201-:7] == 7'd75, fu_data_i[201-:7] == 7'd76, fu_data_i[201-:7] == 7'd77, fu_data_i[201-:7] == 7'd78, fu_data_i[201-:7] == 7'd79, fu_data_i[201-:7] == 7'd80};
	assign div_ready_i = (mul_valid ? 1'b0 : 1'b1);
	assign mult_trans_id_o = (mul_valid ? mul_trans_id : div_trans_id);
	assign result_o = (mul_valid ? mul_result : div_result);
	assign mult_valid_o = div_valid | mul_valid;
	multiplier i_multiplier(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.trans_id_i(fu_data_i[2-:ariane_pkg_TRANS_ID_BITS]),
		.operator_i(fu_data_i[201-:7]),
		.operand_a_i(fu_data_i[194-:64]),
		.operand_b_i(fu_data_i[130-:64]),
		.result_o(mul_result),
		.mult_valid_i(mul_valid_op),
		.mult_valid_o(mul_valid),
		.mult_trans_id_o(mul_trans_id),
		.mult_ready_o()
	);
	reg [63:0] operand_b;
	reg [63:0] operand_a;
	wire [63:0] result;
	wire div_signed;
	wire rem;
	reg word_op_d;
	reg word_op_q;
	assign div_signed = |{fu_data_i[201-:7] == 7'd73, fu_data_i[201-:7] == 7'd75, fu_data_i[201-:7] == 7'd77, fu_data_i[201-:7] == 7'd79};
	assign rem = |{fu_data_i[201-:7] == 7'd77, fu_data_i[201-:7] == 7'd78, fu_data_i[201-:7] == 7'd79, fu_data_i[201-:7] == 7'd80};
	function automatic [63:0] ariane_pkg_sext32;
		input reg [31:0] operand;
		ariane_pkg_sext32 = {{32 {operand[31]}}, operand[31:0]};
	endfunction
	always @(*) begin
		operand_a = 1'sb0;
		operand_b = 1'sb0;
		word_op_d = word_op_q;
		if (mult_valid_i && |{fu_data_i[201-:7] == 7'd73, fu_data_i[201-:7] == 7'd74, fu_data_i[201-:7] == 7'd75, fu_data_i[201-:7] == 7'd76, fu_data_i[201-:7] == 7'd77, fu_data_i[201-:7] == 7'd78, fu_data_i[201-:7] == 7'd79, fu_data_i[201-:7] == 7'd80}) begin
			if (|{fu_data_i[201-:7] == 7'd75, fu_data_i[201-:7] == 7'd76, fu_data_i[201-:7] == 7'd79, fu_data_i[201-:7] == 7'd80}) begin
				if (div_signed) begin
					operand_a = ariane_pkg_sext32(fu_data_i[162:131]);
					operand_b = ariane_pkg_sext32(fu_data_i[98:67]);
				end
				else begin
					operand_a = fu_data_i[162:131];
					operand_b = fu_data_i[98:67];
				end
				word_op_d = 1'b1;
			end
			else begin
				operand_a = fu_data_i[194-:64];
				operand_b = fu_data_i[130-:64];
				word_op_d = 1'b0;
			end
		end
	end
	serdiv #(.WIDTH(riscv_XLEN)) i_div(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.id_i(fu_data_i[2-:ariane_pkg_TRANS_ID_BITS]),
		.op_a_i(operand_a),
		.op_b_i(operand_b),
		.opcode_i({rem, div_signed}),
		.in_vld_i(div_valid_op),
		.in_rdy_o(mult_ready_o),
		.flush_i(flush_i),
		.out_vld_o(div_valid),
		.out_rdy_i(div_ready_i),
		.id_o(div_trans_id),
		.res_o(result)
	);
	assign div_result = (word_op_q ? ariane_pkg_sext32(result) : result);
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			word_op_q <= 1'sb0;
		else
			word_op_q <= word_op_d;
endmodule
module perf_counters (
	clk_i,
	rst_ni,
	debug_mode_i,
	addr_i,
	we_i,
	data_i,
	data_o,
	commit_instr_i,
	commit_ack_i,
	l1_icache_miss_i,
	l1_dcache_miss_i,
	itlb_miss_i,
	dtlb_miss_i,
	sb_full_i,
	if_empty_i,
	ex_i,
	eret_i,
	resolved_branch_i
);
	input wire clk_i;
	input wire rst_ni;
	input wire debug_mode_i;
	input wire [4:0] addr_i;
	input wire we_i;
	localparam riscv_XLEN = 64;
	input wire [63:0] data_i;
	output reg [63:0] data_o;
	localparam ariane_pkg_NR_COMMIT_PORTS = 2;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_VLEN = 64;
	input wire [721:0] commit_instr_i;
	input wire [1:0] commit_ack_i;
	input wire l1_icache_miss_i;
	input wire l1_dcache_miss_i;
	input wire itlb_miss_i;
	input wire dtlb_miss_i;
	input wire sb_full_i;
	input wire if_empty_i;
	input wire [128:0] ex_i;
	input wire eret_i;
	input wire [133:0] resolved_branch_i;
	localparam [6:0] RegOffset = 12'hb03 >> 5;
	reg [(((12'hb10 - 12'hb03) + 1) * 64) + 180415:180416] perf_counter_d;
	reg [(((12'hb10 - 12'hb03) + 1) * 64) + 180415:180416] perf_counter_q;
	always @(*) begin : perf_counters
		perf_counter_d = perf_counter_q;
		data_o = 'b0;
		if (!debug_mode_i) begin
			if (l1_icache_miss_i)
				perf_counter_d[180416+:64] = perf_counter_q[180416+:64] + 1'b1;
			if (l1_dcache_miss_i)
				perf_counter_d[180480+:64] = perf_counter_q[180480+:64] + 1'b1;
			if (itlb_miss_i)
				perf_counter_d[180544+:64] = perf_counter_q[180544+:64] + 1'b1;
			if (dtlb_miss_i)
				perf_counter_d[180608+:64] = perf_counter_q[180608+:64] + 1'b1;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < 1; i = i + 1)
					if (commit_ack_i[i]) begin
						if (commit_instr_i[(i * 361) + 293-:4] == 4'd1)
							perf_counter_d[180672+:64] = perf_counter_q[180672+:64] + 1'b1;
						if (commit_instr_i[(i * 361) + 293-:4] == 4'd2)
							perf_counter_d[180736+:64] = perf_counter_q[180736+:64] + 1'b1;
						if (commit_instr_i[(i * 361) + 293-:4] == 4'd4)
							perf_counter_d[180928+:64] = perf_counter_q[180928+:64] + 1'b1;
						if (((commit_instr_i[(i * 361) + 293-:4] == 4'd4) && (commit_instr_i[(i * 361) + 289-:7] == {7 {1'sb0}})) && ((commit_instr_i[(i * 361) + 270-:6] == 'd1) || (commit_instr_i[(i * 361) + 270-:6] == 'd1)))
							perf_counter_d[180992+:64] = perf_counter_q[180992+:64] + 1'b1;
						if ((commit_instr_i[(i * 361) + 289-:7] == 7'd19) && ((commit_instr_i[(i * 361) + 270-:6] == 'd1) || (commit_instr_i[(i * 361) + 270-:6] == 'd1)))
							perf_counter_d[181056+:64] = perf_counter_q[181056+:64] + 1'b1;
					end
			end
			if (ex_i[0])
				perf_counter_d[180800+:64] = perf_counter_q[180800+:64] + 1'b1;
			if (eret_i)
				perf_counter_d[180864+:64] = perf_counter_q[180864+:64] + 1'b1;
			if (resolved_branch_i[133] && resolved_branch_i[4])
				perf_counter_d[181120+:64] = perf_counter_q[181120+:64] + 1'b1;
			if (sb_full_i)
				perf_counter_d[181184+:64] = perf_counter_q[181184+:64] + 1'b1;
			if (if_empty_i)
				perf_counter_d[181248+:64] = perf_counter_q[181248+:64] + 1'b1;
		end
		data_o = perf_counter_q[{RegOffset, addr_i} * 64+:64];
		if (we_i)
			perf_counter_d[{RegOffset, addr_i} * 64+:64] = data_i;
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			perf_counter_q <= 1'sb0;
		else
			perf_counter_q <= perf_counter_d;
endmodule
module ptw (
	clk_i,
	rst_ni,
	flush_i,
	ptw_active_o,
	walking_instr_o,
	ptw_error_o,
	ptw_access_exception_o,
	enable_translation_i,
	en_ld_st_translation_i,
	lsu_is_store_i,
	req_port_i,
	req_port_o,
	itlb_update_o,
	dtlb_update_o,
	update_vaddr_o,
	asid_i,
	itlb_access_i,
	itlb_hit_i,
	itlb_vaddr_i,
	dtlb_access_i,
	dtlb_hit_i,
	dtlb_vaddr_i,
	satp_ppn_i,
	mxr_i,
	itlb_miss_o,
	dtlb_miss_o,
	pmpcfg_i,
	pmpaddr_i,
	bad_paddr_o
);
	parameter signed [31:0] ASID_WIDTH = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	output wire ptw_active_o;
	output wire walking_instr_o;
	output reg ptw_error_o;
	output reg ptw_access_exception_o;
	input wire enable_translation_i;
	input wire en_ld_st_translation_i;
	input wire lsu_is_store_i;
	input wire [65:0] req_port_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output reg [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_o;
	localparam ariane_pkg_ASID_WIDTH = 16;
	output reg [109:0] itlb_update_o;
	output reg [109:0] dtlb_update_o;
	localparam riscv_VLEN = 64;
	output wire [63:0] update_vaddr_o;
	input wire [ASID_WIDTH - 1:0] asid_i;
	input wire itlb_access_i;
	input wire itlb_hit_i;
	input wire [63:0] itlb_vaddr_i;
	input wire dtlb_access_i;
	input wire dtlb_hit_i;
	input wire [63:0] dtlb_vaddr_i;
	localparam riscv_PPNW = 44;
	input wire [43:0] satp_ppn_i;
	input wire mxr_i;
	output reg itlb_miss_o;
	output reg dtlb_miss_o;
	input wire [127:0] pmpcfg_i;
	input wire [863:0] pmpaddr_i;
	output wire [55:0] bad_paddr_o;
	reg data_rvalid_q;
	reg [63:0] data_rdata_q;
	wire [63:0] pte;
	function automatic [63:0] sv2v_cast_DB804;
		input reg [63:0] inp;
		sv2v_cast_DB804 = inp;
	endfunction
	assign pte = sv2v_cast_DB804(data_rdata_q);
	reg [2:0] state_q;
	reg [2:0] state_d;
	reg [1:0] ptw_lvl_q;
	reg [1:0] ptw_lvl_n;
	reg is_instr_ptw_q;
	reg is_instr_ptw_n;
	reg global_mapping_q;
	reg global_mapping_n;
	reg tag_valid_n;
	reg tag_valid_q;
	reg kill_req_q;
	reg kill_req_d;
	reg [ASID_WIDTH - 1:0] tlb_update_asid_q;
	reg [ASID_WIDTH - 1:0] tlb_update_asid_n;
	reg [63:0] vaddr_q;
	reg [63:0] vaddr_n;
	reg [55:0] ptw_pptr_q;
	reg [55:0] ptw_pptr_n;
	assign update_vaddr_o = vaddr_q;
	assign ptw_active_o = state_q != 3'd0;
	assign walking_instr_o = is_instr_ptw_q;
	wire [12:1] sv2v_tmp_6E983;
	assign sv2v_tmp_6E983 = ptw_pptr_q[11:0];
	always @(*) req_port_o[133-:12] = sv2v_tmp_6E983;
	wire [44:1] sv2v_tmp_30D11;
	assign sv2v_tmp_30D11 = ptw_pptr_q[(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 1:ariane_pkg_DCACHE_INDEX_WIDTH];
	always @(*) req_port_o[121-:44] = sv2v_tmp_30D11;
	wire [1:1] sv2v_tmp_28F77;
	assign sv2v_tmp_28F77 = kill_req_q;
	always @(*) req_port_o[1] = sv2v_tmp_28F77;
	wire [64:1] sv2v_tmp_10C6E;
	assign sv2v_tmp_10C6E = 64'b0000000000000000000000000000000000000000000000000000000000000000;
	always @(*) req_port_o[77-:64] = sv2v_tmp_10C6E;
	localparam [3:0] riscv_MODE_SV = 4'd8;
	localparam riscv_SV = 39;
	wire [27:1] sv2v_tmp_66992;
	assign sv2v_tmp_66992 = {vaddr_q[38:12]};
	always @(*) itlb_update_o[106-:27] = sv2v_tmp_66992;
	wire [27:1] sv2v_tmp_549B3;
	assign sv2v_tmp_549B3 = {vaddr_q[38:12]};
	always @(*) dtlb_update_o[106-:27] = sv2v_tmp_549B3;
	wire [1:1] sv2v_tmp_378A1;
	assign sv2v_tmp_378A1 = ptw_lvl_q == 2'd1;
	always @(*) itlb_update_o[108] = sv2v_tmp_378A1;
	wire [1:1] sv2v_tmp_4A5B3;
	assign sv2v_tmp_4A5B3 = ptw_lvl_q == 2'd0;
	always @(*) itlb_update_o[107] = sv2v_tmp_4A5B3;
	wire [1:1] sv2v_tmp_79E68;
	assign sv2v_tmp_79E68 = ptw_lvl_q == 2'd1;
	always @(*) dtlb_update_o[108] = sv2v_tmp_79E68;
	wire [1:1] sv2v_tmp_F26AE;
	assign sv2v_tmp_F26AE = ptw_lvl_q == 2'd0;
	always @(*) dtlb_update_o[107] = sv2v_tmp_F26AE;
	wire [16:1] sv2v_tmp_61F34;
	assign sv2v_tmp_61F34 = tlb_update_asid_q;
	always @(*) itlb_update_o[79-:16] = sv2v_tmp_61F34;
	wire [16:1] sv2v_tmp_6FDCF;
	assign sv2v_tmp_6FDCF = tlb_update_asid_q;
	always @(*) dtlb_update_o[79-:16] = sv2v_tmp_6FDCF;
	wire [64:1] sv2v_tmp_EC01B;
	assign sv2v_tmp_EC01B = pte | (global_mapping_q << 5);
	always @(*) itlb_update_o[63-:64] = sv2v_tmp_EC01B;
	wire [64:1] sv2v_tmp_ECC9A;
	assign sv2v_tmp_ECC9A = pte | (global_mapping_q << 5);
	always @(*) dtlb_update_o[63-:64] = sv2v_tmp_ECC9A;
	wire [1:1] sv2v_tmp_7C039;
	assign sv2v_tmp_7C039 = tag_valid_q;
	always @(*) req_port_o[0] = sv2v_tmp_7C039;
	wire allow_access;
	assign bad_paddr_o = (ptw_access_exception_o ? ptw_pptr_q : 'b0);
	pmp #(
		.PLEN(riscv_PLEN),
		.PMP_LEN(54),
		.NR_ENTRIES(ArianeCfg[31-:32])
	) i_pmp_ptw(
		.addr_i(ptw_pptr_q),
		.priv_lvl_i(2'b01),
		.access_type_i(3'b001),
		.conf_addr_i(pmpaddr_i),
		.conf_i(pmpcfg_i),
		.allow_o(allow_access)
	);
	always @(*) begin : ptw
		tag_valid_n = 1'b0;
		kill_req_d = 1'b0;
		req_port_o[13] = 1'b0;
		req_port_o[11-:8] = 8'hff;
		req_port_o[3-:2] = 2'b11;
		req_port_o[12] = 1'b0;
		ptw_error_o = 1'b0;
		ptw_access_exception_o = 1'b0;
		itlb_update_o[109] = 1'b0;
		dtlb_update_o[109] = 1'b0;
		is_instr_ptw_n = is_instr_ptw_q;
		ptw_lvl_n = ptw_lvl_q;
		ptw_pptr_n = ptw_pptr_q;
		state_d = state_q;
		global_mapping_n = global_mapping_q;
		tlb_update_asid_n = tlb_update_asid_q;
		vaddr_n = vaddr_q;
		itlb_miss_o = 1'b0;
		dtlb_miss_o = 1'b0;
		case (state_q)
			3'd0: begin
				ptw_lvl_n = 2'd0;
				global_mapping_n = 1'b0;
				is_instr_ptw_n = 1'b0;
				if (((enable_translation_i & itlb_access_i) & ~itlb_hit_i) & ~dtlb_access_i) begin
					ptw_pptr_n = {satp_ppn_i, itlb_vaddr_i[38:30], 3'b000};
					is_instr_ptw_n = 1'b1;
					tlb_update_asid_n = asid_i;
					vaddr_n = itlb_vaddr_i;
					state_d = 3'd1;
					itlb_miss_o = 1'b1;
				end
				else if ((en_ld_st_translation_i & dtlb_access_i) & ~dtlb_hit_i) begin
					ptw_pptr_n = {satp_ppn_i, dtlb_vaddr_i[38:30], 3'b000};
					tlb_update_asid_n = asid_i;
					vaddr_n = dtlb_vaddr_i;
					state_d = 3'd1;
					dtlb_miss_o = 1'b1;
				end
			end
			3'd1: begin
				req_port_o[13] = 1'b1;
				if (req_port_i[65]) begin
					tag_valid_n = 1'b1;
					state_d = 3'd2;
				end
			end
			3'd2:
				if (data_rvalid_q) begin
					if (pte[5])
						global_mapping_n = 1'b1;
					if (!pte[0] || (!pte[1] && pte[2]))
						state_d = 3'd3;
					else begin
						state_d = 3'd0;
						if (pte[1] || pte[3]) begin
							if (is_instr_ptw_q) begin
								if (!pte[3] || !pte[6])
									state_d = 3'd3;
								else
									itlb_update_o[109] = 1'b1;
							end
							else begin
								if (pte[6] && (pte[1] || (pte[3] && mxr_i)))
									dtlb_update_o[109] = 1'b1;
								else
									state_d = 3'd3;
								if (lsu_is_store_i && (!pte[2] || !pte[7])) begin
									dtlb_update_o[109] = 1'b0;
									state_d = 3'd3;
								end
							end
							if ((ptw_lvl_q == 2'd0) && (pte[27:10] != {18 {1'sb0}})) begin
								state_d = 3'd3;
								dtlb_update_o[109] = 1'b0;
								itlb_update_o[109] = 1'b0;
							end
							else if ((ptw_lvl_q == 2'd1) && (pte[18:10] != {9 {1'sb0}})) begin
								state_d = 3'd3;
								dtlb_update_o[109] = 1'b0;
								itlb_update_o[109] = 1'b0;
							end
						end
						else begin
							if (ptw_lvl_q == 2'd0) begin
								ptw_lvl_n = 2'd1;
								ptw_pptr_n = {pte[53-:44], vaddr_q[29:21], 3'b000};
							end
							if (ptw_lvl_q == 2'd1) begin
								ptw_lvl_n = 2'd2;
								ptw_pptr_n = {pte[53-:44], vaddr_q[20:12], 3'b000};
							end
							state_d = 3'd1;
							if (ptw_lvl_q == 2'd2) begin
								ptw_lvl_n = 2'd2;
								state_d = 3'd3;
							end
						end
					end
					if (!allow_access) begin
						itlb_update_o[109] = 1'b0;
						dtlb_update_o[109] = 1'b0;
						ptw_pptr_n = ptw_pptr_q;
						state_d = 3'd4;
					end
				end
			3'd3: begin
				state_d = 3'd0;
				ptw_error_o = 1'b1;
			end
			3'd4: begin
				state_d = 3'd0;
				ptw_access_exception_o = 1'b1;
			end
			default: state_d = 3'd0;
		endcase
		if (flush_i) begin
			if (((state_q == 3'd2) && !data_rvalid_q) || ((state_q == 3'd1) && req_port_i[65])) begin
				tag_valid_n = 1'b1;
				kill_req_d = 1'b1;
			end
			state_d = 3'd0;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			state_q <= 3'd0;
			is_instr_ptw_q <= 1'b0;
			ptw_lvl_q <= 2'd0;
			tag_valid_q <= 1'b0;
			tlb_update_asid_q <= 1'sb0;
			vaddr_q <= 1'sb0;
			ptw_pptr_q <= 1'sb0;
			global_mapping_q <= 1'b0;
			data_rdata_q <= 1'sb0;
			data_rvalid_q <= 1'b0;
			kill_req_q <= 1'b0;
		end
		else begin
			state_q <= state_d;
			ptw_pptr_q <= ptw_pptr_n;
			is_instr_ptw_q <= is_instr_ptw_n;
			ptw_lvl_q <= ptw_lvl_n;
			tag_valid_q <= tag_valid_n;
			tlb_update_asid_q <= tlb_update_asid_n;
			vaddr_q <= vaddr_n;
			global_mapping_q <= global_mapping_n;
			data_rdata_q <= req_port_i[63-:64];
			data_rvalid_q <= req_port_i[64];
			kill_req_q <= kill_req_d;
		end
endmodule
module re_name (
	clk_i,
	rst_ni,
	flush_i,
	flush_unissied_instr_i,
	issue_instr_i,
	issue_instr_valid_i,
	issue_ack_o,
	issue_instr_o,
	issue_instr_valid_o,
	issue_ack_i
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire flush_unissied_instr_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [360:0] issue_instr_i;
	input wire issue_instr_valid_i;
	output wire issue_ack_o;
	output reg [360:0] issue_instr_o;
	output wire issue_instr_valid_o;
	input wire issue_ack_i;
	assign issue_instr_valid_o = issue_instr_valid_i;
	assign issue_ack_o = issue_ack_i;
	reg [31:0] re_name_table_gpr_n;
	reg [31:0] re_name_table_gpr_q;
	reg [31:0] re_name_table_fpr_n;
	reg [31:0] re_name_table_fpr_q;
	localparam ariane_pkg_ENABLE_RENAME = 1'b0;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	function automatic ariane_pkg_is_imm_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd89 <= op) && (7'd90 >= op), (7'd95 <= op) && (7'd98 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_imm_fpr = 1'b1;
			else
				ariane_pkg_is_imm_fpr = 1'b0;
		end
		else
			ariane_pkg_is_imm_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rd_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd81 <= op) && (7'd84 >= op), (7'd89 <= op) && (7'd98 >= op), op == 7'd100, op == 7'd101, op == 7'd102, op == 7'd104, (7'd107 <= op) && (7'd111 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rd_fpr = 1'b1;
			else
				ariane_pkg_is_rd_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rd_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs1_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd91 <= op) && (7'd98 >= op), op == 7'd99, op == 7'd101, op == 7'd102, op == 7'd103, op == 7'd105, op == 7'd106, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs1_fpr = 1'b1;
			else
				ariane_pkg_is_rs1_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs1_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs2_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd85 <= op) && (7'd88 >= op), (7'd89 <= op) && (7'd93 >= op), (7'd95 <= op) && (7'd98 >= op), op == 7'd101, (7'd102 <= op) && (7'd103 >= op), op == 7'd105, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs2_fpr = 1'b1;
			else
				ariane_pkg_is_rs2_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs2_fpr = 1'b0;
	endfunction
	always @(*) begin : sv2v_autoblock_1
		reg name_bit_rs1;
		reg name_bit_rs2;
		reg name_bit_rs3;
		reg name_bit_rd;
		re_name_table_gpr_n = re_name_table_gpr_q;
		re_name_table_fpr_n = re_name_table_fpr_q;
		issue_instr_o = issue_instr_i;
		if (issue_ack_i && !flush_unissied_instr_i) begin
			if (ariane_pkg_is_rd_fpr(issue_instr_i[289-:7]))
				re_name_table_fpr_n[issue_instr_i[270-:6]] = re_name_table_fpr_q[issue_instr_i[270-:6]] ^ 1'b1;
			else
				re_name_table_gpr_n[issue_instr_i[270-:6]] = re_name_table_gpr_q[issue_instr_i[270-:6]] ^ 1'b1;
		end
		name_bit_rs1 = (ariane_pkg_is_rs1_fpr(issue_instr_i[289-:7]) ? re_name_table_fpr_q[issue_instr_i[282-:6]] : re_name_table_gpr_q[issue_instr_i[282-:6]]);
		name_bit_rs2 = (ariane_pkg_is_rs2_fpr(issue_instr_i[289-:7]) ? re_name_table_fpr_q[issue_instr_i[276-:6]] : re_name_table_gpr_q[issue_instr_i[276-:6]]);
		name_bit_rs3 = re_name_table_fpr_q[issue_instr_i[205:201]];
		name_bit_rd = (ariane_pkg_is_rd_fpr(issue_instr_i[289-:7]) ? re_name_table_fpr_q[issue_instr_i[270-:6]] ^ 1'b1 : re_name_table_gpr_q[issue_instr_i[270-:6]] ^ (issue_instr_i[270-:6] != {6 {1'sb0}}));
		issue_instr_o[282-:6] = {ariane_pkg_ENABLE_RENAME & name_bit_rs1, issue_instr_i[281:277]};
		issue_instr_o[276-:6] = {ariane_pkg_ENABLE_RENAME & name_bit_rs2, issue_instr_i[275:271]};
		if (ariane_pkg_is_imm_fpr(issue_instr_i[289-:7]))
			issue_instr_o[264-:64] = {ariane_pkg_ENABLE_RENAME & name_bit_rs3, issue_instr_i[205:201]};
		issue_instr_o[270-:6] = {ariane_pkg_ENABLE_RENAME & name_bit_rd, issue_instr_i[269:265]};
		re_name_table_gpr_n[0] = 1'b0;
		if (flush_i) begin
			re_name_table_gpr_n = 1'sb0;
			re_name_table_fpr_n = 1'sb0;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			re_name_table_gpr_q <= 1'sb0;
			re_name_table_fpr_q <= 1'sb0;
		end
		else begin
			re_name_table_gpr_q <= re_name_table_gpr_n;
			re_name_table_fpr_q <= re_name_table_fpr_n;
		end
endmodule
module scoreboard (
	clk_i,
	rst_ni,
	sb_full_o,
	flush_unissued_instr_i,
	flush_i,
	unresolved_branch_i,
	rd_clobber_gpr_o,
	rd_clobber_fpr_o,
	rs1_i,
	rs1_o,
	rs1_valid_o,
	rs2_i,
	rs2_o,
	rs2_valid_o,
	rs3_i,
	rs3_o,
	rs3_valid_o,
	commit_instr_o,
	commit_ack_i,
	decoded_instr_i,
	decoded_instr_valid_i,
	decoded_instr_ack_o,
	issue_instr_o,
	issue_instr_valid_o,
	issue_ack_i,
	resolved_branch_i,
	trans_id_i,
	wbdata_i,
	ex_i,
	wt_valid_i
);
	parameter [31:0] NR_ENTRIES = 8;
	parameter [31:0] NR_WB_PORTS = 1;
	parameter [31:0] NR_COMMIT_PORTS = 2;
	input wire clk_i;
	input wire rst_ni;
	output wire sb_full_o;
	input wire flush_unissued_instr_i;
	input wire flush_i;
	input wire unresolved_branch_i;
	localparam ariane_pkg_REG_ADDR_SIZE = 6;
	output wire [255:0] rd_clobber_gpr_o;
	output wire [255:0] rd_clobber_fpr_o;
	input wire [5:0] rs1_i;
	localparam riscv_XLEN = 64;
	output wire [63:0] rs1_o;
	output wire rs1_valid_o;
	input wire [5:0] rs2_i;
	output wire [63:0] rs2_o;
	output wire rs2_valid_o;
	input wire [5:0] rs3_i;
	localparam riscv_IS_XLEN64 = 1'b1;
	localparam [0:0] ariane_pkg_RVD = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_RVF = riscv_IS_XLEN64;
	localparam [0:0] ariane_pkg_XF16 = 1'b0;
	localparam [0:0] ariane_pkg_XF16ALT = 1'b0;
	localparam [0:0] ariane_pkg_XF8 = 1'b0;
	localparam ariane_pkg_FLEN = (ariane_pkg_RVD ? 64 : (ariane_pkg_RVF ? 32 : (ariane_pkg_XF16 ? 16 : (ariane_pkg_XF16ALT ? 16 : (ariane_pkg_XF8 ? 8 : 1)))));
	output wire [ariane_pkg_FLEN - 1:0] rs3_o;
	output wire rs3_valid_o;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_VLEN = 64;
	output reg [(NR_COMMIT_PORTS * 361) - 1:0] commit_instr_o;
	input wire [NR_COMMIT_PORTS - 1:0] commit_ack_i;
	input wire [360:0] decoded_instr_i;
	input wire decoded_instr_valid_i;
	output reg decoded_instr_ack_o;
	output reg [360:0] issue_instr_o;
	output reg issue_instr_valid_o;
	input wire issue_ack_i;
	input wire [133:0] resolved_branch_i;
	input wire [(NR_WB_PORTS * 3) - 1:0] trans_id_i;
	input wire [(NR_WB_PORTS * 64) - 1:0] wbdata_i;
	input wire [(NR_WB_PORTS * 129) - 1:0] ex_i;
	input wire [NR_WB_PORTS - 1:0] wt_valid_i;
	localparam [31:0] BITS_ENTRIES = $clog2(NR_ENTRIES);
	reg [(NR_ENTRIES * 363) - 1:0] mem_q;
	reg [(NR_ENTRIES * 363) - 1:0] mem_n;
	wire issue_full;
	reg issue_en;
	wire [BITS_ENTRIES - 1:0] issue_cnt_n;
	reg [BITS_ENTRIES - 1:0] issue_cnt_q;
	wire [BITS_ENTRIES - 1:0] issue_pointer_n;
	reg [BITS_ENTRIES - 1:0] issue_pointer_q;
	wire [(NR_COMMIT_PORTS * BITS_ENTRIES) - 1:0] commit_pointer_n;
	reg [(NR_COMMIT_PORTS * BITS_ENTRIES) - 1:0] commit_pointer_q;
	wire [$clog2(NR_COMMIT_PORTS):0] num_commit;
	assign issue_full = &issue_cnt_q;
	assign sb_full_o = issue_full;
	always @(*) begin : commit_ports
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < NR_COMMIT_PORTS; i = i + 1)
				begin
					commit_instr_o[i * 361+:361] = mem_q[(commit_pointer_q[i * BITS_ENTRIES+:BITS_ENTRIES] * 363) + 360-:361];
					commit_instr_o[(i * 361) + 296-:3] = commit_pointer_q[i * BITS_ENTRIES+:BITS_ENTRIES];
				end
		end
	end
	always @(*) begin
		issue_instr_o = decoded_instr_i;
		issue_instr_o[296-:3] = issue_pointer_q;
		issue_instr_valid_o = (decoded_instr_valid_i & ~unresolved_branch_i) & ~issue_full;
		decoded_instr_ack_o = issue_ack_i & ~issue_full;
	end
	localparam [0:0] ariane_pkg_FP_PRESENT = (((ariane_pkg_RVF | ariane_pkg_RVD) | ariane_pkg_XF16) | ariane_pkg_XF16ALT) | ariane_pkg_XF8;
	function automatic ariane_pkg_is_rd_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd81 <= op) && (7'd84 >= op), (7'd89 <= op) && (7'd98 >= op), op == 7'd100, op == 7'd101, op == 7'd102, op == 7'd104, (7'd107 <= op) && (7'd111 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rd_fpr = 1'b1;
			else
				ariane_pkg_is_rd_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rd_fpr = 1'b0;
	endfunction
	always @(*) begin : issue_fifo
		mem_n = mem_q;
		issue_en = 1'b0;
		if ((decoded_instr_valid_i && decoded_instr_ack_o) && !flush_unissued_instr_i) begin
			issue_en = 1'b1;
			mem_n[issue_pointer_q * 363+:363] = {1'b1, ariane_pkg_is_rd_fpr(decoded_instr_i[289-:7]), decoded_instr_i};
		end
		begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < NR_ENTRIES; i = i + 1)
				if ((mem_q[(i * 363) + 293-:4] == 4'd0) && mem_q[(i * 363) + 362])
					mem_n[(i * 363) + 200] = 1'b1;
		end
		begin : sv2v_autoblock_3
			reg [31:0] i;
			for (i = 0; i < NR_WB_PORTS; i = i + 1)
				if (wt_valid_i[i] && mem_q[(trans_id_i[i * 3+:3] * 363) + 362]) begin
					mem_n[(trans_id_i[i * 3+:3] * 363) + 200] = 1'b1;
					mem_n[(trans_id_i[i * 3+:3] * 363) + 264-:64] = wbdata_i[i * 64+:64];
					mem_n[(trans_id_i[i * 3+:3] * 363) + 64-:riscv_VLEN] = resolved_branch_i[68-:64];
					if (ex_i[(i * 129) + 0])
						mem_n[(trans_id_i[i * 3+:3] * 363) + 196-:129] = ex_i[0 + (i * 129)+:129];
					else if (|{mem_q[(trans_id_i[i * 3+:3] * 363) + 293-:4] == 4'd7, mem_q[(trans_id_i[i * 3+:3] * 363) + 293-:4] == 4'd8})
						mem_n[(trans_id_i[i * 3+:3] * 363) + 196-:64] = ex_i[(i * 129) + 128-:64];
				end
		end
		begin : sv2v_autoblock_4
			reg [BITS_ENTRIES - 1:0] i;
			for (i = 0; i < NR_COMMIT_PORTS; i = i + 1)
				if (commit_ack_i[i]) begin
					mem_n[(commit_pointer_q[i * BITS_ENTRIES+:BITS_ENTRIES] * 363) + 362] = 1'b0;
					mem_n[(commit_pointer_q[i * BITS_ENTRIES+:BITS_ENTRIES] * 363) + 200] = 1'b0;
				end
		end
		if (flush_i) begin : sv2v_autoblock_5
			reg [31:0] i;
			for (i = 0; i < NR_ENTRIES; i = i + 1)
				begin
					mem_n[(i * 363) + 362] = 1'b0;
					mem_n[(i * 363) + 200] = 1'b0;
					mem_n[(i * 363) + 68] = 1'b0;
				end
		end
	end
	popcount #(.INPUT_WIDTH(NR_COMMIT_PORTS)) i_popcount(
		.data_i(commit_ack_i),
		.popcount_o(num_commit)
	);
	assign issue_cnt_n = (flush_i ? {BITS_ENTRIES {1'sb0}} : (issue_cnt_q - num_commit) + issue_en);
	assign commit_pointer_n[0+:BITS_ENTRIES] = (flush_i ? {BITS_ENTRIES * 1 {1'sb0}} : commit_pointer_q[0+:BITS_ENTRIES] + num_commit);
	assign issue_pointer_n = (flush_i ? {BITS_ENTRIES {1'sb0}} : issue_pointer_q + issue_en);
	genvar k;
	generate
		for (k = 1; k < NR_COMMIT_PORTS; k = k + 1) begin : gen_cnt_incr
			assign commit_pointer_n[k * BITS_ENTRIES+:BITS_ENTRIES] = (flush_i ? {BITS_ENTRIES * 1 {1'sb0}} : commit_pointer_n[0+:BITS_ENTRIES] + $unsigned(k));
		end
	endgenerate
	reg [(NR_ENTRIES >= 0 ? (64 * (NR_ENTRIES + 1)) - 1 : (64 * (1 - NR_ENTRIES)) + (NR_ENTRIES - 1)):(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES + 0)] gpr_clobber_vld;
	reg [(NR_ENTRIES >= 0 ? (64 * (NR_ENTRIES + 1)) - 1 : (64 * (1 - NR_ENTRIES)) + (NR_ENTRIES - 1)):(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES + 0)] fpr_clobber_vld;
	reg [(NR_ENTRIES >= 0 ? ((NR_ENTRIES + 1) * 4) - 1 : ((1 - NR_ENTRIES) * 4) + ((NR_ENTRIES * 4) - 1)):(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES * 4)] clobber_fu;
	always @(*) begin : clobber_assign
		gpr_clobber_vld = 1'sb0;
		fpr_clobber_vld = 1'sb0;
		clobber_fu[(NR_ENTRIES >= 0 ? NR_ENTRIES : NR_ENTRIES - NR_ENTRIES) * 4+:4] = 4'd0;
		begin : sv2v_autoblock_6
			reg [31:0] i;
			for (i = 0; i < 64; i = i + 1)
				begin
					gpr_clobber_vld[(i * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)) + (NR_ENTRIES >= 0 ? NR_ENTRIES : NR_ENTRIES - NR_ENTRIES)] = 1'b1;
					fpr_clobber_vld[(i * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)) + (NR_ENTRIES >= 0 ? NR_ENTRIES : NR_ENTRIES - NR_ENTRIES)] = 1'b1;
				end
		end
		begin : sv2v_autoblock_7
			reg [31:0] i;
			for (i = 0; i < NR_ENTRIES; i = i + 1)
				begin
					gpr_clobber_vld[(mem_q[(i * 363) + 270-:6] * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)) + (NR_ENTRIES >= 0 ? i : NR_ENTRIES - i)] = mem_q[(i * 363) + 362] & ~mem_q[(i * 363) + 361];
					fpr_clobber_vld[(mem_q[(i * 363) + 270-:6] * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)) + (NR_ENTRIES >= 0 ? i : NR_ENTRIES - i)] = mem_q[(i * 363) + 362] & mem_q[(i * 363) + 361];
					clobber_fu[(NR_ENTRIES >= 0 ? i : NR_ENTRIES - i) * 4+:4] = mem_q[(i * 363) + 293-:4];
				end
		end
		gpr_clobber_vld[(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES) + 0+:(NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)] = 1'sb0;
	end
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	generate
		for (k = 0; k < 64; k = k + 1) begin : gen_sel_clobbers
			localparam [31:0] sv2v_uu_i_sel_gpr_clobbers_NumIn = NR_ENTRIES + 1;
			localparam [$clog2(sv2v_cast_32(NR_ENTRIES + 1)) - 1:0] sv2v_uu_i_sel_gpr_clobbers_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_88014 #(
				.NumIn(NR_ENTRIES + 1),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_gpr_clobbers(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_gpr_clobbers_ext_rr_i_0),
				.req_i(gpr_clobber_vld[(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES) + (k * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES))+:(NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)]),
				.gnt_o(),
				.data_i(clobber_fu),
				.gnt_i(1'b1),
				.req_o(),
				.data_o(rd_clobber_gpr_o[k * 4+:4]),
				.idx_o()
			);
			localparam [31:0] sv2v_uu_i_sel_fpr_clobbers_NumIn = NR_ENTRIES + 1;
			localparam [$clog2(sv2v_cast_32(NR_ENTRIES + 1)) - 1:0] sv2v_uu_i_sel_fpr_clobbers_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_88014 #(
				.NumIn(NR_ENTRIES + 1),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1)
			) i_sel_fpr_clobbers(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.rr_i(sv2v_uu_i_sel_fpr_clobbers_ext_rr_i_0),
				.req_i(fpr_clobber_vld[(NR_ENTRIES >= 0 ? 0 : NR_ENTRIES) + (k * (NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES))+:(NR_ENTRIES >= 0 ? NR_ENTRIES + 1 : 1 - NR_ENTRIES)]),
				.gnt_o(),
				.data_i(clobber_fu),
				.gnt_i(1'b1),
				.req_o(),
				.data_o(rd_clobber_fpr_o[k * 4+:4]),
				.idx_o()
			);
		end
	endgenerate
	wire [(NR_ENTRIES + NR_WB_PORTS) - 1:0] rs1_fwd_req;
	wire [(NR_ENTRIES + NR_WB_PORTS) - 1:0] rs2_fwd_req;
	wire [(NR_ENTRIES + NR_WB_PORTS) - 1:0] rs3_fwd_req;
	wire [((NR_ENTRIES + NR_WB_PORTS) * 64) - 1:0] rs_data;
	wire rs1_valid;
	wire rs2_valid;
	function automatic ariane_pkg_is_imm_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd89 <= op) && (7'd90 >= op), (7'd95 <= op) && (7'd98 >= op), (7'd118 <= op) && (7'd121 >= op)})
				ariane_pkg_is_imm_fpr = 1'b1;
			else
				ariane_pkg_is_imm_fpr = 1'b0;
		end
		else
			ariane_pkg_is_imm_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs1_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd91 <= op) && (7'd98 >= op), op == 7'd99, op == 7'd101, op == 7'd102, op == 7'd103, op == 7'd105, op == 7'd106, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs1_fpr = 1'b1;
			else
				ariane_pkg_is_rs1_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs1_fpr = 1'b0;
	endfunction
	function automatic ariane_pkg_is_rs2_fpr;
		input reg [6:0] op;
		if (ariane_pkg_FP_PRESENT) begin
			if (|{(7'd85 <= op) && (7'd88 >= op), (7'd89 <= op) && (7'd93 >= op), (7'd95 <= op) && (7'd98 >= op), op == 7'd101, (7'd102 <= op) && (7'd103 >= op), op == 7'd105, (7'd107 <= op) && (7'd121 >= op)})
				ariane_pkg_is_rs2_fpr = 1'b1;
			else
				ariane_pkg_is_rs2_fpr = 1'b0;
		end
		else
			ariane_pkg_is_rs2_fpr = 1'b0;
	endfunction
	generate
		for (k = 0; $unsigned(k) < NR_WB_PORTS; k = k + 1) begin : gen_rs_wb
			assign rs1_fwd_req[k] = (((mem_q[(trans_id_i[k * 3+:3] * 363) + 270-:6] == rs1_i) & wt_valid_i[k]) & ~ex_i[(k * 129) + 0]) & (mem_q[(trans_id_i[k * 3+:3] * 363) + 361] == ariane_pkg_is_rs1_fpr(issue_instr_o[289-:7]));
			assign rs2_fwd_req[k] = (((mem_q[(trans_id_i[k * 3+:3] * 363) + 270-:6] == rs2_i) & wt_valid_i[k]) & ~ex_i[(k * 129) + 0]) & (mem_q[(trans_id_i[k * 3+:3] * 363) + 361] == ariane_pkg_is_rs2_fpr(issue_instr_o[289-:7]));
			assign rs3_fwd_req[k] = (((mem_q[(trans_id_i[k * 3+:3] * 363) + 270-:6] == rs3_i) & wt_valid_i[k]) & ~ex_i[(k * 129) + 0]) & (mem_q[(trans_id_i[k * 3+:3] * 363) + 361] == ariane_pkg_is_imm_fpr(issue_instr_o[289-:7]));
			assign rs_data[k * 64+:64] = wbdata_i[k * 64+:64];
		end
		for (k = 0; $unsigned(k) < NR_ENTRIES; k = k + 1) begin : gen_rs_entries
			assign rs1_fwd_req[k + NR_WB_PORTS] = (((mem_q[(k * 363) + 270-:6] == rs1_i) & mem_q[(k * 363) + 362]) & mem_q[(k * 363) + 200]) & (mem_q[(k * 363) + 361] == ariane_pkg_is_rs1_fpr(issue_instr_o[289-:7]));
			assign rs2_fwd_req[k + NR_WB_PORTS] = (((mem_q[(k * 363) + 270-:6] == rs2_i) & mem_q[(k * 363) + 362]) & mem_q[(k * 363) + 200]) & (mem_q[(k * 363) + 361] == ariane_pkg_is_rs2_fpr(issue_instr_o[289-:7]));
			assign rs3_fwd_req[k + NR_WB_PORTS] = (((mem_q[(k * 363) + 270-:6] == rs3_i) & mem_q[(k * 363) + 362]) & mem_q[(k * 363) + 200]) & (mem_q[(k * 363) + 361] == ariane_pkg_is_imm_fpr(issue_instr_o[289-:7]));
			assign rs_data[(k + NR_WB_PORTS) * 64+:64] = mem_q[(k * 363) + 264-:64];
		end
	endgenerate
	assign rs1_valid_o = rs1_valid & (|rs1_i | ariane_pkg_is_rs1_fpr(issue_instr_o[289-:7]));
	assign rs2_valid_o = rs2_valid & (|rs2_i | ariane_pkg_is_rs2_fpr(issue_instr_o[289-:7]));
	localparam [31:0] sv2v_uu_i_sel_rs1_NumIn = NR_ENTRIES + NR_WB_PORTS;
	localparam [$clog2(sv2v_uu_i_sel_rs1_NumIn) - 1:0] sv2v_uu_i_sel_rs1_ext_rr_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NR_ENTRIES + NR_WB_PORTS),
		.DataWidth(riscv_XLEN),
		.ExtPrio(1'b1),
		.AxiVldRdy(1'b1)
	) i_sel_rs1(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.rr_i(sv2v_uu_i_sel_rs1_ext_rr_i_0),
		.req_i(rs1_fwd_req),
		.gnt_o(),
		.data_i(rs_data),
		.gnt_i(1'b1),
		.req_o(rs1_valid),
		.data_o(rs1_o),
		.idx_o()
	);
	localparam [31:0] sv2v_uu_i_sel_rs2_NumIn = NR_ENTRIES + NR_WB_PORTS;
	localparam [$clog2(sv2v_uu_i_sel_rs2_NumIn) - 1:0] sv2v_uu_i_sel_rs2_ext_rr_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NR_ENTRIES + NR_WB_PORTS),
		.DataWidth(riscv_XLEN),
		.ExtPrio(1'b1),
		.AxiVldRdy(1'b1)
	) i_sel_rs2(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.rr_i(sv2v_uu_i_sel_rs2_ext_rr_i_0),
		.req_i(rs2_fwd_req),
		.gnt_o(),
		.data_i(rs_data),
		.gnt_i(1'b1),
		.req_o(rs2_valid),
		.data_o(rs2_o),
		.idx_o()
	);
	wire [63:0] rs3;
	localparam [31:0] sv2v_uu_i_sel_rs3_NumIn = NR_ENTRIES + NR_WB_PORTS;
	localparam [$clog2(sv2v_uu_i_sel_rs3_NumIn) - 1:0] sv2v_uu_i_sel_rs3_ext_rr_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NR_ENTRIES + NR_WB_PORTS),
		.DataWidth(riscv_XLEN),
		.ExtPrio(1'b1),
		.AxiVldRdy(1'b1)
	) i_sel_rs3(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.rr_i(sv2v_uu_i_sel_rs3_ext_rr_i_0),
		.req_i(rs3_fwd_req),
		.gnt_o(),
		.data_i(rs_data),
		.gnt_i(1'b1),
		.req_o(rs3_valid_o),
		.data_o(rs3),
		.idx_o()
	);
	assign rs3_o = rs3[ariane_pkg_FLEN - 1:0];
	always @(posedge clk_i or negedge rst_ni) begin : regs
		if (!rst_ni) begin
			mem_q <= {NR_ENTRIES {363'd0}};
			issue_cnt_q <= 1'sb0;
			commit_pointer_q <= 1'sb0;
			issue_pointer_q <= 1'sb0;
		end
		else begin
			issue_cnt_q <= issue_cnt_n;
			issue_pointer_q <= issue_pointer_n;
			mem_q <= mem_n;
			commit_pointer_q <= commit_pointer_n;
		end
	end
endmodule
module serdiv (
	clk_i,
	rst_ni,
	id_i,
	op_a_i,
	op_b_i,
	opcode_i,
	in_vld_i,
	in_rdy_o,
	flush_i,
	out_vld_o,
	out_rdy_i,
	id_o,
	res_o
);
	parameter WIDTH = 64;
	input wire clk_i;
	input wire rst_ni;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	input wire [2:0] id_i;
	input wire [WIDTH - 1:0] op_a_i;
	input wire [WIDTH - 1:0] op_b_i;
	input wire [1:0] opcode_i;
	input wire in_vld_i;
	output reg in_rdy_o;
	input wire flush_i;
	output reg out_vld_o;
	input wire out_rdy_i;
	output wire [2:0] id_o;
	output wire [WIDTH - 1:0] res_o;
	reg [1:0] state_d;
	reg [1:0] state_q;
	reg [WIDTH - 1:0] res_q;
	wire [WIDTH - 1:0] res_d;
	reg [WIDTH - 1:0] op_a_q;
	wire [WIDTH - 1:0] op_a_d;
	reg [WIDTH - 1:0] op_b_q;
	wire [WIDTH - 1:0] op_b_d;
	wire op_a_sign;
	wire op_b_sign;
	wire op_b_zero;
	reg op_b_zero_q;
	wire op_b_zero_d;
	reg [2:0] id_q;
	wire [2:0] id_d;
	wire rem_sel_d;
	reg rem_sel_q;
	wire comp_inv_d;
	reg comp_inv_q;
	wire res_inv_d;
	reg res_inv_q;
	wire [WIDTH - 1:0] add_mux;
	wire [WIDTH - 1:0] add_out;
	wire [WIDTH - 1:0] add_tmp;
	wire [WIDTH - 1:0] b_mux;
	wire [WIDTH - 1:0] out_mux;
	reg [$clog2(WIDTH + 1) - 1:0] cnt_q;
	wire [$clog2(WIDTH + 1) - 1:0] cnt_d;
	wire cnt_zero;
	wire [WIDTH - 1:0] lzc_a_input;
	wire [WIDTH - 1:0] lzc_b_input;
	wire [WIDTH - 1:0] op_b;
	wire [$clog2(WIDTH) - 1:0] lzc_a_result;
	wire [$clog2(WIDTH) - 1:0] lzc_b_result;
	wire [$clog2(WIDTH + 1) - 1:0] shift_a;
	wire [$clog2(WIDTH + 1):0] div_shift;
	reg a_reg_en;
	reg b_reg_en;
	reg res_reg_en;
	wire ab_comp;
	wire pm_sel;
	reg load_en;
	wire lzc_a_no_one;
	wire lzc_b_no_one;
	wire div_res_zero_d;
	reg div_res_zero_q;
	assign op_b_zero = op_b_i == 0;
	assign op_a_sign = op_a_i[WIDTH - 1];
	assign op_b_sign = op_b_i[WIDTH - 1];
	assign lzc_a_input = (opcode_i[0] & op_a_sign ? {~op_a_i, 1'b0} : op_a_i);
	assign lzc_b_input = (opcode_i[0] & op_b_sign ? ~op_b_i : op_b_i);
	lzc #(
		.MODE(1),
		.WIDTH(WIDTH)
	) i_lzc_a(
		.in_i(lzc_a_input),
		.cnt_o(lzc_a_result),
		.empty_o(lzc_a_no_one)
	);
	lzc #(
		.MODE(1),
		.WIDTH(WIDTH)
	) i_lzc_b(
		.in_i(lzc_b_input),
		.cnt_o(lzc_b_result),
		.empty_o(lzc_b_no_one)
	);
	assign shift_a = (lzc_a_no_one ? WIDTH : lzc_a_result);
	assign div_shift = (lzc_b_no_one ? WIDTH : lzc_b_result - shift_a);
	assign op_b = op_b_i <<< $unsigned(div_shift);
	assign div_res_zero_d = (load_en ? $signed(div_shift) < 0 : div_res_zero_q);
	assign pm_sel = load_en & ~(opcode_i[0] & (op_a_sign ^ op_b_sign));
	assign add_mux = (load_en ? op_a_i : op_b_q);
	assign b_mux = (load_en ? op_b : {comp_inv_q, op_b_q[WIDTH - 1:1]});
	assign out_mux = (rem_sel_q ? op_a_q : res_q);
	assign res_o = (res_inv_q ? -$signed(out_mux) : out_mux);
	assign ab_comp = ((op_a_q == op_b_q) | ((op_a_q > op_b_q) ^ comp_inv_q)) & (|op_a_q | op_b_zero_q);
	assign add_tmp = (load_en ? 0 : op_a_q);
	assign add_out = (pm_sel ? add_tmp + add_mux : add_tmp - $signed(add_mux));
	assign cnt_zero = cnt_q == 0;
	assign cnt_d = (load_en ? div_shift : (~cnt_zero ? cnt_q - 1 : cnt_q));
	always @(*) begin : p_fsm
		state_d = state_q;
		in_rdy_o = 1'b0;
		out_vld_o = 1'b0;
		load_en = 1'b0;
		a_reg_en = 1'b0;
		b_reg_en = 1'b0;
		res_reg_en = 1'b0;
		case (state_q)
			2'd0: begin
				in_rdy_o = 1'b1;
				if (in_vld_i) begin
					in_rdy_o = 1'b0;
					a_reg_en = 1'b1;
					b_reg_en = 1'b1;
					load_en = 1'b1;
					state_d = 2'd1;
				end
			end
			2'd1: begin
				if (~div_res_zero_q) begin
					a_reg_en = ab_comp;
					b_reg_en = 1'b1;
					res_reg_en = 1'b1;
				end
				if (div_res_zero_q) begin
					out_vld_o = 1'b1;
					state_d = 2'd2;
					if (out_rdy_i)
						state_d = 2'd0;
				end
				else if (cnt_zero)
					state_d = 2'd2;
			end
			2'd2: begin
				out_vld_o = 1'b1;
				if (out_rdy_i)
					state_d = 2'd0;
			end
			default: state_d = 2'd0;
		endcase
		if (flush_i) begin
			in_rdy_o = 1'b0;
			out_vld_o = 1'b0;
			a_reg_en = 1'b0;
			b_reg_en = 1'b0;
			load_en = 1'b0;
			state_d = 2'd0;
		end
	end
	assign rem_sel_d = (load_en ? opcode_i[1] : rem_sel_q);
	assign comp_inv_d = (load_en ? opcode_i[0] & op_b_sign : comp_inv_q);
	assign op_b_zero_d = (load_en ? op_b_zero : op_b_zero_q);
	assign res_inv_d = (load_en ? ((~op_b_zero | opcode_i[1]) & opcode_i[0]) & (op_a_sign ^ op_b_sign) : res_inv_q);
	assign id_d = (load_en ? id_i : id_q);
	assign id_o = id_q;
	assign op_a_d = (a_reg_en ? add_out : op_a_q);
	assign op_b_d = (b_reg_en ? b_mux : op_b_q);
	assign res_d = (load_en ? {WIDTH {1'sb0}} : (res_reg_en ? {res_q[WIDTH - 2:0], ab_comp} : res_q));
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (~rst_ni) begin
			state_q <= 2'd0;
			op_a_q <= 1'sb0;
			op_b_q <= 1'sb0;
			res_q <= 1'sb0;
			cnt_q <= 1'sb0;
			id_q <= 1'sb0;
			rem_sel_q <= 1'b0;
			comp_inv_q <= 1'b0;
			res_inv_q <= 1'b0;
			op_b_zero_q <= 1'b0;
			div_res_zero_q <= 1'b0;
		end
		else begin
			state_q <= state_d;
			op_a_q <= op_a_d;
			op_b_q <= op_b_d;
			res_q <= res_d;
			cnt_q <= cnt_d;
			id_q <= id_d;
			rem_sel_q <= rem_sel_d;
			comp_inv_q <= comp_inv_d;
			res_inv_q <= res_inv_d;
			op_b_zero_q <= op_b_zero_d;
			div_res_zero_q <= div_res_zero_d;
		end
	end
endmodule
module store_buffer (
	clk_i,
	rst_ni,
	flush_i,
	no_st_pending_o,
	store_buffer_empty_o,
	page_offset_i,
	page_offset_matches_o,
	commit_i,
	commit_ready_o,
	ready_o,
	valid_i,
	valid_without_flush_i,
	paddr_i,
	data_i,
	be_i,
	data_size_i,
	req_port_i,
	req_port_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	output reg no_st_pending_o;
	output wire store_buffer_empty_o;
	input wire [11:0] page_offset_i;
	output reg page_offset_matches_o;
	input wire commit_i;
	output reg commit_ready_o;
	output reg ready_o;
	input wire valid_i;
	input wire valid_without_flush_i;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	input wire [55:0] paddr_i;
	input wire [63:0] data_i;
	input wire [7:0] be_i;
	input wire [1:0] data_size_i;
	input wire [65:0] req_port_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output reg [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_o;
	localparam [31:0] ariane_pkg_DEPTH_SPEC = 4;
	reg [523:0] speculative_queue_n;
	reg [523:0] speculative_queue_q;
	localparam [31:0] ariane_pkg_DEPTH_COMMIT = 4;
	reg [523:0] commit_queue_n;
	reg [523:0] commit_queue_q;
	reg [2:0] speculative_status_cnt_n;
	reg [2:0] speculative_status_cnt_q;
	reg [2:0] commit_status_cnt_n;
	reg [2:0] commit_status_cnt_q;
	reg [1:0] speculative_read_pointer_n;
	reg [1:0] speculative_read_pointer_q;
	reg [1:0] speculative_write_pointer_n;
	reg [1:0] speculative_write_pointer_q;
	reg [1:0] commit_read_pointer_n;
	reg [1:0] commit_read_pointer_q;
	reg [1:0] commit_write_pointer_n;
	reg [1:0] commit_write_pointer_q;
	assign store_buffer_empty_o = (speculative_status_cnt_q == 0) & no_st_pending_o;
	always @(*) begin : core_if
		reg [ariane_pkg_DEPTH_SPEC:0] speculative_status_cnt;
		speculative_status_cnt = speculative_status_cnt_q;
		ready_o = (speculative_status_cnt_q < 3) || commit_i;
		speculative_status_cnt_n = speculative_status_cnt_q;
		speculative_read_pointer_n = speculative_read_pointer_q;
		speculative_write_pointer_n = speculative_write_pointer_q;
		speculative_queue_n = speculative_queue_q;
		if (valid_i) begin
			speculative_queue_n[(speculative_write_pointer_q * 131) + 130-:56] = paddr_i;
			speculative_queue_n[(speculative_write_pointer_q * 131) + 74-:64] = data_i;
			speculative_queue_n[(speculative_write_pointer_q * 131) + 10-:8] = be_i;
			speculative_queue_n[(speculative_write_pointer_q * 131) + 2-:2] = data_size_i;
			speculative_queue_n[(speculative_write_pointer_q * 131) + 0] = 1'b1;
			speculative_write_pointer_n = speculative_write_pointer_q + 1'b1;
			speculative_status_cnt = speculative_status_cnt + 1;
		end
		if (commit_i) begin
			speculative_queue_n[(speculative_read_pointer_q * 131) + 0] = 1'b0;
			speculative_read_pointer_n = speculative_read_pointer_q + 1'b1;
			speculative_status_cnt = speculative_status_cnt - 1;
		end
		speculative_status_cnt_n = speculative_status_cnt;
		if (flush_i) begin
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < ariane_pkg_DEPTH_SPEC; i = i + 1)
					speculative_queue_n[(i * 131) + 0] = 1'b0;
			end
			speculative_write_pointer_n = speculative_read_pointer_q;
			speculative_status_cnt_n = 'b0;
		end
	end
	wire [1:1] sv2v_tmp_A682E;
	assign sv2v_tmp_A682E = 1'b0;
	always @(*) req_port_o[1] = sv2v_tmp_A682E;
	wire [1:1] sv2v_tmp_19E1C;
	assign sv2v_tmp_19E1C = 1'b1;
	always @(*) req_port_o[12] = sv2v_tmp_19E1C;
	wire [1:1] sv2v_tmp_F170F;
	assign sv2v_tmp_F170F = 1'b0;
	always @(*) req_port_o[0] = sv2v_tmp_F170F;
	wire [12:1] sv2v_tmp_6FE53;
	assign sv2v_tmp_6FE53 = commit_queue_q[(commit_read_pointer_q * 131) + 86-:12];
	always @(*) req_port_o[133-:12] = sv2v_tmp_6FE53;
	wire [44:1] sv2v_tmp_7A7D5;
	assign sv2v_tmp_7A7D5 = commit_queue_q[(commit_read_pointer_q * 131) + (74 + (ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_INDEX_WIDTH))-:(74 + (ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_INDEX_WIDTH)) - 86];
	always @(*) req_port_o[121-:44] = sv2v_tmp_7A7D5;
	wire [64:1] sv2v_tmp_8BEAD;
	assign sv2v_tmp_8BEAD = (req_port_o[124] == 1'b0 ? {commit_queue_q[(commit_read_pointer_q * 131) + 74-:64]} : {commit_queue_q[(commit_read_pointer_q * 131) + 74-:64]});
	always @(*) req_port_o[77-:64] = sv2v_tmp_8BEAD;
	wire [8:1] sv2v_tmp_6B135;
	assign sv2v_tmp_6B135 = commit_queue_q[(commit_read_pointer_q * 131) + 10-:8];
	always @(*) req_port_o[11-:8] = sv2v_tmp_6B135;
	wire [2:1] sv2v_tmp_13B79;
	assign sv2v_tmp_13B79 = commit_queue_q[(commit_read_pointer_q * 131) + 2-:2];
	always @(*) req_port_o[3-:2] = sv2v_tmp_13B79;
	always @(*) begin : store_if
		reg [ariane_pkg_DEPTH_COMMIT:0] commit_status_cnt;
		commit_status_cnt = commit_status_cnt_q;
		commit_ready_o = commit_status_cnt_q < ariane_pkg_DEPTH_COMMIT;
		no_st_pending_o = commit_status_cnt_q == 0;
		commit_read_pointer_n = commit_read_pointer_q;
		commit_write_pointer_n = commit_write_pointer_q;
		commit_queue_n = commit_queue_q;
		req_port_o[13] = 1'b0;
		if (commit_queue_q[(commit_read_pointer_q * 131) + 0]) begin
			req_port_o[13] = 1'b1;
			if (req_port_i[65]) begin
				commit_queue_n[(commit_read_pointer_q * 131) + 0] = 1'b0;
				commit_read_pointer_n = commit_read_pointer_q + 1'b1;
				commit_status_cnt = commit_status_cnt - 1;
			end
		end
		if (commit_i) begin
			commit_queue_n[0 + (commit_write_pointer_q * 131)+:131] = speculative_queue_q[0 + (speculative_read_pointer_q * 131)+:131];
			commit_write_pointer_n = commit_write_pointer_n + 1'b1;
			commit_status_cnt = commit_status_cnt + 1;
		end
		commit_status_cnt_n = commit_status_cnt;
	end
	always @(*) begin : sv2v_autoblock_2
		reg [0:1] _sv2v_jump;
		_sv2v_jump = 2'b00;
		begin : address_checker
			page_offset_matches_o = 1'b0;
			begin : sv2v_autoblock_3
				reg [31:0] i;
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < ariane_pkg_DEPTH_COMMIT; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if ((page_offset_i[11:3] == commit_queue_q[(i * 131) + 86-:9]) && commit_queue_q[(i * 131) + 0]) begin
								page_offset_matches_o = 1'b1;
								_sv2v_jump = 2'b10;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				begin : sv2v_autoblock_5
					reg [31:0] i;
					begin : sv2v_autoblock_6
						reg [31:0] _sv2v_value_on_break;
						for (i = 0; i < ariane_pkg_DEPTH_SPEC; i = i + 1)
							if (_sv2v_jump < 2'b10) begin
								_sv2v_jump = 2'b00;
								if ((page_offset_i[11:3] == speculative_queue_q[(i * 131) + 86-:9]) && speculative_queue_q[(i * 131) + 0]) begin
									page_offset_matches_o = 1'b1;
									_sv2v_jump = 2'b10;
								end
								_sv2v_value_on_break = i;
							end
						if (!(_sv2v_jump < 2'b10))
							i = _sv2v_value_on_break;
						if (_sv2v_jump != 2'b11)
							_sv2v_jump = 2'b00;
					end
				end
				if (_sv2v_jump == 2'b00) begin
					if ((page_offset_i[11:3] == paddr_i[11:3]) && valid_without_flush_i)
						page_offset_matches_o = 1'b1;
				end
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_spec
		if (~rst_ni) begin
			speculative_queue_q <= {ariane_pkg_DEPTH_SPEC {131'd0}};
			speculative_read_pointer_q <= 1'sb0;
			speculative_write_pointer_q <= 1'sb0;
			speculative_status_cnt_q <= 1'sb0;
		end
		else begin
			speculative_queue_q <= speculative_queue_n;
			speculative_read_pointer_q <= speculative_read_pointer_n;
			speculative_write_pointer_q <= speculative_write_pointer_n;
			speculative_status_cnt_q <= speculative_status_cnt_n;
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_commit
		if (~rst_ni) begin
			commit_queue_q <= {ariane_pkg_DEPTH_COMMIT {131'd0}};
			commit_read_pointer_q <= 1'sb0;
			commit_write_pointer_q <= 1'sb0;
			commit_status_cnt_q <= 1'sb0;
		end
		else begin
			commit_queue_q <= commit_queue_n;
			commit_read_pointer_q <= commit_read_pointer_n;
			commit_write_pointer_q <= commit_write_pointer_n;
			commit_status_cnt_q <= commit_status_cnt_n;
		end
	end
endmodule
module store_unit (
	clk_i,
	rst_ni,
	flush_i,
	no_st_pending_o,
	store_buffer_empty_o,
	valid_i,
	lsu_ctrl_i,
	pop_st_o,
	commit_i,
	commit_ready_o,
	amo_valid_commit_i,
	valid_o,
	trans_id_o,
	result_o,
	ex_o,
	translation_req_o,
	vaddr_o,
	paddr_i,
	ex_i,
	dtlb_hit_i,
	page_offset_i,
	page_offset_matches_o,
	amo_req_o,
	amo_resp_i,
	req_port_i,
	req_port_o
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	output wire no_st_pending_o;
	output wire store_buffer_empty_o;
	input wire valid_i;
	localparam ariane_pkg_NR_SB_ENTRIES = 8;
	localparam ariane_pkg_TRANS_ID_BITS = 3;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [151:0] lsu_ctrl_i;
	output reg pop_st_o;
	input wire commit_i;
	output wire commit_ready_o;
	input wire amo_valid_commit_i;
	output reg valid_o;
	output wire [2:0] trans_id_o;
	output wire [63:0] result_o;
	output reg [128:0] ex_o;
	output reg translation_req_o;
	output wire [63:0] vaddr_o;
	localparam riscv_PLEN = 56;
	input wire [55:0] paddr_i;
	input wire [128:0] ex_i;
	input wire dtlb_hit_i;
	input wire [11:0] page_offset_i;
	output wire page_offset_matches_o;
	output wire [134:0] amo_req_o;
	input wire [64:0] amo_resp_i;
	input wire [65:0] req_port_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output wire [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_o;
	assign result_o = 1'sb0;
	reg [1:0] state_d;
	reg [1:0] state_q;
	wire st_ready;
	reg st_valid;
	reg st_valid_without_flush;
	wire instr_is_amo;
	function automatic ariane_pkg_is_amo;
		input reg [6:0] op;
		if ((7'd46 <= op) && (7'd67 >= op))
			ariane_pkg_is_amo = 1'b1;
		else
			ariane_pkg_is_amo = 1'b0;
	endfunction
	assign instr_is_amo = ariane_pkg_is_amo(lsu_ctrl_i[9-:7]);
	reg [63:0] st_data_n;
	reg [63:0] st_data_q;
	reg [7:0] st_be_n;
	reg [7:0] st_be_q;
	reg [1:0] st_data_size_n;
	reg [1:0] st_data_size_q;
	reg [3:0] amo_op_d;
	reg [3:0] amo_op_q;
	reg [2:0] trans_id_n;
	reg [2:0] trans_id_q;
	assign vaddr_o = lsu_ctrl_i[150-:64];
	assign trans_id_o = trans_id_q;
	always @(*) begin : store_control
		translation_req_o = 1'b0;
		valid_o = 1'b0;
		st_valid = 1'b0;
		st_valid_without_flush = 1'b0;
		pop_st_o = 1'b0;
		ex_o = ex_i;
		trans_id_n = lsu_ctrl_i[2-:ariane_pkg_TRANS_ID_BITS];
		state_d = state_q;
		case (state_q)
			2'd0:
				if (valid_i) begin
					state_d = 2'd1;
					translation_req_o = 1'b1;
					pop_st_o = 1'b1;
					if (!dtlb_hit_i) begin
						state_d = 2'd2;
						pop_st_o = 1'b0;
					end
					if (!st_ready) begin
						state_d = 2'd3;
						pop_st_o = 1'b0;
					end
				end
			2'd1: begin
				valid_o = 1'b1;
				if (!flush_i)
					st_valid = 1'b1;
				st_valid_without_flush = 1'b1;
				if (valid_i && !instr_is_amo) begin
					translation_req_o = 1'b1;
					state_d = 2'd1;
					pop_st_o = 1'b1;
					if (!dtlb_hit_i) begin
						state_d = 2'd2;
						pop_st_o = 1'b0;
					end
					if (!st_ready) begin
						state_d = 2'd3;
						pop_st_o = 1'b0;
					end
				end
				else
					state_d = 2'd0;
			end
			2'd3: begin
				translation_req_o = 1'b1;
				if (st_ready && dtlb_hit_i)
					state_d = 2'd0;
			end
			2'd2: begin
				translation_req_o = 1'b1;
				if (dtlb_hit_i)
					state_d = 2'd0;
			end
		endcase
		if (ex_i[0] && (state_q != 2'd0)) begin
			pop_st_o = 1'b1;
			st_valid = 1'b0;
			state_d = 2'd0;
			valid_o = 1'b1;
		end
		if (flush_i)
			state_d = 2'd0;
	end
	localparam riscv_IS_XLEN64 = 1'b1;
	function automatic [63:0] ariane_pkg_data_align;
		input reg [2:0] addr;
		input reg [63:0] data;
		reg [2:0] addr_tmp;
		reg [63:0] data_tmp;
		begin
			addr_tmp = {addr[2] && riscv_IS_XLEN64, addr[1:0]};
			data_tmp = {64 {1'b0}};
			case (addr_tmp)
				3'b000: data_tmp[63:0] = {data[63:0]};
				3'b001: data_tmp[63:0] = {data[55:0], data[63:56]};
				3'b010: data_tmp[63:0] = {data[47:0], data[63:48]};
				3'b011: data_tmp[63:0] = {data[39:0], data[63:40]};
				3'b100: data_tmp = {data[31:0], data[63:32]};
				3'b101: data_tmp = {data[23:0], data[63:24]};
				3'b110: data_tmp = {data[15:0], data[63:16]};
				3'b111: data_tmp = {data[7:0], data[63:8]};
			endcase
			ariane_pkg_data_align = data_tmp[63:0];
		end
	endfunction
	function automatic [1:0] ariane_pkg_extract_transfer_size;
		input reg [6:0] op;
		case (op)
			7'd35, 7'd36, 7'd81, 7'd85, 7'd47, 7'd49, 7'd59, 7'd60, 7'd61, 7'd62, 7'd63, 7'd64, 7'd65, 7'd66, 7'd67: ariane_pkg_extract_transfer_size = 2'b11;
			7'd37, 7'd38, 7'd39, 7'd82, 7'd86, 7'd46, 7'd48, 7'd50, 7'd51, 7'd52, 7'd53, 7'd54, 7'd55, 7'd56, 7'd57, 7'd58: ariane_pkg_extract_transfer_size = 2'b10;
			7'd40, 7'd41, 7'd42, 7'd83, 7'd87: ariane_pkg_extract_transfer_size = 2'b01;
			7'd43, 7'd45, 7'd44, 7'd84, 7'd88: ariane_pkg_extract_transfer_size = 2'b00;
			default: ariane_pkg_extract_transfer_size = 2'b11;
		endcase
	endfunction
	always @(*) begin
		st_be_n = lsu_ctrl_i[21-:8];
		st_data_n = (instr_is_amo ? lsu_ctrl_i[85:22] : ariane_pkg_data_align(lsu_ctrl_i[89:87], {lsu_ctrl_i[85:22]}));
		st_data_size_n = ariane_pkg_extract_transfer_size(lsu_ctrl_i[9-:7]);
		case (lsu_ctrl_i[9-:7])
			7'd46, 7'd47: amo_op_d = 4'b0001;
			7'd48, 7'd49: amo_op_d = 4'b0010;
			7'd50, 7'd59: amo_op_d = 4'b0011;
			7'd51, 7'd60: amo_op_d = 4'b0100;
			7'd52, 7'd61: amo_op_d = 4'b0101;
			7'd53, 7'd62: amo_op_d = 4'b0110;
			7'd54, 7'd63: amo_op_d = 4'b0111;
			7'd55, 7'd64: amo_op_d = 4'b1000;
			7'd56, 7'd65: amo_op_d = 4'b1001;
			7'd57, 7'd66: amo_op_d = 4'b1010;
			7'd58, 7'd67: amo_op_d = 4'b1011;
			default: amo_op_d = 4'b0000;
		endcase
	end
	wire store_buffer_valid;
	wire amo_buffer_valid;
	wire store_buffer_ready;
	wire amo_buffer_ready;
	assign store_buffer_valid = st_valid & (amo_op_q == 4'b0000);
	assign amo_buffer_valid = st_valid & (amo_op_q != 4'b0000);
	assign st_ready = store_buffer_ready & amo_buffer_ready;
	store_buffer store_buffer_i(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.no_st_pending_o(no_st_pending_o),
		.store_buffer_empty_o(store_buffer_empty_o),
		.page_offset_i(page_offset_i),
		.page_offset_matches_o(page_offset_matches_o),
		.commit_i(commit_i),
		.commit_ready_o(commit_ready_o),
		.ready_o(store_buffer_ready),
		.valid_i(store_buffer_valid),
		.valid_without_flush_i(st_valid_without_flush),
		.paddr_i(paddr_i),
		.data_i(st_data_q),
		.be_i(st_be_q),
		.data_size_i(st_data_size_q),
		.req_port_i(req_port_i),
		.req_port_o(req_port_o)
	);
	amo_buffer i_amo_buffer(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.valid_i(amo_buffer_valid),
		.ready_o(amo_buffer_ready),
		.paddr_i(paddr_i),
		.amo_op_i(amo_op_q),
		.data_i(st_data_q),
		.data_size_i(st_data_size_q),
		.amo_req_o(amo_req_o),
		.amo_resp_i(amo_resp_i),
		.amo_valid_commit_i(amo_valid_commit_i),
		.no_st_pending_i(no_st_pending_o)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			state_q <= 2'd0;
			st_be_q <= 1'sb0;
			st_data_q <= 1'sb0;
			st_data_size_q <= 1'sb0;
			trans_id_q <= 1'sb0;
			amo_op_q <= 4'b0000;
		end
		else begin
			state_q <= state_d;
			st_be_q <= st_be_n;
			st_data_q <= st_data_n;
			trans_id_q <= trans_id_n;
			st_data_size_q <= st_data_size_n;
			amo_op_q <= amo_op_d;
		end
endmodule
module tlb (
	clk_i,
	rst_ni,
	flush_i,
	update_i,
	lu_access_i,
	lu_asid_i,
	lu_vaddr_i,
	lu_content_o,
	asid_to_be_flushed_i,
	vaddr_to_be_flushed_i,
	lu_is_2M_o,
	lu_is_1G_o,
	lu_hit_o
);
	parameter [31:0] TLB_ENTRIES = 4;
	parameter [31:0] ASID_WIDTH = 1;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam riscv_XLEN = 64;
	localparam ariane_pkg_ASID_WIDTH = 16;
	localparam riscv_PLEN = 56;
	input wire [109:0] update_i;
	input wire lu_access_i;
	input wire [ASID_WIDTH - 1:0] lu_asid_i;
	localparam riscv_VLEN = 64;
	input wire [63:0] lu_vaddr_i;
	output reg [63:0] lu_content_o;
	input wire [ASID_WIDTH - 1:0] asid_to_be_flushed_i;
	input wire [63:0] vaddr_to_be_flushed_i;
	output reg lu_is_2M_o;
	output reg lu_is_1G_o;
	output reg lu_hit_o;
	localparam riscv_VPN2 = 8;
	reg [((ASID_WIDTH + 29) >= 0 ? (TLB_ENTRIES * (ASID_WIDTH + 30)) - 1 : (TLB_ENTRIES * (1 - (ASID_WIDTH + 29))) + (ASID_WIDTH + 28)):((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] tags_q;
	reg [((ASID_WIDTH + 29) >= 0 ? (TLB_ENTRIES * (ASID_WIDTH + 30)) - 1 : (TLB_ENTRIES * (1 - (ASID_WIDTH + 29))) + (ASID_WIDTH + 28)):((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] tags_n;
	reg [(TLB_ENTRIES * 64) - 1:0] content_q;
	reg [(TLB_ENTRIES * 64) - 1:0] content_n;
	reg [8:0] vpn0;
	reg [8:0] vpn1;
	reg [riscv_VPN2:0] vpn2;
	reg [TLB_ENTRIES - 1:0] lu_hit;
	reg [TLB_ENTRIES - 1:0] replace_en;
	function automatic [43:0] sv2v_cast_768E8;
		input reg [43:0] inp;
		sv2v_cast_768E8 = inp;
	endfunction
	always @(*) begin : translation
		vpn0 = lu_vaddr_i[20:12];
		vpn1 = lu_vaddr_i[29:21];
		vpn2 = lu_vaddr_i[38:30];
		lu_hit = {TLB_ENTRIES {1'd0}};
		lu_hit_o = 1'b0;
		lu_content_o = {10'd0, sv2v_cast_768E8(0), 10'h000};
		lu_is_1G_o = 1'b0;
		lu_is_2M_o = 1'b0;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				if ((tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] && ((lu_asid_i == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29)) : (((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))) - 1)-:((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))]) || content_q[(i * 64) + 5])) && (vpn2 == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 29 : ASID_WIDTH + 0) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 29 : ASID_WIDTH + 0)) + 8)-:9])) begin
					if (tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 1 : ASID_WIDTH + 28)]) begin
						lu_is_1G_o = 1'b1;
						lu_content_o = content_q[0 + (i * 64)+:64];
						lu_hit_o = 1'b1;
						lu_hit[i] = 1'b1;
					end
					else if (vpn1 == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 20 : ASID_WIDTH + 9) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 20 : ASID_WIDTH + 9)) + 8)-:9]) begin
						if (tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 2 : ASID_WIDTH + 27)] || (vpn0 == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 11 : ASID_WIDTH + 18) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 11 : ASID_WIDTH + 18)) + 8)-:9])) begin
							lu_is_2M_o = tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 2 : ASID_WIDTH + 27)];
							lu_content_o = content_q[0 + (i * 64)+:64];
							lu_hit_o = 1'b1;
							lu_hit[i] = 1'b1;
						end
					end
				end
		end
	end
	wire asid_to_be_flushed_is0;
	wire vaddr_to_be_flushed_is0;
	reg [TLB_ENTRIES - 1:0] vaddr_vpn0_match;
	reg [TLB_ENTRIES - 1:0] vaddr_vpn1_match;
	reg [TLB_ENTRIES - 1:0] vaddr_vpn2_match;
	assign asid_to_be_flushed_is0 = ~(|asid_to_be_flushed_i);
	assign vaddr_to_be_flushed_is0 = ~(|vaddr_to_be_flushed_i);
	function automatic [ASID_WIDTH - 1:0] sv2v_cast_E5F2C;
		input reg [ASID_WIDTH - 1:0] inp;
		sv2v_cast_E5F2C = inp;
	endfunction
	function automatic [8:0] sv2v_cast_8667A;
		input reg [8:0] inp;
		sv2v_cast_8667A = inp;
	endfunction
	always @(*) begin : update_flush
		tags_n = tags_q;
		content_n = content_q;
		begin : sv2v_autoblock_2
			reg [31:0] i;
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin
					vaddr_vpn0_match[i] = vaddr_to_be_flushed_i[20:12] == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 11 : ASID_WIDTH + 18) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 11 : ASID_WIDTH + 18)) + 8)-:9];
					vaddr_vpn1_match[i] = vaddr_to_be_flushed_i[29:21] == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 20 : ASID_WIDTH + 9) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 20 : ASID_WIDTH + 9)) + 8)-:9];
					vaddr_vpn2_match[i] = vaddr_to_be_flushed_i[38:30] == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 29 : ASID_WIDTH + 0) : ((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 29 : ASID_WIDTH + 0)) + 8)-:9];
					if (flush_i) begin
						if (asid_to_be_flushed_is0 && vaddr_to_be_flushed_is0)
							tags_n[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] = 1'b0;
						else if ((asid_to_be_flushed_is0 && ((((vaddr_vpn0_match[i] && vaddr_vpn1_match[i]) && vaddr_vpn2_match[i]) || (vaddr_vpn2_match[i] && tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 1 : ASID_WIDTH + 28)])) || ((vaddr_vpn1_match[i] && vaddr_vpn2_match[i]) && tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 2 : ASID_WIDTH + 27)]))) && ~vaddr_to_be_flushed_is0)
							tags_n[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] = 1'b0;
						else if ((((!content_q[(i * 64) + 5] && ((((vaddr_vpn0_match[i] && vaddr_vpn1_match[i]) && vaddr_vpn2_match[i]) || (vaddr_vpn2_match[i] && tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 1 : ASID_WIDTH + 28)])) || ((vaddr_vpn1_match[i] && vaddr_vpn2_match[i]) && tags_q[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 2 : ASID_WIDTH + 27)]))) && (asid_to_be_flushed_i == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29)) : (((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))) - 1)-:((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))])) && !vaddr_to_be_flushed_is0) && !asid_to_be_flushed_is0)
							tags_n[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] = 1'b0;
						else if (((!content_q[(i * 64) + 5] && vaddr_to_be_flushed_is0) && (asid_to_be_flushed_i == tags_q[((ASID_WIDTH + 29) >= 0 ? (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29)) : (((i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 29 : (ASID_WIDTH + 29) - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))) - 1)-:((ASID_WIDTH + 29) >= 30 ? ASID_WIDTH : 31 - (ASID_WIDTH + 29))])) && !asid_to_be_flushed_is0)
							tags_n[(i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))) + ((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29)] = 1'b0;
					end
					else if (update_i[109] & replace_en[i]) begin
						tags_n[((ASID_WIDTH + 29) >= 0 ? 0 : ASID_WIDTH + 29) + (i * ((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29)))+:((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29))] = {sv2v_cast_E5F2C(update_i[79-:16]), sv2v_cast_8667A(update_i[106:98]), update_i[97:89], update_i[88:80], update_i[108], update_i[107], 1'b1};
						content_n[0 + (i * 64)+:64] = update_i[63-:64];
					end
				end
		end
	end
	reg [(2 * (TLB_ENTRIES - 1)) - 1:0] plru_tree_q;
	reg [(2 * (TLB_ENTRIES - 1)) - 1:0] plru_tree_n;
	always @(*) begin : plru_replacement
		plru_tree_n = plru_tree_q;
		begin : sv2v_autoblock_3
			reg [31:0] i;
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin : sv2v_autoblock_4
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					if (lu_hit[i] & lu_access_i) begin : sv2v_autoblock_5
						reg [31:0] lvl;
						for (lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl = lvl + 1)
							begin
								idx_base = $unsigned((2 ** lvl) - 1);
								shift = $clog2(TLB_ENTRIES) - lvl;
								new_index = ~((i >> (shift - 1)) & 32'b00000000000000000000000000000001);
								plru_tree_n[idx_base + (i >> shift)] = new_index[0];
							end
					end
				end
		end
		begin : sv2v_autoblock_6
			reg [31:0] i;
			for (i = 0; i < TLB_ENTRIES; i = i + 1)
				begin : sv2v_autoblock_7
					reg en;
					reg [31:0] idx_base;
					reg [31:0] shift;
					reg [31:0] new_index;
					en = 1'b1;
					begin : sv2v_autoblock_8
						reg [31:0] lvl;
						for (lvl = 0; lvl < $clog2(TLB_ENTRIES); lvl = lvl + 1)
							begin
								idx_base = $unsigned((2 ** lvl) - 1);
								shift = $clog2(TLB_ENTRIES) - lvl;
								new_index = (i >> (shift - 1)) & 32'b00000000000000000000000000000001;
								if (new_index[0])
									en = en & plru_tree_q[idx_base + (i >> shift)];
								else
									en = en & ~plru_tree_q[idx_base + (i >> shift)];
							end
					end
					replace_en[i] = en;
				end
		end
	end
	function automatic [((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29)) - 1:0] sv2v_cast_296FB;
		input reg [((ASID_WIDTH + 29) >= 0 ? ASID_WIDTH + 30 : 1 - (ASID_WIDTH + 29)) - 1:0] inp;
		sv2v_cast_296FB = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			tags_q <= {TLB_ENTRIES {sv2v_cast_296FB(0)}};
			content_q <= {TLB_ENTRIES {64'd0}};
			plru_tree_q <= {2 * (TLB_ENTRIES - 1) {1'd0}};
		end
		else begin
			tags_q <= tags_n;
			content_q <= content_n;
			plru_tree_q <= plru_tree_n;
		end
endmodule
module fpnew_cast_multi_5BCFE_D3186 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [31:0] AuxType_AUX_BITS = 0;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	parameter [0:4] FpFmtConfig = 1'sb1;
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	parameter [0:3] IntFmtConfig = 1'sb1;
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		input reg [1:0] ifmt;
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		input reg [0:3] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_2
				reg signed [31:0] ifmt;
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					if (cfg[ifmt])
						res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_maximum(fpnew_pkg_max_fp_width(FpFmtConfig), fpnew_pkg_max_int_width(IntFmtConfig));
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	input wire clk_i;
	input wire rst_ni;
	input wire [WIDTH - 1:0] operands_i;
	input wire [4:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	input wire [2:0] src_fmt_i;
	input wire [2:0] dst_fmt_i;
	input wire [1:0] int_fmt_i;
	input wire [2:0] tag_i;
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	function automatic [31:0] fpnew_pkg_exp_bits;
		input reg [2:0] fmt;
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		input reg [2:0] fmt;
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		input reg [0:4] cfg;
		reg [63:0] res;
		begin
			res = 1'sb0;
			begin : sv2v_autoblock_3
				reg [31:0] fmt;
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	localparam [31:0] SUPER_BIAS = (2 ** (SUPER_EXP_BITS - 1)) - 1;
	localparam [31:0] INT_MAN_WIDTH = fpnew_pkg_maximum(SUPER_MAN_BITS + 1, MAX_INT_WIDTH);
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(INT_MAN_WIDTH);
	localparam [31:0] INT_EXP_WIDTH = fpnew_pkg_maximum($clog2(MAX_INT_WIDTH), fpnew_pkg_maximum(SUPER_EXP_BITS, $clog2(SUPER_BIAS + SUPER_MAN_BITS))) + 1;
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	wire [WIDTH - 1:0] operands_q;
	wire [4:0] is_boxed_q;
	wire op_mod_q;
	wire [2:0] src_fmt_q;
	wire [2:0] dst_fmt_q;
	wire [1:0] int_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * WIDTH) + ((NUM_INP_REGS * WIDTH) - 1) : ((NUM_INP_REGS + 1) * WIDTH) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * WIDTH : 0)] inp_pipe_operands_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)] inp_pipe_is_boxed_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] inp_pipe_int_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_tag_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	wire [WIDTH * 1:1] sv2v_tmp_6E45B;
	assign sv2v_tmp_6E45B = operands_i;
	always @(*) inp_pipe_operands_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6E45B;
	wire [5:1] sv2v_tmp_C47E1;
	assign sv2v_tmp_C47E1 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS] = sv2v_tmp_C47E1;
	wire [3:1] sv2v_tmp_45ED9;
	assign sv2v_tmp_45ED9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_45ED9;
	wire [4:1] sv2v_tmp_AD1FB;
	assign sv2v_tmp_AD1FB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_AD1FB;
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	wire [3:1] sv2v_tmp_CB295;
	assign sv2v_tmp_CB295 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_CB295;
	wire [3:1] sv2v_tmp_6AF63;
	assign sv2v_tmp_6AF63 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6AF63;
	wire [2:1] sv2v_tmp_CA55F;
	assign sv2v_tmp_CA55F = int_fmt_i;
	always @(*) inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_CA55F;
	wire [3:1] sv2v_tmp_F99B7;
	assign sv2v_tmp_F99B7 = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_F99B7;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_AA86B;
	assign sv2v_tmp_AA86B = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_AA86B;
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	assign in_ready_o = inp_pipe_ready[0];
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			wire reg_ena;
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * WIDTH+:WIDTH] : inp_pipe_operands_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * WIDTH+:WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= 1'sb0;
				else
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS+:NUM_FORMATS] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS+:NUM_FORMATS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign operands_q = inp_pipe_operands_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * WIDTH+:WIDTH];
	assign is_boxed_q = inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS+:NUM_FORMATS];
	assign op_mod_q = inp_pipe_op_mod_q[NUM_INP_REGS];
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign int_fmt_q = inp_pipe_int_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	wire src_is_int;
	wire dst_is_int;
	assign src_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(12);
	assign dst_is_int = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(11);
	wire [INT_MAN_WIDTH - 1:0] encoded_mant;
	wire [4:0] fmt_sign;
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_exponent;
	wire [(NUM_FORMATS * INT_MAN_WIDTH) - 1:0] fmt_mantissa;
	wire signed [(NUM_FORMATS * INT_EXP_WIDTH) - 1:0] fmt_shift_compensation;
	wire [39:0] info;
	reg [(NUM_INT_FORMATS * INT_MAN_WIDTH) - 1:0] ifmt_input_val;
	wire int_sign;
	wire [INT_MAN_WIDTH - 1:0] int_value;
	wire [INT_MAN_WIDTH - 1:0] int_mantissa;
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [0:0] sv2v_cast_1_signed;
		input reg signed [0:0] inp;
		sv2v_cast_1_signed = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(1)
				) i_fpnew_classifier(
					.operands_i(operands_q[FP_WIDTH - 1:0]),
					.is_boxed_i(is_boxed_q[fmt]),
					.info_o(info[fmt * 8+:8])
				);
				assign fmt_sign[fmt] = operands_q[FP_WIDTH - 1];
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed({1'b0, operands_q[MAN_BITS+:EXP_BITS]});
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {info[(fmt * 8) + 7], operands_q[MAN_BITS - 1:0]};
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = $signed((INT_MAN_WIDTH - 1) - MAN_BITS);
			end
			else begin : inactive_format
				assign info[fmt * 8+:8] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				assign fmt_sign[fmt] = fpnew_pkg_DONT_CARE;
				assign fmt_exponent[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
				assign fmt_mantissa[fmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				assign fmt_shift_compensation[fmt * INT_EXP_WIDTH+:INT_EXP_WIDTH] = {INT_EXP_WIDTH {sv2v_cast_1_signed(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	genvar ifmt;
	function automatic [0:0] sv2v_cast_1;
		input reg [0:0] inp;
		sv2v_cast_1 = inp;
	endfunction
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_sign_extend_int
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				always @(*) begin : sign_ext_input
					ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = {INT_MAN_WIDTH {sv2v_cast_1(operands_q[INT_WIDTH - 1] & ~op_mod_q)}};
					ifmt_input_val[(ifmt * INT_MAN_WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = operands_q[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_5B946;
				assign sv2v_tmp_5B946 = {INT_MAN_WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_input_val[ifmt * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_5B946;
			end
		end
	endgenerate
	assign int_value = ifmt_input_val[int_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	assign int_sign = int_value[INT_MAN_WIDTH - 1] & ~op_mod_q;
	assign int_mantissa = (int_sign ? $unsigned(-int_value) : int_value);
	assign encoded_mant = (src_is_int ? int_mantissa : fmt_mantissa[src_fmt_q * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
	wire signed [INT_EXP_WIDTH - 1:0] src_bias;
	wire signed [INT_EXP_WIDTH - 1:0] src_exp;
	wire signed [INT_EXP_WIDTH - 1:0] src_subnormal;
	wire signed [INT_EXP_WIDTH - 1:0] src_offset;
	function automatic [31:0] fpnew_pkg_bias;
		input reg [2:0] fmt;
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	assign src_bias = $signed(fpnew_pkg_bias(src_fmt_q));
	assign src_exp = fmt_exponent[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	assign src_subnormal = $signed({1'b0, info[(src_fmt_q * 8) + 6]});
	assign src_offset = fmt_shift_compensation[src_fmt_q * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	wire input_sign;
	wire signed [INT_EXP_WIDTH - 1:0] input_exp;
	wire [INT_MAN_WIDTH - 1:0] input_mant;
	wire mant_is_zero;
	wire signed [INT_EXP_WIDTH - 1:0] fp_input_exp;
	wire signed [INT_EXP_WIDTH - 1:0] int_input_exp;
	wire [LZC_RESULT_WIDTH - 1:0] renorm_shamt;
	wire [LZC_RESULT_WIDTH:0] renorm_shamt_sgn;
	lzc #(
		.WIDTH(INT_MAN_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(encoded_mant),
		.cnt_o(renorm_shamt),
		.empty_o(mant_is_zero)
	);
	assign renorm_shamt_sgn = $signed({1'b0, renorm_shamt});
	assign input_sign = (src_is_int ? int_sign : fmt_sign[src_fmt_q]);
	assign input_mant = encoded_mant << renorm_shamt;
	assign fp_input_exp = $signed((((src_exp + src_subnormal) - src_bias) - renorm_shamt_sgn) + src_offset);
	assign int_input_exp = $signed((INT_MAN_WIDTH - 1) - renorm_shamt_sgn);
	assign input_exp = (src_is_int ? int_input_exp : fp_input_exp);
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp;
	assign destination_exp = input_exp + $signed(fpnew_pkg_bias(dst_fmt_q));
	wire input_sign_q;
	wire signed [INT_EXP_WIDTH - 1:0] input_exp_q;
	wire [INT_MAN_WIDTH - 1:0] input_mant_q;
	wire signed [INT_EXP_WIDTH - 1:0] destination_exp_q;
	wire src_is_int_q;
	wire dst_is_int_q;
	wire [7:0] info_q;
	wire mant_is_zero_q;
	wire op_mod_q2;
	wire [2:0] rnd_mode_q;
	wire [2:0] src_fmt_q2;
	wire [2:0] dst_fmt_q2;
	wire [1:0] int_fmt_q2;
	reg [0:NUM_MID_REGS] mid_pipe_input_sign_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_input_exp_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_MAN_WIDTH) + ((NUM_MID_REGS * INT_MAN_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_MAN_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_MAN_WIDTH : 0)] mid_pipe_input_mant_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * INT_EXP_WIDTH) + ((NUM_MID_REGS * INT_EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * INT_EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * INT_EXP_WIDTH : 0)] mid_pipe_dest_exp_q;
	reg [0:NUM_MID_REGS] mid_pipe_src_is_int_q;
	reg [0:NUM_MID_REGS] mid_pipe_dst_is_int_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 8) + ((NUM_MID_REGS * 8) - 1) : ((NUM_MID_REGS + 1) * 8) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 8 : 0)] mid_pipe_info_q;
	reg [0:NUM_MID_REGS] mid_pipe_mant_zero_q;
	reg [0:NUM_MID_REGS] mid_pipe_op_mod_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_src_fmt_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_INT_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_INT_FORMAT_BITS : 0)] mid_pipe_int_fmt_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_tag_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	wire [1:1] sv2v_tmp_3DFAC;
	assign sv2v_tmp_3DFAC = input_sign;
	always @(*) mid_pipe_input_sign_q[0] = sv2v_tmp_3DFAC;
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_9AB08;
	assign sv2v_tmp_9AB08 = input_exp;
	always @(*) mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_9AB08;
	wire [INT_MAN_WIDTH * 1:1] sv2v_tmp_3BE44;
	assign sv2v_tmp_3BE44 = input_mant;
	always @(*) mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH] = sv2v_tmp_3BE44;
	wire [INT_EXP_WIDTH * 1:1] sv2v_tmp_F626F;
	assign sv2v_tmp_F626F = destination_exp;
	always @(*) mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH] = sv2v_tmp_F626F;
	wire [1:1] sv2v_tmp_3D9F8;
	assign sv2v_tmp_3D9F8 = src_is_int;
	always @(*) mid_pipe_src_is_int_q[0] = sv2v_tmp_3D9F8;
	wire [1:1] sv2v_tmp_4E95C;
	assign sv2v_tmp_4E95C = dst_is_int;
	always @(*) mid_pipe_dst_is_int_q[0] = sv2v_tmp_4E95C;
	wire [8:1] sv2v_tmp_48E57;
	assign sv2v_tmp_48E57 = info[src_fmt_q * 8+:8];
	always @(*) mid_pipe_info_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 8+:8] = sv2v_tmp_48E57;
	wire [1:1] sv2v_tmp_4351A;
	assign sv2v_tmp_4351A = mant_is_zero;
	always @(*) mid_pipe_mant_zero_q[0] = sv2v_tmp_4351A;
	wire [1:1] sv2v_tmp_88AB6;
	assign sv2v_tmp_88AB6 = op_mod_q;
	always @(*) mid_pipe_op_mod_q[0] = sv2v_tmp_88AB6;
	wire [3:1] sv2v_tmp_32E16;
	assign sv2v_tmp_32E16 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_32E16;
	wire [3:1] sv2v_tmp_DE9EA;
	assign sv2v_tmp_DE9EA = src_fmt_q;
	always @(*) mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_DE9EA;
	wire [3:1] sv2v_tmp_FC1E4;
	assign sv2v_tmp_FC1E4 = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_FC1E4;
	wire [2:1] sv2v_tmp_2AE08;
	assign sv2v_tmp_2AE08 = int_fmt_q;
	always @(*) mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] = sv2v_tmp_2AE08;
	wire [3:1] sv2v_tmp_BC8FE;
	assign sv2v_tmp_BC8FE = inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_tag_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_BC8FE;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_A8626;
	assign sv2v_tmp_A8626 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_A8626;
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			wire reg_ena;
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_input_sign_q[i + 1] <= 1'sb0;
				else
					mid_pipe_input_sign_q[i + 1] <= (reg_ena ? mid_pipe_input_sign_q[i] : mid_pipe_input_sign_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= 1'sb0;
				else
					mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH] <= (reg_ena ? mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_MAN_WIDTH+:INT_MAN_WIDTH] : mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_MAN_WIDTH+:INT_MAN_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH] <= (reg_ena ? mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * INT_EXP_WIDTH+:INT_EXP_WIDTH] : mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * INT_EXP_WIDTH+:INT_EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_src_is_int_q[i + 1] <= 1'sb0;
				else
					mid_pipe_src_is_int_q[i + 1] <= (reg_ena ? mid_pipe_src_is_int_q[i] : mid_pipe_src_is_int_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_dst_is_int_q[i + 1] <= 1'sb0;
				else
					mid_pipe_dst_is_int_q[i + 1] <= (reg_ena ? mid_pipe_dst_is_int_q[i] : mid_pipe_dst_is_int_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= 1'sb0;
				else
					mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8] <= (reg_ena ? mid_pipe_info_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 8+:8] : mid_pipe_info_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 8+:8]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_mant_zero_q[i + 1] <= 1'sb0;
				else
					mid_pipe_mant_zero_q[i + 1] <= (reg_ena ? mid_pipe_mant_zero_q[i] : mid_pipe_mant_zero_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					mid_pipe_op_mod_q[i + 1] <= (reg_ena ? mid_pipe_op_mod_q[i] : mid_pipe_op_mod_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= sv2v_cast_87CC5(0);
				else
					mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] <= (reg_ena ? mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS] : mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign input_sign_q = mid_pipe_input_sign_q[NUM_MID_REGS];
	assign input_exp_q = mid_pipe_input_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	assign input_mant_q = mid_pipe_input_mant_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_MAN_WIDTH+:INT_MAN_WIDTH];
	assign destination_exp_q = mid_pipe_dest_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * INT_EXP_WIDTH+:INT_EXP_WIDTH];
	assign src_is_int_q = mid_pipe_src_is_int_q[NUM_MID_REGS];
	assign dst_is_int_q = mid_pipe_dst_is_int_q[NUM_MID_REGS];
	assign info_q = mid_pipe_info_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 8+:8];
	assign mant_is_zero_q = mid_pipe_mant_zero_q[NUM_MID_REGS];
	assign op_mod_q2 = mid_pipe_op_mod_q[NUM_MID_REGS];
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	assign src_fmt_q2 = mid_pipe_src_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign int_fmt_q2 = mid_pipe_int_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_INT_FORMAT_BITS+:fpnew_pkg_INT_FORMAT_BITS];
	reg [INT_EXP_WIDTH - 1:0] final_exp;
	reg [2 * INT_MAN_WIDTH:0] preshift_mant;
	wire [2 * INT_MAN_WIDTH:0] destination_mant;
	wire [SUPER_MAN_BITS - 1:0] final_mant;
	wire [MAX_INT_WIDTH - 1:0] final_int;
	reg [$clog2(INT_MAN_WIDTH + 1) - 1:0] denorm_shamt;
	wire [1:0] fp_round_sticky_bits;
	wire [1:0] int_round_sticky_bits;
	wire [1:0] round_sticky_bits;
	reg of_before_round;
	reg uf_before_round;
	always @(*) begin : cast_value
		final_exp = $unsigned(destination_exp_q);
		preshift_mant = 1'sb0;
		denorm_shamt = SUPER_MAN_BITS - fpnew_pkg_man_bits(dst_fmt_q2);
		of_before_round = 1'b0;
		uf_before_round = 1'b0;
		preshift_mant = input_mant_q << (INT_MAN_WIDTH + 1);
		if (dst_is_int_q) begin
			denorm_shamt = $unsigned((MAX_INT_WIDTH - 1) - input_exp_q);
			if (input_exp_q >= $signed((fpnew_pkg_int_width(int_fmt_q2) - 1) + op_mod_q2)) begin
				denorm_shamt = 1'sb0;
				of_before_round = 1'b1;
			end
			else if (input_exp_q < -1) begin
				denorm_shamt = MAX_INT_WIDTH + 1;
				uf_before_round = 1'b1;
			end
		end
		else if ((destination_exp_q >= ($signed(2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1)) || (~src_is_int_q && info_q[4])) begin
			final_exp = $unsigned((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 2);
			preshift_mant = 1'sb1;
			of_before_round = 1'b1;
		end
		else if ((destination_exp_q < 1) && (destination_exp_q >= -$signed(fpnew_pkg_man_bits(dst_fmt_q2)))) begin
			final_exp = 1'sb0;
			denorm_shamt = $unsigned((denorm_shamt + 1) - destination_exp_q);
			uf_before_round = 1'b1;
		end
		else if (destination_exp_q < -$signed(fpnew_pkg_man_bits(dst_fmt_q2))) begin
			final_exp = 1'sb0;
			denorm_shamt = $unsigned((denorm_shamt + 2) + fpnew_pkg_man_bits(dst_fmt_q2));
			uf_before_round = 1'b1;
		end
	end
	localparam NUM_FP_STICKY = ((2 * INT_MAN_WIDTH) - SUPER_MAN_BITS) - 1;
	localparam NUM_INT_STICKY = (2 * INT_MAN_WIDTH) - MAX_INT_WIDTH;
	assign destination_mant = preshift_mant >> denorm_shamt;
	assign {final_mant, fp_round_sticky_bits[1]} = destination_mant[(2 * INT_MAN_WIDTH) - 1-:SUPER_MAN_BITS + 1];
	assign {final_int, int_round_sticky_bits[1]} = destination_mant[2 * INT_MAN_WIDTH-:MAX_INT_WIDTH + 1];
	assign fp_round_sticky_bits[0] = |{destination_mant[NUM_FP_STICKY - 1:0]};
	assign int_round_sticky_bits[0] = |{destination_mant[NUM_INT_STICKY - 1:0]};
	assign round_sticky_bits = (dst_is_int_q ? int_round_sticky_bits : fp_round_sticky_bits);
	wire [WIDTH - 1:0] pre_round_abs;
	wire of_after_round;
	wire uf_after_round;
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_pre_round_abs;
	reg [4:0] fmt_of_after_round;
	reg [4:0] fmt_uf_after_round;
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_pre_round_abs;
	wire rounded_sign;
	wire [WIDTH - 1:0] rounded_abs;
	wire result_true_zero;
	wire [WIDTH - 1:0] rounded_int_res;
	wire rounded_int_res_zero;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				always @(*) begin : assemble_result
					fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = {final_exp[EXP_BITS - 1:0], final_mant[MAN_BITS - 1:0]};
				end
			end
			else begin : inactive_format
				wire [WIDTH * 1:1] sv2v_tmp_C33E0;
				assign sv2v_tmp_C33E0 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_pre_round_abs[fmt * WIDTH+:WIDTH] = sv2v_tmp_C33E0;
			end
		end
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_int_res_sign_ext
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				always @(*) begin : assemble_result
					ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = {WIDTH {final_int[INT_WIDTH - 1]}};
					ifmt_pre_round_abs[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = final_int[INT_WIDTH - 1:0];
				end
			end
			else begin : inactive_format
				wire [WIDTH * 1:1] sv2v_tmp_F6FA8;
				assign sv2v_tmp_F6FA8 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_pre_round_abs[ifmt * WIDTH+:WIDTH] = sv2v_tmp_F6FA8;
			end
		end
	endgenerate
	assign pre_round_abs = (dst_is_int_q ? ifmt_pre_round_abs[int_fmt_q2 * WIDTH+:WIDTH] : fmt_pre_round_abs[dst_fmt_q2 * WIDTH+:WIDTH]);
	fpnew_rounding #(.AbsWidth(WIDTH)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(input_sign_q),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(1'b0),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_true_zero)
	);
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				always @(*) begin : post_process
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = (src_is_int_q & mant_is_zero_q ? {FP_WIDTH * 1 {1'sb0}} : {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]});
				end
			end
			else begin : inactive_format
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				wire [WIDTH * 1:1] sv2v_tmp_649FB;
				assign sv2v_tmp_649FB = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_649FB;
			end
		end
	endgenerate
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	assign rounded_int_res = (rounded_sign ? $unsigned(-rounded_abs) : rounded_abs);
	assign rounded_int_res_zero = rounded_int_res == {WIDTH {1'sb0}};
	wire [WIDTH - 1:0] fp_special_result;
	wire [4:0] fp_special_status;
	wire fp_result_is_special;
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			if (FpFmtConfig[fmt]) begin : active_format
				always @(*) begin : special_results
					reg [FP_WIDTH - 1:0] special_res;
					special_res = (info_q[5] ? input_sign_q << (FP_WIDTH - 1) : {1'b0, QNAN_EXPONENT, QNAN_MANTISSA});
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				wire [WIDTH * 1:1] sv2v_tmp_B718F;
				assign sv2v_tmp_B718F = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_B718F;
			end
		end
	endgenerate
	assign fp_result_is_special = ~src_is_int_q & ((info_q[5] | info_q[3]) | ~info_q[0]);
	assign fp_special_status = {info_q[2], 4'b0000};
	assign fp_special_result = fmt_special_result[dst_fmt_q2 * WIDTH+:WIDTH];
	wire [WIDTH - 1:0] int_special_result;
	wire [4:0] int_special_status;
	wire int_result_is_special;
	reg [(NUM_INT_FORMATS * WIDTH) - 1:0] ifmt_special_result;
	generate
		for (ifmt = 0; ifmt < sv2v_cast_32_signed(NUM_INT_FORMATS); ifmt = ifmt + 1) begin : gen_special_results_int
			localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
			if (IntFmtConfig[ifmt]) begin : active_format
				always @(*) begin : special_results
					reg [INT_WIDTH - 1:0] special_res;
					special_res[INT_WIDTH - 2:0] = 1'sb1;
					special_res[INT_WIDTH - 1] = op_mod_q2;
					if (input_sign_q && !info_q[3])
						special_res = ~special_res;
					ifmt_special_result[ifmt * WIDTH+:WIDTH] = {WIDTH {special_res[INT_WIDTH - 1]}};
					ifmt_special_result[(ifmt * WIDTH) + (INT_WIDTH - 1)-:INT_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				wire [WIDTH * 1:1] sv2v_tmp_99B6D;
				assign sv2v_tmp_99B6D = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) ifmt_special_result[ifmt * WIDTH+:WIDTH] = sv2v_tmp_99B6D;
			end
		end
	endgenerate
	assign int_result_is_special = (((info_q[3] | info_q[4]) | of_before_round) | ~info_q[0]) | ((input_sign_q & op_mod_q2) & ~rounded_int_res_zero);
	assign int_special_status = 5'b10000;
	assign int_special_result = ifmt_special_result[int_fmt_q2 * WIDTH+:WIDTH];
	wire [4:0] int_regular_status;
	wire [4:0] fp_regular_status;
	wire [WIDTH - 1:0] fp_result;
	wire [WIDTH - 1:0] int_result;
	wire [4:0] fp_status;
	wire [4:0] int_status;
	assign fp_regular_status[4] = src_is_int_q & (of_before_round | of_after_round);
	assign fp_regular_status[3] = 1'b0;
	assign fp_regular_status[2] = ~src_is_int_q & (~info_q[4] & (of_before_round | of_after_round));
	assign fp_regular_status[1] = uf_after_round & fp_regular_status[0];
	assign fp_regular_status[0] = (src_is_int_q ? |fp_round_sticky_bits : |fp_round_sticky_bits | (~info_q[4] & (of_before_round | of_after_round)));
	assign int_regular_status = {4'b0000, |int_round_sticky_bits};
	assign fp_result = (fp_result_is_special ? fp_special_result : fmt_result[dst_fmt_q2 * WIDTH+:WIDTH]);
	assign fp_status = (fp_result_is_special ? fp_special_status : fp_regular_status);
	assign int_result = (int_result_is_special ? int_special_result : rounded_int_res);
	assign int_status = (int_result_is_special ? int_special_status : int_regular_status);
	wire [WIDTH - 1:0] result_d;
	wire [4:0] status_d;
	wire extension_bit;
	assign result_d = (dst_is_int_q ? int_result : fp_result);
	assign status_d = (dst_is_int_q ? int_status : fp_status);
	assign extension_bit = (dst_is_int_q ? int_result[WIDTH - 1] : 1'b1);
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	reg [0:NUM_OUT_REGS] out_pipe_ext_bit_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 3) + ((NUM_OUT_REGS * 3) - 1) : ((NUM_OUT_REGS + 1) * 3) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 3 : 0)] out_pipe_tag_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	wire [WIDTH * 1:1] sv2v_tmp_4086F;
	assign sv2v_tmp_4086F = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_4086F;
	wire [5:1] sv2v_tmp_B7C45;
	assign sv2v_tmp_B7C45 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_B7C45;
	wire [1:1] sv2v_tmp_8F736;
	assign sv2v_tmp_8F736 = extension_bit;
	always @(*) out_pipe_ext_bit_q[0] = sv2v_tmp_8F736;
	wire [3:1] sv2v_tmp_1DCFD;
	assign sv2v_tmp_1DCFD = mid_pipe_tag_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 3+:3] = sv2v_tmp_1DCFD;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_3BE1D;
	assign sv2v_tmp_3BE1D = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_3BE1D;
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			wire reg_ena;
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_ext_bit_q[i + 1] <= 1'sb0;
				else
					out_pipe_ext_bit_q[i + 1] <= (reg_ena ? out_pipe_ext_bit_q[i] : out_pipe_ext_bit_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 3+:3] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	assign extension_bit_o = out_pipe_ext_bit_q[NUM_OUT_REGS];
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 3+:3];
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_classifier (
	operands_i,
	is_boxed_i,
	info_o
);
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	parameter [31:0] NumOperands = 1;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	input wire [(NumOperands * WIDTH) - 1:0] operands_i;
	input wire [NumOperands - 1:0] is_boxed_i;
	output reg [(NumOperands * 8) - 1:0] info_o;
	function automatic [31:0] fpnew_pkg_exp_bits;
		input reg [2:0] fmt;
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	function automatic [31:0] fpnew_pkg_man_bits;
		input reg [2:0] fmt;
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	genvar op;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (op = 0; op < sv2v_cast_32_signed(NumOperands); op = op + 1) begin : gen_num_values
			reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] value;
			reg is_boxed;
			reg is_normal;
			reg is_inf;
			reg is_nan;
			reg is_signalling;
			reg is_quiet;
			reg is_zero;
			reg is_subnormal;
			always @(*) begin : classify_input
				value = operands_i[op * WIDTH+:WIDTH];
				is_boxed = is_boxed_i[op];
				is_normal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] != {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}});
				is_zero = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}});
				is_subnormal = (is_boxed && (value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb0}})) && !is_zero;
				is_inf = is_boxed && ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] == {MAN_BITS * 1 {1'sb0}}));
				is_nan = !is_boxed || ((value[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)] == {((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1) * 1 {1'sb1}}) && (value[MAN_BITS - 1-:MAN_BITS] != {MAN_BITS * 1 {1'sb0}}));
				is_signalling = (is_boxed && is_nan) && (value[(MAN_BITS - 1) - ((MAN_BITS - 1) - (MAN_BITS - 1))] == 1'b0);
				is_quiet = is_nan && !is_signalling;
				info_o[(op * 8) + 7] = is_normal;
				info_o[(op * 8) + 6] = is_subnormal;
				info_o[(op * 8) + 5] = is_zero;
				info_o[(op * 8) + 4] = is_inf;
				info_o[(op * 8) + 3] = is_nan;
				info_o[(op * 8) + 2] = is_signalling;
				info_o[(op * 8) + 1] = is_quiet;
				info_o[op * 8] = is_boxed;
			end
		end
	endgenerate
endmodule
module fpnew_divsqrt_multi_C04AD_31CA4 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [31:0] AuxType_AUX_BITS = 0;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	parameter [0:4] FpFmtConfig = 1'sb1;
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd1;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	input wire clk_i;
	input wire rst_ni;
	input wire [(2 * WIDTH) - 1:0] operands_i;
	input wire [9:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire [2:0] dst_fmt_i;
	input wire [2:0] tag_i;
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	localparam NUM_OUT_REGS = ((PipeConfig == 2'd1) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	wire [(2 * WIDTH) - 1:0] operands_q;
	wire [2:0] rnd_mode_q;
	wire [3:0] op_q;
	wire [2:0] dst_fmt_q;
	wire in_valid_q;
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_tag_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	wire [2 * WIDTH:1] sv2v_tmp_83757;
	assign sv2v_tmp_83757 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_83757;
	wire [3:1] sv2v_tmp_857E9;
	assign sv2v_tmp_857E9 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_857E9;
	wire [4:1] sv2v_tmp_4BFFB;
	assign sv2v_tmp_4BFFB = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_4BFFB;
	wire [3:1] sv2v_tmp_54055;
	assign sv2v_tmp_54055 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_54055;
	wire [3:1] sv2v_tmp_0DF27;
	assign sv2v_tmp_0DF27 = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_0DF27;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_CDB25;
	assign sv2v_tmp_CDB25 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_CDB25;
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	assign in_ready_o = inp_pipe_ready[0];
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			wire reg_ena;
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2];
	assign rnd_mode_q = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	assign op_q = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS];
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign in_valid_q = inp_pipe_valid_q[NUM_INP_REGS];
	reg [1:0] divsqrt_fmt;
	reg [127:0] divsqrt_operands;
	reg input_is_fp8;
	always @(*) begin : translate_fmt
		case (dst_fmt_q)
			sv2v_cast_0BC43('d0): divsqrt_fmt = 2'b00;
			sv2v_cast_0BC43('d1): divsqrt_fmt = 2'b01;
			sv2v_cast_0BC43('d2): divsqrt_fmt = 2'b10;
			sv2v_cast_0BC43('d4): divsqrt_fmt = 2'b11;
			default: divsqrt_fmt = 2'b10;
		endcase
		input_is_fp8 = FpFmtConfig[sv2v_cast_0BC43('d3)] & (dst_fmt_q == sv2v_cast_0BC43('d3));
		divsqrt_operands[0+:64] = (input_is_fp8 ? operands_q[0+:WIDTH] << 8 : operands_q[0+:WIDTH]);
		divsqrt_operands[64+:64] = (input_is_fp8 ? operands_q[WIDTH+:WIDTH] << 8 : operands_q[WIDTH+:WIDTH]);
	end
	reg in_ready;
	wire div_valid;
	wire sqrt_valid;
	wire unit_ready;
	wire unit_done;
	wire op_starting;
	reg out_valid;
	wire out_ready;
	reg hold_result;
	reg data_is_held;
	reg unit_busy;
	reg [1:0] state_q;
	reg [1:0] state_d;
	assign inp_pipe_ready[NUM_INP_REGS] = in_ready;
	assign div_valid = ((in_valid_q & (op_q == sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	assign sqrt_valid = ((in_valid_q & (op_q != sv2v_cast_A53F3(4))) & in_ready) & ~flush_i;
	assign op_starting = div_valid | sqrt_valid;
	always @(*) begin : flag_fsm
		in_ready = 1'b0;
		out_valid = 1'b0;
		hold_result = 1'b0;
		data_is_held = 1'b0;
		unit_busy = 1'b0;
		state_d = state_q;
		case (state_q)
			2'd0: begin
				in_ready = 1'b1;
				if (in_valid_q && unit_ready)
					state_d = 2'd1;
			end
			2'd1: begin
				unit_busy = 1'b1;
				if (unit_done) begin
					out_valid = 1'b1;
					if (out_ready) begin
						state_d = 2'd0;
						if (in_valid_q && unit_ready) begin
							in_ready = 1'b1;
							state_d = 2'd1;
						end
					end
					else begin
						hold_result = 1'b1;
						state_d = 2'd2;
					end
				end
			end
			2'd2: begin
				unit_busy = 1'b1;
				data_is_held = 1'b1;
				out_valid = 1'b1;
				if (out_ready) begin
					state_d = 2'd0;
					if (in_valid_q && unit_ready) begin
						in_ready = 1'b1;
						state_d = 2'd1;
					end
				end
			end
			default: state_d = 2'd0;
		endcase
		if (flush_i) begin
			unit_busy = 1'b0;
			out_valid = 1'b0;
			state_d = 2'd0;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			state_q <= 2'd0;
		else
			state_q <= state_d;
	reg result_is_fp8_q;
	reg [2:0] result_tag_q;
	reg [AuxType_AUX_BITS - 1:0] result_aux_q;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			result_is_fp8_q <= 1'sb0;
		else
			result_is_fp8_q <= (op_starting ? input_is_fp8 : result_is_fp8_q);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			result_tag_q <= 1'sb0;
		else
			result_tag_q <= (op_starting ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3] : result_tag_q);
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni)
			result_aux_q <= 1'sb0;
		else
			result_aux_q <= (op_starting ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : result_aux_q);
	wire [63:0] unit_result;
	wire [WIDTH - 1:0] adjusted_result;
	reg [WIDTH - 1:0] held_result_q;
	wire [4:0] unit_status;
	reg [4:0] held_status_q;
	localparam [5:0] sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0 = 1'sb0;
	div_sqrt_top_mvp i_divsqrt_lei(
		.Clk_CI(clk_i),
		.Rst_RBI(rst_ni),
		.Div_start_SI(div_valid),
		.Sqrt_start_SI(sqrt_valid),
		.Operand_a_DI(divsqrt_operands[0+:64]),
		.Operand_b_DI(divsqrt_operands[64+:64]),
		.RM_SI(rnd_mode_q),
		.Precision_ctl_SI(sv2v_uu_i_divsqrt_lei_ext_Precision_ctl_SI_0),
		.Format_sel_SI(divsqrt_fmt),
		.Kill_SI(flush_i),
		.Result_DO(unit_result),
		.Fflags_SO(unit_status),
		.Ready_SO(unit_ready),
		.Done_SO(unit_done)
	);
	assign adjusted_result = (result_is_fp8_q ? unit_result >> 8 : unit_result);
	always @(posedge clk_i) held_result_q <= (hold_result ? adjusted_result : held_result_q);
	always @(posedge clk_i) held_status_q <= (hold_result ? unit_status : held_status_q);
	wire [WIDTH - 1:0] result_d;
	wire [4:0] status_d;
	assign result_d = (data_is_held ? held_result_q : adjusted_result);
	assign status_d = (data_is_held ? held_status_q : unit_status);
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 3) + ((NUM_OUT_REGS * 3) - 1) : ((NUM_OUT_REGS + 1) * 3) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 3 : 0)] out_pipe_tag_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	wire [WIDTH * 1:1] sv2v_tmp_6C30D;
	assign sv2v_tmp_6C30D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_6C30D;
	wire [5:1] sv2v_tmp_2ED07;
	assign sv2v_tmp_2ED07 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2ED07;
	wire [3:1] sv2v_tmp_77C11;
	assign sv2v_tmp_77C11 = result_tag_q;
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 3+:3] = sv2v_tmp_77C11;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_7E003;
	assign sv2v_tmp_7E003 = result_aux_q;
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_7E003;
	wire [1:1] sv2v_tmp_D06FD;
	assign sv2v_tmp_D06FD = out_valid;
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_D06FD;
	assign out_ready = out_pipe_ready[0];
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			wire reg_ena;
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 3+:3] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	assign extension_bit_o = 1'b1;
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 3+:3];
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	assign busy_o = |{inp_pipe_valid_q, unit_busy, out_pipe_valid_q};
endmodule
module fpnew_fma_multi_FF0B0_361DB (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [31:0] AuxType_AUX_BITS = 0;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	parameter [0:4] FpFmtConfig = 1'sb1;
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	input wire clk_i;
	input wire rst_ni;
	input wire [(3 * WIDTH) - 1:0] operands_i;
	input wire [14:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	input wire [2:0] src_fmt_i;
	input wire [2:0] dst_fmt_i;
	input wire [2:0] tag_i;
	input wire [AuxType_AUX_BITS - 1:0] aux_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire [AuxType_AUX_BITS - 1:0] aux_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	function automatic [31:0] fpnew_pkg_exp_bits;
		input reg [2:0] fmt;
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	function automatic [31:0] fpnew_pkg_man_bits;
		input reg [2:0] fmt;
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	function automatic [63:0] fpnew_pkg_super_format;
		input reg [0:4] cfg;
		reg [63:0] res;
		begin
			res = 1'sb0;
			begin : sv2v_autoblock_2
				reg [31:0] fmt;
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					if (cfg[fmt]) begin
						res[63-:32] = $unsigned(fpnew_pkg_maximum(res[63-:32], fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt))));
						res[31-:32] = $unsigned(fpnew_pkg_maximum(res[31-:32], fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt))));
					end
			end
			fpnew_pkg_super_format = res;
		end
	endfunction
	localparam [63:0] SUPER_FORMAT = fpnew_pkg_super_format(FpFmtConfig);
	localparam [31:0] SUPER_EXP_BITS = SUPER_FORMAT[63-:32];
	localparam [31:0] SUPER_MAN_BITS = SUPER_FORMAT[31-:32];
	localparam [31:0] PRECISION_BITS = SUPER_MAN_BITS + 1;
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	localparam [31:0] EXP_WIDTH = fpnew_pkg_maximum(SUPER_EXP_BITS + 2, LZC_RESULT_WIDTH);
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	wire [(3 * WIDTH) - 1:0] operands_q;
	wire [2:0] src_fmt_q;
	wire [2:0] dst_fmt_q;
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0)) + 1) * 3) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)) + 1) * 3) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) * 3 : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) * 3)] inp_pipe_is_boxed_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_src_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] inp_pipe_dst_fmt_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_tag_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * AuxType_AUX_BITS) + ((NUM_INP_REGS * AuxType_AUX_BITS) - 1) : ((NUM_INP_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * AuxType_AUX_BITS : 0)] inp_pipe_aux_q;
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	wire [3 * WIDTH:1] sv2v_tmp_5DCC9;
	assign sv2v_tmp_5DCC9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_5DCC9;
	wire [15:1] sv2v_tmp_7F60B;
	assign sv2v_tmp_7F60B = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] = sv2v_tmp_7F60B;
	wire [3:1] sv2v_tmp_700C1;
	assign sv2v_tmp_700C1 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_700C1;
	wire [4:1] sv2v_tmp_3923B;
	assign sv2v_tmp_3923B = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_3923B;
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	wire [3:1] sv2v_tmp_6B115;
	assign sv2v_tmp_6B115 = src_fmt_i;
	always @(*) inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_6B115;
	wire [3:1] sv2v_tmp_B8677;
	assign sv2v_tmp_B8677 = dst_fmt_i;
	always @(*) inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_B8677;
	wire [3:1] sv2v_tmp_8D5DD;
	assign sv2v_tmp_8D5DD = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_8D5DD;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_08A77;
	assign sv2v_tmp_08A77 = aux_i;
	always @(*) inp_pipe_aux_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_08A77;
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	assign in_ready_o = inp_pipe_ready[0];
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [AuxType_AUX_BITS - 1:0] sv2v_cast_14358;
		input reg [AuxType_AUX_BITS - 1:0] inp;
		sv2v_cast_14358 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			wire reg_ena;
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= 1'sb0;
				else
					inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] <= (reg_ena ? inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15] : inp_pipe_is_boxed_q[3 * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * NUM_FORMATS) + 4) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1)))+:15]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : inp_pipe_aux_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign operands_q = inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3];
	assign src_fmt_q = inp_pipe_src_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign dst_fmt_q = inp_pipe_dst_fmt_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	wire [14:0] fmt_sign;
	wire signed [(15 * SUPER_EXP_BITS) - 1:0] fmt_exponent;
	wire [(15 * SUPER_MAN_BITS) - 1:0] fmt_mantissa;
	wire [119:0] info_q;
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic signed [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6_signed;
		input reg signed [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6_signed = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_52F63;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_52F63 = inp;
	endfunction
	function automatic [7:0] sv2v_cast_8;
		input reg [7:0] inp;
		sv2v_cast_8 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : fmt_init_inputs
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				wire [(3 * FP_WIDTH) - 1:0] trimmed_ops;
				fpnew_classifier #(
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.NumOperands(3)
				) i_fpnew_classifier(
					.operands_i(trimmed_ops),
					.is_boxed_i(inp_pipe_is_boxed_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt : (0 >= NUM_INP_REGS ? NUM_INP_REGS * NUM_FORMATS : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * NUM_FORMATS) + fmt) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * NUM_FORMATS) + ((NUM_INP_REGS * NUM_FORMATS) - 1) : ((NUM_INP_REGS + 1) * NUM_FORMATS) - 1))) * 3+:3]),
					.info_o(info_q[8 * (fmt * 3)+:24])
				);
				genvar op;
				for (op = 0; op < 3; op = op + 1) begin : gen_operands
					assign trimmed_ops[op * fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))+:fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH];
					assign fmt_sign[(fmt * 3) + op] = operands_q[(op * WIDTH) + (FP_WIDTH - 1)];
					assign fmt_exponent[((fmt * 3) + op) * SUPER_EXP_BITS+:SUPER_EXP_BITS] = $signed({1'b0, operands_q[(op * WIDTH) + MAN_BITS+:EXP_BITS]});
					assign fmt_mantissa[((fmt * 3) + op) * SUPER_MAN_BITS+:SUPER_MAN_BITS] = {info_q[(((fmt * 3) + op) * 8) + 7], operands_q[(op * WIDTH) + (MAN_BITS - 1)-:MAN_BITS]} << (SUPER_MAN_BITS - MAN_BITS);
				end
			end
			else begin : inactive_format
				assign info_q[8 * (fmt * 3)+:24] = {3 {sv2v_cast_8(fpnew_pkg_DONT_CARE)}};
				assign fmt_sign[fmt * 3+:3] = fpnew_pkg_DONT_CARE;
				assign fmt_exponent[SUPER_EXP_BITS * (fmt * 3)+:SUPER_EXP_BITS * 3] = {3 {sv2v_cast_A3BB6_signed(fpnew_pkg_DONT_CARE)}};
				assign fmt_mantissa[SUPER_MAN_BITS * (fmt * 3)+:SUPER_MAN_BITS * 3] = {3 {sv2v_cast_52F63(fpnew_pkg_DONT_CARE)}};
			end
		end
	endgenerate
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_a;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_b;
	reg [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] operand_c;
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	function automatic [31:0] fpnew_pkg_bias;
		input reg [2:0] fmt;
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_A3BB6;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_A3BB6 = inp;
	endfunction
	function automatic [SUPER_MAN_BITS - 1:0] sv2v_cast_FC661;
		input reg [SUPER_MAN_BITS - 1:0] inp;
		sv2v_cast_FC661 = inp;
	endfunction
	function automatic [SUPER_EXP_BITS - 1:0] sv2v_cast_705CC;
		input reg [SUPER_EXP_BITS - 1:0] inp;
		sv2v_cast_705CC = inp;
	endfunction
	always @(*) begin : op_select
		operand_a = {fmt_sign[src_fmt_q * 3], fmt_exponent[(src_fmt_q * 3) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[(src_fmt_q * 3) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		operand_b = {fmt_sign[(src_fmt_q * 3) + 1], fmt_exponent[((src_fmt_q * 3) + 1) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((src_fmt_q * 3) + 1) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		operand_c = {fmt_sign[(dst_fmt_q * 3) + 2], fmt_exponent[((dst_fmt_q * 3) + 2) * SUPER_EXP_BITS+:SUPER_EXP_BITS], fmt_mantissa[((dst_fmt_q * 3) + 2) * SUPER_MAN_BITS+:SUPER_MAN_BITS]};
		info_a = info_q[(src_fmt_q * 3) * 8+:8];
		info_b = info_q[((src_fmt_q * 3) + 1) * 8+:8];
		info_c = info_q[((dst_fmt_q * 3) + 2) * 8+:8];
		operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1): operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] = ~operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				operand_a = {1'b0, sv2v_cast_A3BB6(fpnew_pkg_bias(src_fmt_q)), sv2v_cast_FC661(1'sb0)};
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				operand_c = {1'b1, sv2v_cast_705CC(1'sb0), sv2v_cast_FC661(1'sb0)};
				info_c = 8'b00100001;
			end
			default: begin
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_A3BB6(fpnew_pkg_DONT_CARE), sv2v_cast_52F63(fpnew_pkg_DONT_CARE)};
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	wire any_operand_inf;
	wire any_operand_nan;
	wire signalling_nan;
	wire effective_subtraction;
	wire tentative_sign;
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	assign effective_subtraction = (operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))]) ^ operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	assign tentative_sign = operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))];
	wire [WIDTH - 1:0] special_result;
	wire [4:0] special_status;
	wire result_is_special;
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_special_result;
	reg [24:0] fmt_special_status;
	reg [4:0] fmt_result_is_special;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_special_results
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			localparam [EXP_BITS - 1:0] QNAN_EXPONENT = 1'sb1;
			localparam [MAN_BITS - 1:0] QNAN_MANTISSA = 2 ** (MAN_BITS - 1);
			localparam [MAN_BITS - 1:0] ZERO_MANTISSA = 1'sb0;
			if (FpFmtConfig[fmt]) begin : active_format
				always @(*) begin : special_results
					reg [FP_WIDTH - 1:0] special_res;
					special_res = {1'b0, QNAN_EXPONENT, QNAN_MANTISSA};
					fmt_special_status[fmt * 5+:5] = 1'sb0;
					fmt_result_is_special[fmt] = 1'b0;
					if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
						fmt_result_is_special[fmt] = 1'b1;
						fmt_special_status[(fmt * 5) + 4] = 1'b1;
					end
					else if (any_operand_nan) begin
						fmt_result_is_special[fmt] = 1'b1;
						fmt_special_status[(fmt * 5) + 4] = signalling_nan;
					end
					else if (any_operand_inf) begin
						fmt_result_is_special[fmt] = 1'b1;
						if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
							fmt_special_status[(fmt * 5) + 4] = 1'b1;
						else if (info_a[4] || info_b[4])
							special_res = {operand_a[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))] ^ operand_b[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
						else if (info_c[4])
							special_res = {operand_c[1 + (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))], QNAN_EXPONENT, ZERO_MANTISSA};
					end
					fmt_special_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					fmt_special_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = special_res;
				end
			end
			else begin : inactive_format
				wire [WIDTH * 1:1] sv2v_tmp_7740B;
				assign sv2v_tmp_7740B = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_special_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_7740B;
			end
		end
	endgenerate
	assign result_is_special = fmt_result_is_special[dst_fmt_q];
	assign special_status = fmt_special_status[dst_fmt_q * 5+:5];
	assign special_result = fmt_special_result[dst_fmt_q * WIDTH+:WIDTH];
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	assign exponent_a = $signed({1'b0, operand_a[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	assign exponent_b = $signed({1'b0, operand_b[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	assign exponent_c = $signed({1'b0, operand_c[SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)-:((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) >= (SUPER_MAN_BITS + 0) ? ((SUPER_EXP_BITS + (SUPER_MAN_BITS - 1)) - (SUPER_MAN_BITS + 0)) + 1 : ((SUPER_MAN_BITS + 0) - (SUPER_EXP_BITS + (SUPER_MAN_BITS - 1))) + 1)]});
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(fpnew_pkg_bias(dst_fmt_q)) : $signed(((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - (2 * $signed(fpnew_pkg_bias(src_fmt_q)))) + $signed(fpnew_pkg_bias(dst_fmt_q))));
	assign exponent_difference = exponent_addend - exponent_product;
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	always @(*) begin : addend_shift_amount
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			addend_shamt = 0;
	end
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	wire [(2 * PRECISION_BITS) - 1:0] product;
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	assign mantissa_a = {info_a[7], operand_a[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	assign mantissa_b = {info_b[7], operand_b[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	assign mantissa_c = {info_c[7], operand_c[SUPER_MAN_BITS - 1-:SUPER_MAN_BITS]};
	assign product = mantissa_a * mantissa_b;
	assign product_shifted = product << 2;
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	wire sticky_before_add;
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	wire inject_carry_in;
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	assign sticky_before_add = |addend_sticky_bits;
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	wire sum_carry;
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	wire final_sign;
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	wire effective_subtraction_q;
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	wire sticky_before_add_q;
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	wire final_sign_q;
	wire [2:0] dst_fmt_q2;
	wire [2:0] rnd_mode_q;
	wire result_is_special_q;
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) - 1:0] special_result_q;
	wire [4:0] special_status_q;
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS) + ((NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS) - 1) : ((NUM_MID_REGS + 1) * fpnew_pkg_FP_FORMAT_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * fpnew_pkg_FP_FORMAT_BITS : 0)] mid_pipe_dst_fmt_q;
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) + ((NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) : 0)] mid_pipe_spec_res_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_tag_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * AuxType_AUX_BITS) + ((NUM_MID_REGS * AuxType_AUX_BITS) - 1) : ((NUM_MID_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * AuxType_AUX_BITS : 0)] mid_pipe_aux_q;
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_8565A;
	assign sv2v_tmp_8565A = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_8565A;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_F1167;
	assign sv2v_tmp_F1167 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_F1167;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_19629;
	assign sv2v_tmp_19629 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_19629;
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_037F4;
	assign sv2v_tmp_037F4 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_037F4;
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_74CB3;
	assign sv2v_tmp_74CB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_74CB3;
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	wire [3:1] sv2v_tmp_2170E;
	assign sv2v_tmp_2170E = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_2170E;
	wire [3:1] sv2v_tmp_8A4AE;
	assign sv2v_tmp_8A4AE = dst_fmt_q;
	always @(*) mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] = sv2v_tmp_8A4AE;
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	wire [((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS) * 1:1] sv2v_tmp_1ADE6;
	assign sv2v_tmp_1ADE6 = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] = sv2v_tmp_1ADE6;
	wire [5:1] sv2v_tmp_1A1E3;
	assign sv2v_tmp_1A1E3 = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_1A1E3;
	wire [3:1] sv2v_tmp_D1C94;
	assign sv2v_tmp_D1C94 = inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_tag_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_D1C94;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_89EE4;
	assign sv2v_tmp_89EE4 = inp_pipe_aux_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) mid_pipe_aux_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_89EE4;
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			wire reg_ena;
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= sv2v_cast_0BC43(0);
				else
					mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] <= (reg_ena ? mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS] : mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= 1'sb0;
				else
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : mid_pipe_aux_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	assign dst_fmt_q2 = mid_pipe_dst_fmt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * fpnew_pkg_FP_FORMAT_BITS+:fpnew_pkg_FP_FORMAT_BITS];
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + SUPER_EXP_BITS) + SUPER_MAN_BITS)+:(1 + SUPER_EXP_BITS) + SUPER_MAN_BITS];
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	wire lzc_zeroes;
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	reg [PRECISION_BITS:0] final_mantissa;
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	wire sticky_after_norm;
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	always @(*) begin : norm_shift_amount
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
				norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
				normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
			end
			else begin
				norm_shamt = $unsigned($signed((PRECISION_BITS + 2) + exponent_product_q));
				normalized_exponent = 0;
			end
		end
		else begin
			norm_shamt = addend_shamt_q;
			normalized_exponent = tentative_exponent_q;
		end
	end
	assign sum_shifted = sum_q << norm_shamt;
	always @(*) begin : small_norm
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		final_exponent = normalized_exponent;
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			final_exponent = normalized_exponent - 1;
		end
		else
			final_exponent = 1'sb0;
	end
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	wire pre_round_sign;
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] pre_round_abs;
	wire [1:0] round_sticky_bits;
	wire of_before_round;
	wire of_after_round;
	wire uf_before_round;
	wire uf_after_round;
	wire [(NUM_FORMATS * (SUPER_EXP_BITS + SUPER_MAN_BITS)) - 1:0] fmt_pre_round_abs;
	wire [9:0] fmt_round_sticky_bits;
	reg [4:0] fmt_of_after_round;
	reg [4:0] fmt_uf_after_round;
	wire rounded_sign;
	wire [(SUPER_EXP_BITS + SUPER_MAN_BITS) - 1:0] rounded_abs;
	wire result_zero;
	assign of_before_round = final_exponent >= ((2 ** fpnew_pkg_exp_bits(dst_fmt_q2)) - 1);
	assign uf_before_round = final_exponent == 0;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_res_assemble
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			wire [EXP_BITS - 1:0] pre_round_exponent;
			wire [MAN_BITS - 1:0] pre_round_mantissa;
			if (FpFmtConfig[fmt]) begin : active_format
				assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : final_exponent[EXP_BITS - 1:0]);
				assign pre_round_mantissa = (of_before_round ? {fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt)) {1'sb1}} : final_mantissa[SUPER_MAN_BITS-:MAN_BITS]);
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {pre_round_exponent, pre_round_mantissa};
				assign fmt_round_sticky_bits[(fmt * 2) + 1] = final_mantissa[SUPER_MAN_BITS - MAN_BITS] | of_before_round;
				if (MAN_BITS < SUPER_MAN_BITS) begin : narrow_sticky
					assign fmt_round_sticky_bits[fmt * 2] = (|final_mantissa[(SUPER_MAN_BITS - MAN_BITS) - 1:0] | sticky_after_norm) | of_before_round;
				end
				else begin : normal_sticky
					assign fmt_round_sticky_bits[fmt * 2] = sticky_after_norm | of_before_round;
				end
			end
			else begin : inactive_format
				assign fmt_pre_round_abs[fmt * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS] = {SUPER_EXP_BITS + SUPER_MAN_BITS {fpnew_pkg_DONT_CARE}};
				assign fmt_round_sticky_bits[fmt * 2+:2] = {2 {fpnew_pkg_DONT_CARE}};
			end
		end
	endgenerate
	assign pre_round_sign = final_sign_q;
	assign pre_round_abs = fmt_pre_round_abs[dst_fmt_q2 * (SUPER_EXP_BITS + SUPER_MAN_BITS)+:SUPER_EXP_BITS + SUPER_MAN_BITS];
	assign round_sticky_bits = fmt_round_sticky_bits[dst_fmt_q2 * 2+:2];
	fpnew_rounding #(.AbsWidth(SUPER_EXP_BITS + SUPER_MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	reg [(NUM_FORMATS * WIDTH) - 1:0] fmt_result;
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_sign_inject
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(sv2v_cast_0BC43(fmt));
			localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(sv2v_cast_0BC43(fmt));
			if (FpFmtConfig[fmt]) begin : active_format
				always @(*) begin : post_process
					fmt_uf_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
					fmt_of_after_round[fmt] = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
					fmt_result[fmt * WIDTH+:WIDTH] = 1'sb1;
					fmt_result[(fmt * WIDTH) + (FP_WIDTH - 1)-:FP_WIDTH] = {rounded_sign, rounded_abs[(EXP_BITS + MAN_BITS) - 1:0]};
				end
			end
			else begin : inactive_format
				wire [1:1] sv2v_tmp_4A747;
				assign sv2v_tmp_4A747 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_uf_after_round[fmt] = sv2v_tmp_4A747;
				wire [1:1] sv2v_tmp_90681;
				assign sv2v_tmp_90681 = fpnew_pkg_DONT_CARE;
				always @(*) fmt_of_after_round[fmt] = sv2v_tmp_90681;
				wire [WIDTH * 1:1] sv2v_tmp_143A7;
				assign sv2v_tmp_143A7 = {WIDTH {fpnew_pkg_DONT_CARE}};
				always @(*) fmt_result[fmt * WIDTH+:WIDTH] = sv2v_tmp_143A7;
			end
		end
	endgenerate
	assign uf_after_round = fmt_uf_after_round[dst_fmt_q2];
	assign of_after_round = fmt_of_after_round[dst_fmt_q2];
	wire [WIDTH - 1:0] regular_result;
	wire [4:0] regular_status;
	assign regular_result = fmt_result[dst_fmt_q2 * WIDTH+:WIDTH];
	assign regular_status[4] = 1'b0;
	assign regular_status[3] = 1'b0;
	assign regular_status[2] = of_before_round | of_after_round;
	assign regular_status[1] = uf_after_round & regular_status[0];
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	wire [WIDTH - 1:0] result_d;
	wire [4:0] status_d;
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * WIDTH) + ((NUM_OUT_REGS * WIDTH) - 1) : ((NUM_OUT_REGS + 1) * WIDTH) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * WIDTH : 0)] out_pipe_result_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 3) + ((NUM_OUT_REGS * 3) - 1) : ((NUM_OUT_REGS + 1) * 3) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 3 : 0)] out_pipe_tag_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * AuxType_AUX_BITS) + ((NUM_OUT_REGS * AuxType_AUX_BITS) - 1) : ((NUM_OUT_REGS + 1) * AuxType_AUX_BITS) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * AuxType_AUX_BITS : 0)] out_pipe_aux_q;
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	wire [WIDTH * 1:1] sv2v_tmp_1212D;
	assign sv2v_tmp_1212D = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * WIDTH+:WIDTH] = sv2v_tmp_1212D;
	wire [5:1] sv2v_tmp_F691B;
	assign sv2v_tmp_F691B = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_F691B;
	wire [3:1] sv2v_tmp_AE3D3;
	assign sv2v_tmp_AE3D3 = mid_pipe_tag_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 3+:3] = sv2v_tmp_AE3D3;
	wire [AuxType_AUX_BITS * 1:1] sv2v_tmp_44007;
	assign sv2v_tmp_44007 = mid_pipe_aux_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	always @(*) out_pipe_aux_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS] = sv2v_tmp_44007;
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			wire reg_ena;
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= 1'sb0;
				else
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * WIDTH+:WIDTH] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * WIDTH+:WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 3+:3] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= sv2v_cast_14358(1'sb0);
				else
					out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS] <= (reg_ena ? out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * AuxType_AUX_BITS+:AuxType_AUX_BITS] : out_pipe_aux_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * AuxType_AUX_BITS+:AuxType_AUX_BITS]);
		end
	endgenerate
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * WIDTH+:WIDTH];
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	assign extension_bit_o = 1'b1;
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 3+:3];
	assign aux_o = out_pipe_aux_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * AuxType_AUX_BITS+:AuxType_AUX_BITS];
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_fma_F8EAE (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	input wire clk_i;
	input wire rst_ni;
	input wire [(3 * WIDTH) - 1:0] operands_i;
	input wire [2:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	input wire [2:0] tag_i;
	input wire aux_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire aux_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	function automatic [31:0] fpnew_pkg_exp_bits;
		input reg [2:0] fmt;
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	function automatic [31:0] fpnew_pkg_man_bits;
		input reg [2:0] fmt;
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	function automatic [31:0] fpnew_pkg_bias;
		input reg [2:0] fmt;
		fpnew_pkg_bias = $unsigned((2 ** (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] - 1)) - 1);
	endfunction
	localparam [31:0] BIAS = fpnew_pkg_bias(FpFormat);
	localparam [31:0] PRECISION_BITS = MAN_BITS + 1;
	localparam [31:0] LOWER_SUM_WIDTH = (2 * PRECISION_BITS) + 3;
	localparam [31:0] LZC_RESULT_WIDTH = $clog2(LOWER_SUM_WIDTH);
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	localparam [31:0] EXP_WIDTH = $unsigned(fpnew_pkg_maximum(EXP_BITS + 2, LZC_RESULT_WIDTH));
	localparam [31:0] SHIFT_AMOUNT_WIDTH = $clog2((3 * PRECISION_BITS) + 3);
	localparam NUM_INP_REGS = (PipeConfig == 2'd0 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 3 : 0));
	localparam NUM_MID_REGS = (PipeConfig == 2'd2 ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 2) / 3 : 0));
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 3 : 0));
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) * WIDTH)] inp_pipe_operands_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_is_boxed_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_tag_q;
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	wire [3 * WIDTH:1] sv2v_tmp_BC8B9;
	assign sv2v_tmp_BC8B9 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] = sv2v_tmp_BC8B9;
	wire [3:1] sv2v_tmp_FE389;
	assign sv2v_tmp_FE389 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_FE389;
	wire [3:1] sv2v_tmp_E1339;
	assign sv2v_tmp_E1339 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_E1339;
	wire [4:1] sv2v_tmp_CBA8F;
	assign sv2v_tmp_CBA8F = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_CBA8F;
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	wire [3:1] sv2v_tmp_31E69;
	assign sv2v_tmp_31E69 = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_31E69;
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	assign in_ready_o = inp_pipe_ready[0];
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			wire reg_ena;
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= 1'sb0;
				else
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 1'sb0;
				else
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	wire [23:0] info_q;
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(3)
	) i_class_inputs(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1)))+:WIDTH * 3]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3]),
		.info_o(info_q)
	);
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_c;
	reg [7:0] info_a;
	reg [7:0] info_b;
	reg [7:0] info_c;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_60B87;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_60B87 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_F33EE;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F33EE = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	always @(*) begin : op_select
		operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		operand_c = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3) + 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1))) * WIDTH+:WIDTH];
		info_a = info_q[0+:8];
		info_b = info_q[8+:8];
		info_c = info_q[16+:8];
		operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] = operand_c[1 + (EXP_BITS + (MAN_BITS - 1))] ^ inp_pipe_op_mod_q[NUM_INP_REGS];
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(0):
				;
			sv2v_cast_A53F3(1): operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] = ~operand_a[1 + (EXP_BITS + (MAN_BITS - 1))];
			sv2v_cast_A53F3(2): begin
				operand_a = {1'b0, sv2v_cast_91364(BIAS), sv2v_cast_60B87(1'sb0)};
				info_a = 8'b10000001;
			end
			sv2v_cast_A53F3(3): begin
				operand_c = {1'b1, sv2v_cast_F33EE(1'sb0), sv2v_cast_60B87(1'sb0)};
				info_c = 8'b00100001;
			end
			default: begin
				operand_a = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				operand_b = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				operand_c = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				info_a = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				info_b = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				info_c = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
			end
		endcase
	end
	wire any_operand_inf;
	wire any_operand_nan;
	wire signalling_nan;
	wire effective_subtraction;
	wire tentative_sign;
	assign any_operand_inf = |{info_a[4], info_b[4], info_c[4]};
	assign any_operand_nan = |{info_a[3], info_b[3], info_c[3]};
	assign signalling_nan = |{info_a[2], info_b[2], info_c[2]};
	assign effective_subtraction = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]) ^ operand_c[1 + (EXP_BITS + (MAN_BITS - 1))];
	assign tentative_sign = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))];
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result;
	reg [4:0] special_status;
	reg result_is_special;
	always @(*) begin : special_cases
		special_result = {1'b0, sv2v_cast_F33EE(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		special_status = 1'sb0;
		result_is_special = 1'b0;
		if ((info_a[4] && info_b[5]) || (info_a[5] && info_b[4])) begin
			result_is_special = 1'b1;
			special_status[4] = 1'b1;
		end
		else if (any_operand_nan) begin
			result_is_special = 1'b1;
			special_status[4] = signalling_nan;
		end
		else if (any_operand_inf) begin
			result_is_special = 1'b1;
			if (((info_a[4] || info_b[4]) && info_c[4]) && effective_subtraction)
				special_status[4] = 1'b1;
			else if (info_a[4] || info_b[4])
				special_result = {operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ^ operand_b[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
			else if (info_c[4])
				special_result = {operand_c[1 + (EXP_BITS + (MAN_BITS - 1))], sv2v_cast_F33EE(1'sb1), sv2v_cast_60B87(1'sb0)};
		end
	end
	wire signed [EXP_WIDTH - 1:0] exponent_a;
	wire signed [EXP_WIDTH - 1:0] exponent_b;
	wire signed [EXP_WIDTH - 1:0] exponent_c;
	wire signed [EXP_WIDTH - 1:0] exponent_addend;
	wire signed [EXP_WIDTH - 1:0] exponent_product;
	wire signed [EXP_WIDTH - 1:0] exponent_difference;
	wire signed [EXP_WIDTH - 1:0] tentative_exponent;
	assign exponent_a = $signed({1'b0, operand_a[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	assign exponent_b = $signed({1'b0, operand_b[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	assign exponent_c = $signed({1'b0, operand_c[EXP_BITS + (MAN_BITS - 1)-:((EXP_BITS + (MAN_BITS - 1)) >= (MAN_BITS + 0) ? ((EXP_BITS + (MAN_BITS - 1)) - (MAN_BITS + 0)) + 1 : ((MAN_BITS + 0) - (EXP_BITS + (MAN_BITS - 1))) + 1)]});
	assign exponent_addend = $signed(exponent_c + $signed({1'b0, ~info_c[7]}));
	assign exponent_product = (info_a[5] || info_b[5] ? 2 - $signed(BIAS) : $signed((((exponent_a + info_a[6]) + exponent_b) + info_b[6]) - $signed(BIAS)));
	assign exponent_difference = exponent_addend - exponent_product;
	assign tentative_exponent = (exponent_difference > 0 ? exponent_addend : exponent_product);
	reg [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt;
	always @(*) begin : addend_shift_amount
		if (exponent_difference <= $signed((-2 * PRECISION_BITS) - 1))
			addend_shamt = (3 * PRECISION_BITS) + 4;
		else if (exponent_difference <= $signed(PRECISION_BITS + 2))
			addend_shamt = $unsigned(($signed(PRECISION_BITS) + 3) - exponent_difference);
		else
			addend_shamt = 0;
	end
	wire [PRECISION_BITS - 1:0] mantissa_a;
	wire [PRECISION_BITS - 1:0] mantissa_b;
	wire [PRECISION_BITS - 1:0] mantissa_c;
	wire [(2 * PRECISION_BITS) - 1:0] product;
	wire [(3 * PRECISION_BITS) + 3:0] product_shifted;
	assign mantissa_a = {info_a[7], operand_a[MAN_BITS - 1-:MAN_BITS]};
	assign mantissa_b = {info_b[7], operand_b[MAN_BITS - 1-:MAN_BITS]};
	assign mantissa_c = {info_c[7], operand_c[MAN_BITS - 1-:MAN_BITS]};
	assign product = mantissa_a * mantissa_b;
	assign product_shifted = product << 2;
	wire [(3 * PRECISION_BITS) + 3:0] addend_after_shift;
	wire [PRECISION_BITS - 1:0] addend_sticky_bits;
	wire sticky_before_add;
	wire [(3 * PRECISION_BITS) + 3:0] addend_shifted;
	wire inject_carry_in;
	assign {addend_after_shift, addend_sticky_bits} = (mantissa_c << ((3 * PRECISION_BITS) + 4)) >> addend_shamt;
	assign sticky_before_add = |addend_sticky_bits;
	assign addend_shifted = (effective_subtraction ? ~addend_after_shift : addend_after_shift);
	assign inject_carry_in = effective_subtraction & ~sticky_before_add;
	wire [(3 * PRECISION_BITS) + 4:0] sum_raw;
	wire sum_carry;
	wire [(3 * PRECISION_BITS) + 3:0] sum;
	wire final_sign;
	assign sum_raw = (product_shifted + addend_shifted) + inject_carry_in;
	assign sum_carry = sum_raw[(3 * PRECISION_BITS) + 4];
	assign sum = (effective_subtraction && ~sum_carry ? -sum_raw : sum_raw);
	assign final_sign = (effective_subtraction && (sum_carry == tentative_sign) ? 1'b1 : (effective_subtraction ? 1'b0 : tentative_sign));
	wire effective_subtraction_q;
	wire signed [EXP_WIDTH - 1:0] exponent_product_q;
	wire signed [EXP_WIDTH - 1:0] exponent_difference_q;
	wire signed [EXP_WIDTH - 1:0] tentative_exponent_q;
	wire [SHIFT_AMOUNT_WIDTH - 1:0] addend_shamt_q;
	wire sticky_before_add_q;
	wire [(3 * PRECISION_BITS) + 3:0] sum_q;
	wire final_sign_q;
	wire [2:0] rnd_mode_q;
	wire result_is_special_q;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] special_result_q;
	wire [4:0] special_status_q;
	reg [0:NUM_MID_REGS] mid_pipe_eff_sub_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_prod_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_exp_diff_q;
	reg signed [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * EXP_WIDTH) + ((NUM_MID_REGS * EXP_WIDTH) - 1) : ((NUM_MID_REGS + 1) * EXP_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * EXP_WIDTH : 0)] mid_pipe_tent_exp_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH) + ((NUM_MID_REGS * SHIFT_AMOUNT_WIDTH) - 1) : ((NUM_MID_REGS + 1) * SHIFT_AMOUNT_WIDTH) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * SHIFT_AMOUNT_WIDTH : 0)] mid_pipe_add_shamt_q;
	reg [0:NUM_MID_REGS] mid_pipe_sticky_q;
	reg [(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? ((1 - NUM_MID_REGS) * ((3 * PRECISION_BITS) + 4)) + ((NUM_MID_REGS * ((3 * PRECISION_BITS) + 4)) - 1) : ((1 - NUM_MID_REGS) * (1 - ((3 * PRECISION_BITS) + 3))) + ((((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) - 1)) : (((3 * PRECISION_BITS) + 3) >= 0 ? ((NUM_MID_REGS + 1) * ((3 * PRECISION_BITS) + 4)) - 1 : ((NUM_MID_REGS + 1) * (1 - ((3 * PRECISION_BITS) + 3))) + ((3 * PRECISION_BITS) + 2))):(0 >= NUM_MID_REGS ? (((3 * PRECISION_BITS) + 3) >= 0 ? NUM_MID_REGS * ((3 * PRECISION_BITS) + 4) : ((3 * PRECISION_BITS) + 3) + (NUM_MID_REGS * (1 - ((3 * PRECISION_BITS) + 3)))) : (((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3))] mid_pipe_sum_q;
	reg [0:NUM_MID_REGS] mid_pipe_final_sign_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_rnd_mode_q;
	reg [0:NUM_MID_REGS] mid_pipe_res_is_spec_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_MID_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] mid_pipe_spec_res_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 5) + ((NUM_MID_REGS * 5) - 1) : ((NUM_MID_REGS + 1) * 5) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 5 : 0)] mid_pipe_spec_stat_q;
	reg [(0 >= NUM_MID_REGS ? ((1 - NUM_MID_REGS) * 3) + ((NUM_MID_REGS * 3) - 1) : ((NUM_MID_REGS + 1) * 3) - 1):(0 >= NUM_MID_REGS ? NUM_MID_REGS * 3 : 0)] mid_pipe_tag_q;
	reg [0:NUM_MID_REGS] mid_pipe_aux_q;
	reg [0:NUM_MID_REGS] mid_pipe_valid_q;
	wire [0:NUM_MID_REGS] mid_pipe_ready;
	wire [1:1] sv2v_tmp_56A72;
	assign sv2v_tmp_56A72 = effective_subtraction;
	always @(*) mid_pipe_eff_sub_q[0] = sv2v_tmp_56A72;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_2D21E;
	assign sv2v_tmp_2D21E = exponent_product;
	always @(*) mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_2D21E;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_00793;
	assign sv2v_tmp_00793 = exponent_difference;
	always @(*) mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_00793;
	wire [EXP_WIDTH * 1:1] sv2v_tmp_B4C85;
	assign sv2v_tmp_B4C85 = tentative_exponent;
	always @(*) mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH] = sv2v_tmp_B4C85;
	wire [SHIFT_AMOUNT_WIDTH * 1:1] sv2v_tmp_83404;
	assign sv2v_tmp_83404 = addend_shamt;
	always @(*) mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] = sv2v_tmp_83404;
	wire [1:1] sv2v_tmp_6F5F7;
	assign sv2v_tmp_6F5F7 = sticky_before_add;
	always @(*) mid_pipe_sticky_q[0] = sv2v_tmp_6F5F7;
	wire [(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)) * 1:1] sv2v_tmp_CEAB3;
	assign sv2v_tmp_CEAB3 = sum;
	always @(*) mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] = sv2v_tmp_CEAB3;
	wire [1:1] sv2v_tmp_D7BD0;
	assign sv2v_tmp_D7BD0 = final_sign;
	always @(*) mid_pipe_final_sign_q[0] = sv2v_tmp_D7BD0;
	wire [3:1] sv2v_tmp_A74E2;
	assign sv2v_tmp_A74E2 = inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_A74E2;
	wire [1:1] sv2v_tmp_7DEC5;
	assign sv2v_tmp_7DEC5 = result_is_special;
	always @(*) mid_pipe_res_is_spec_q[0] = sv2v_tmp_7DEC5;
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_4A83E;
	assign sv2v_tmp_4A83E = special_result;
	always @(*) mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_4A83E;
	wire [5:1] sv2v_tmp_EC01B;
	assign sv2v_tmp_EC01B = special_status;
	always @(*) mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 5+:5] = sv2v_tmp_EC01B;
	wire [3:1] sv2v_tmp_46358;
	assign sv2v_tmp_46358 = inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) mid_pipe_tag_q[(0 >= NUM_MID_REGS ? 0 : NUM_MID_REGS) * 3+:3] = sv2v_tmp_46358;
	wire [1:1] sv2v_tmp_CDA0E;
	assign sv2v_tmp_CDA0E = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) mid_pipe_aux_q[0] = sv2v_tmp_CDA0E;
	wire [1:1] sv2v_tmp_CB10A;
	assign sv2v_tmp_CB10A = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) mid_pipe_valid_q[0] = sv2v_tmp_CB10A;
	assign inp_pipe_ready[NUM_INP_REGS] = mid_pipe_ready[0];
	generate
		for (i = 0; i < NUM_MID_REGS; i = i + 1) begin : gen_inside_pipeline
			wire reg_ena;
			assign mid_pipe_ready[i] = mid_pipe_ready[i + 1] | ~mid_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_valid_q[i + 1] <= 1'b0;
				else
					mid_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (mid_pipe_ready[i] ? mid_pipe_valid_q[i] : mid_pipe_valid_q[i + 1]));
			assign reg_ena = mid_pipe_ready[i] & mid_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_eff_sub_q[i + 1] <= 1'sb0;
				else
					mid_pipe_eff_sub_q[i + 1] <= (reg_ena ? mid_pipe_eff_sub_q[i] : mid_pipe_eff_sub_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= 1'sb0;
				else
					mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH] <= (reg_ena ? mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * EXP_WIDTH+:EXP_WIDTH] : mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * EXP_WIDTH+:EXP_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= 1'sb0;
				else
					mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] <= (reg_ena ? mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH] : mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_sticky_q[i + 1] <= 1'sb0;
				else
					mid_pipe_sticky_q[i + 1] <= (reg_ena ? mid_pipe_sticky_q[i] : mid_pipe_sticky_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= 1'sb0;
				else
					mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] <= (reg_ena ? mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))] : mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_final_sign_q[i + 1] <= 1'sb0;
				else
					mid_pipe_final_sign_q[i + 1] <= (reg_ena ? mid_pipe_final_sign_q[i] : mid_pipe_final_sign_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_res_is_spec_q[i + 1] <= 1'sb0;
				else
					mid_pipe_res_is_spec_q[i + 1] <= (reg_ena ? mid_pipe_res_is_spec_q[i] : mid_pipe_res_is_spec_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5] <= (reg_ena ? mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 5+:5] : mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3] <= (reg_ena ? mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i : NUM_MID_REGS - i) * 3+:3] : mid_pipe_tag_q[(0 >= NUM_MID_REGS ? i + 1 : NUM_MID_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					mid_pipe_aux_q[i + 1] <= 1'b0;
				else
					mid_pipe_aux_q[i + 1] <= (reg_ena ? mid_pipe_aux_q[i] : mid_pipe_aux_q[i + 1]);
		end
	endgenerate
	assign effective_subtraction_q = mid_pipe_eff_sub_q[NUM_MID_REGS];
	assign exponent_product_q = mid_pipe_exp_prod_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign exponent_difference_q = mid_pipe_exp_diff_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign tentative_exponent_q = mid_pipe_tent_exp_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * EXP_WIDTH+:EXP_WIDTH];
	assign addend_shamt_q = mid_pipe_add_shamt_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * SHIFT_AMOUNT_WIDTH+:SHIFT_AMOUNT_WIDTH];
	assign sticky_before_add_q = mid_pipe_sticky_q[NUM_MID_REGS];
	assign sum_q = mid_pipe_sum_q[(((3 * PRECISION_BITS) + 3) >= 0 ? 0 : (3 * PRECISION_BITS) + 3) + ((0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * (((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3)))+:(((3 * PRECISION_BITS) + 3) >= 0 ? (3 * PRECISION_BITS) + 4 : 1 - ((3 * PRECISION_BITS) + 3))];
	assign final_sign_q = mid_pipe_final_sign_q[NUM_MID_REGS];
	assign rnd_mode_q = mid_pipe_rnd_mode_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	assign result_is_special_q = mid_pipe_res_is_spec_q[NUM_MID_REGS];
	assign special_result_q = mid_pipe_spec_res_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	assign special_status_q = mid_pipe_spec_stat_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 5+:5];
	wire [LOWER_SUM_WIDTH - 1:0] sum_lower;
	wire [LZC_RESULT_WIDTH - 1:0] leading_zero_count;
	wire signed [LZC_RESULT_WIDTH:0] leading_zero_count_sgn;
	wire lzc_zeroes;
	reg [SHIFT_AMOUNT_WIDTH - 1:0] norm_shamt;
	reg signed [EXP_WIDTH - 1:0] normalized_exponent;
	wire [(3 * PRECISION_BITS) + 4:0] sum_shifted;
	reg [PRECISION_BITS:0] final_mantissa;
	reg [(2 * PRECISION_BITS) + 2:0] sum_sticky_bits;
	wire sticky_after_norm;
	reg signed [EXP_WIDTH - 1:0] final_exponent;
	assign sum_lower = sum_q[LOWER_SUM_WIDTH - 1:0];
	lzc #(
		.WIDTH(LOWER_SUM_WIDTH),
		.MODE(1)
	) i_lzc(
		.in_i(sum_lower),
		.cnt_o(leading_zero_count),
		.empty_o(lzc_zeroes)
	);
	assign leading_zero_count_sgn = $signed({1'b0, leading_zero_count});
	always @(*) begin : norm_shift_amount
		if ((exponent_difference_q <= 0) || (effective_subtraction_q && (exponent_difference_q <= 2))) begin
			if ((((exponent_product_q - leading_zero_count_sgn) + 1) >= 0) && !lzc_zeroes) begin
				norm_shamt = (PRECISION_BITS + 2) + leading_zero_count;
				normalized_exponent = (exponent_product_q - leading_zero_count_sgn) + 1;
			end
			else begin
				norm_shamt = $unsigned(($signed(PRECISION_BITS) + 2) + exponent_product_q);
				normalized_exponent = 0;
			end
		end
		else begin
			norm_shamt = addend_shamt_q;
			normalized_exponent = tentative_exponent_q;
		end
	end
	assign sum_shifted = sum_q << norm_shamt;
	always @(*) begin : small_norm
		{final_mantissa, sum_sticky_bits} = sum_shifted;
		final_exponent = normalized_exponent;
		if (sum_shifted[(3 * PRECISION_BITS) + 4]) begin
			{final_mantissa, sum_sticky_bits} = sum_shifted >> 1;
			final_exponent = normalized_exponent + 1;
		end
		else if (sum_shifted[(3 * PRECISION_BITS) + 3])
			;
		else if (normalized_exponent > 1) begin
			{final_mantissa, sum_sticky_bits} = sum_shifted << 1;
			final_exponent = normalized_exponent - 1;
		end
		else
			final_exponent = 1'sb0;
	end
	assign sticky_after_norm = |{sum_sticky_bits} | sticky_before_add_q;
	wire pre_round_sign;
	wire [EXP_BITS - 1:0] pre_round_exponent;
	wire [MAN_BITS - 1:0] pre_round_mantissa;
	wire [(EXP_BITS + MAN_BITS) - 1:0] pre_round_abs;
	wire [1:0] round_sticky_bits;
	wire of_before_round;
	wire of_after_round;
	wire uf_before_round;
	wire uf_after_round;
	wire result_zero;
	wire rounded_sign;
	wire [(EXP_BITS + MAN_BITS) - 1:0] rounded_abs;
	assign of_before_round = final_exponent >= ((2 ** EXP_BITS) - 1);
	assign uf_before_round = final_exponent == 0;
	assign pre_round_sign = final_sign_q;
	assign pre_round_exponent = (of_before_round ? (2 ** EXP_BITS) - 2 : $unsigned(final_exponent[EXP_BITS - 1:0]));
	assign pre_round_mantissa = (of_before_round ? {MAN_BITS {1'sb1}} : final_mantissa[MAN_BITS:1]);
	assign pre_round_abs = {pre_round_exponent, pre_round_mantissa};
	assign round_sticky_bits = (of_before_round ? 2'b11 : {final_mantissa[0], sticky_after_norm});
	fpnew_rounding #(.AbsWidth(EXP_BITS + MAN_BITS)) i_fpnew_rounding(
		.abs_value_i(pre_round_abs),
		.sign_i(pre_round_sign),
		.round_sticky_bits_i(round_sticky_bits),
		.rnd_mode_i(rnd_mode_q),
		.effective_subtraction_i(effective_subtraction_q),
		.abs_rounded_o(rounded_abs),
		.sign_o(rounded_sign),
		.exact_zero_o(result_zero)
	);
	assign uf_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb0}};
	assign of_after_round = rounded_abs[(EXP_BITS + MAN_BITS) - 1:MAN_BITS] == {(((EXP_BITS + MAN_BITS) - 1) >= MAN_BITS ? (((EXP_BITS + MAN_BITS) - 1) - MAN_BITS) + 1 : (MAN_BITS - ((EXP_BITS + MAN_BITS) - 1)) + 1) * 1 {1'sb1}};
	wire [WIDTH - 1:0] regular_result;
	wire [4:0] regular_status;
	assign regular_result = {rounded_sign, rounded_abs};
	assign regular_status[4] = 1'b0;
	assign regular_status[3] = 1'b0;
	assign regular_status[2] = of_before_round | of_after_round;
	assign regular_status[1] = uf_after_round & regular_status[0];
	assign regular_status[0] = (|round_sticky_bits | of_before_round) | of_after_round;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	wire [4:0] status_d;
	assign result_d = (result_is_special_q ? special_result_q : regular_result);
	assign status_d = (result_is_special_q ? special_status_q : regular_status);
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 3) + ((NUM_OUT_REGS * 3) - 1) : ((NUM_OUT_REGS + 1) * 3) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 3 : 0)] out_pipe_tag_q;
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_0252C;
	assign sv2v_tmp_0252C = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_0252C;
	wire [5:1] sv2v_tmp_2A843;
	assign sv2v_tmp_2A843 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_2A843;
	wire [3:1] sv2v_tmp_2A8B3;
	assign sv2v_tmp_2A8B3 = mid_pipe_tag_q[(0 >= NUM_MID_REGS ? NUM_MID_REGS : NUM_MID_REGS - NUM_MID_REGS) * 3+:3];
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 3+:3] = sv2v_tmp_2A8B3;
	wire [1:1] sv2v_tmp_9E262;
	assign sv2v_tmp_9E262 = mid_pipe_aux_q[NUM_MID_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_9E262;
	wire [1:1] sv2v_tmp_25EE6;
	assign sv2v_tmp_25EE6 = mid_pipe_valid_q[NUM_MID_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_25EE6;
	assign mid_pipe_ready[NUM_MID_REGS] = out_pipe_ready[0];
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			wire reg_ena;
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 3+:3] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	assign extension_bit_o = 1'b1;
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 3+:3];
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	assign busy_o = |{inp_pipe_valid_q, mid_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_noncomp_CF7FE (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	tag_i,
	aux_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	class_mask_o,
	is_class_o,
	tag_o,
	aux_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] WIDTH = fpnew_pkg_fp_width(FpFormat);
	input wire clk_i;
	input wire rst_ni;
	input wire [(2 * WIDTH) - 1:0] operands_i;
	input wire [1:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	input wire [2:0] tag_i;
	input wire aux_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [9:0] class_mask_o;
	output wire is_class_o;
	output wire [2:0] tag_o;
	output wire aux_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	function automatic [31:0] fpnew_pkg_exp_bits;
		input reg [2:0] fmt;
		fpnew_pkg_exp_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32];
	endfunction
	localparam [31:0] EXP_BITS = fpnew_pkg_exp_bits(FpFormat);
	function automatic [31:0] fpnew_pkg_man_bits;
		input reg [2:0] fmt;
		fpnew_pkg_man_bits = fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32];
	endfunction
	localparam [31:0] MAN_BITS = fpnew_pkg_man_bits(FpFormat);
	localparam NUM_INP_REGS = ((PipeConfig == 2'd0) || (PipeConfig == 2'd2) ? NumPipeRegs : (PipeConfig == 2'd3 ? (NumPipeRegs + 1) / 2 : 0));
	localparam NUM_OUT_REGS = (PipeConfig == 2'd1 ? NumPipeRegs : (PipeConfig == 2'd3 ? NumPipeRegs / 2 : 0));
	reg [((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) - (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH) - 1) : ((((0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)) + 1) * WIDTH) + (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH) - 1)):((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) * WIDTH : (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) * WIDTH)] inp_pipe_operands_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0)] inp_pipe_is_boxed_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_rnd_mode_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * fpnew_pkg_OP_BITS) + ((NUM_INP_REGS * fpnew_pkg_OP_BITS) - 1) : ((NUM_INP_REGS + 1) * fpnew_pkg_OP_BITS) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * fpnew_pkg_OP_BITS : 0)] inp_pipe_op_q;
	reg [0:NUM_INP_REGS] inp_pipe_op_mod_q;
	reg [(0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 3) + ((NUM_INP_REGS * 3) - 1) : ((NUM_INP_REGS + 1) * 3) - 1):(0 >= NUM_INP_REGS ? NUM_INP_REGS * 3 : 0)] inp_pipe_tag_q;
	reg [0:NUM_INP_REGS] inp_pipe_aux_q;
	reg [0:NUM_INP_REGS] inp_pipe_valid_q;
	wire [0:NUM_INP_REGS] inp_pipe_ready;
	wire [2 * WIDTH:1] sv2v_tmp_D1067;
	assign sv2v_tmp_D1067 = operands_i;
	always @(*) inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] = sv2v_tmp_D1067;
	wire [2:1] sv2v_tmp_86D63;
	assign sv2v_tmp_86D63 = is_boxed_i;
	always @(*) inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 2+:2] = sv2v_tmp_86D63;
	wire [3:1] sv2v_tmp_62109;
	assign sv2v_tmp_62109 = rnd_mode_i;
	always @(*) inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_62109;
	wire [4:1] sv2v_tmp_0B797;
	assign sv2v_tmp_0B797 = op_i;
	always @(*) inp_pipe_op_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] = sv2v_tmp_0B797;
	wire [1:1] sv2v_tmp_D1C37;
	assign sv2v_tmp_D1C37 = op_mod_i;
	always @(*) inp_pipe_op_mod_q[0] = sv2v_tmp_D1C37;
	wire [3:1] sv2v_tmp_785B5;
	assign sv2v_tmp_785B5 = tag_i;
	always @(*) inp_pipe_tag_q[(0 >= NUM_INP_REGS ? 0 : NUM_INP_REGS) * 3+:3] = sv2v_tmp_785B5;
	wire [1:1] sv2v_tmp_8D189;
	assign sv2v_tmp_8D189 = aux_i;
	always @(*) inp_pipe_aux_q[0] = sv2v_tmp_8D189;
	wire [1:1] sv2v_tmp_73AEA;
	assign sv2v_tmp_73AEA = in_valid_i;
	always @(*) inp_pipe_valid_q[0] = sv2v_tmp_73AEA;
	assign in_ready_o = inp_pipe_ready[0];
	genvar i;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	generate
		for (i = 0; i < NUM_INP_REGS; i = i + 1) begin : gen_input_pipeline
			wire reg_ena;
			assign inp_pipe_ready[i] = inp_pipe_ready[i + 1] | ~inp_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_valid_q[i + 1] <= 1'b0;
				else
					inp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (inp_pipe_ready[i] ? inp_pipe_valid_q[i] : inp_pipe_valid_q[i + 1]));
			assign reg_ena = inp_pipe_ready[i] & inp_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= 1'sb0;
				else
					inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] <= (reg_ena ? inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2 : ((0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2] : inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2 : ((0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= 1'sb0;
				else
					inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2] <= (reg_ena ? inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 2+:2] : inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 2+:2]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= sv2v_cast_A53F3(0);
				else
					inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] <= (reg_ena ? inp_pipe_op_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] : inp_pipe_op_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_op_mod_q[i + 1] <= 1'sb0;
				else
					inp_pipe_op_mod_q[i + 1] <= (reg_ena ? inp_pipe_op_mod_q[i] : inp_pipe_op_mod_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3] <= (reg_ena ? inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i : NUM_INP_REGS - i) * 3+:3] : inp_pipe_tag_q[(0 >= NUM_INP_REGS ? i + 1 : NUM_INP_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					inp_pipe_aux_q[i + 1] <= 1'b0;
				else
					inp_pipe_aux_q[i + 1] <= (reg_ena ? inp_pipe_aux_q[i] : inp_pipe_aux_q[i + 1]);
		end
	endgenerate
	wire [15:0] info_q;
	fpnew_classifier #(
		.FpFormat(FpFormat),
		.NumOperands(2)
	) i_class_a(
		.operands_i(inp_pipe_operands_q[WIDTH * ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1)))+:WIDTH * 2]),
		.is_boxed_i(inp_pipe_is_boxed_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2+:2]),
		.info_o(info_q)
	);
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_a;
	wire [((1 + EXP_BITS) + MAN_BITS) - 1:0] operand_b;
	wire [7:0] info_a;
	wire [7:0] info_b;
	assign operand_a = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? (0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - (((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	assign operand_b = inp_pipe_operands_q[((0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1) >= (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) ? ((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1 : (0 >= NUM_INP_REGS ? NUM_INP_REGS * 2 : 0) - ((((0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 2) + 1) - (0 >= NUM_INP_REGS ? ((1 - NUM_INP_REGS) * 2) + ((NUM_INP_REGS * 2) - 1) : ((NUM_INP_REGS + 1) * 2) - 1))) * WIDTH+:WIDTH];
	assign info_a = info_q[0+:8];
	assign info_b = info_q[8+:8];
	wire any_operand_inf;
	wire any_operand_nan;
	wire signalling_nan;
	assign any_operand_inf = |{info_a[4], info_b[4]};
	assign any_operand_nan = |{info_a[3], info_b[3]};
	assign signalling_nan = |{info_a[2], info_b[2]};
	wire operands_equal;
	wire operand_a_smaller;
	assign operands_equal = (operand_a == operand_b) || (info_a[5] && info_b[5]);
	assign operand_a_smaller = (operand_a < operand_b) ^ (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] || operand_b[1 + (EXP_BITS + (MAN_BITS - 1))]);
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] sgnj_result;
	wire [4:0] sgnj_status;
	wire sgnj_extension_bit;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic [EXP_BITS - 1:0] sv2v_cast_F2D56;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_F2D56 = inp;
	endfunction
	function automatic [MAN_BITS - 1:0] sv2v_cast_14681;
		input reg [MAN_BITS - 1:0] inp;
		sv2v_cast_14681 = inp;
	endfunction
	function automatic [EXP_BITS - 1:0] sv2v_cast_91364;
		input reg [EXP_BITS - 1:0] inp;
		sv2v_cast_91364 = inp;
	endfunction
	always @(*) begin : sign_injections
		reg sign_a;
		reg sign_b;
		sgnj_result = operand_a;
		if (!info_a[0])
			sgnj_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		sign_a = operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] & info_a[0];
		sign_b = operand_b[1 + (EXP_BITS + (MAN_BITS - 1))] & info_b[0];
		case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
			3'b000: sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_b;
			3'b001: sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = ~sign_b;
			3'b010: sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] = sign_a ^ sign_b;
			3'b011: sgnj_result = operand_a;
			default: sgnj_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
		endcase
	end
	assign sgnj_status = 1'sb0;
	assign sgnj_extension_bit = (inp_pipe_op_mod_q[NUM_INP_REGS] ? sgnj_result[1 + (EXP_BITS + (MAN_BITS - 1))] : 1'b1);
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] minmax_result;
	reg [4:0] minmax_status;
	wire minmax_extension_bit;
	always @(*) begin : min_max
		minmax_status = 1'sb0;
		minmax_status[4] = signalling_nan;
		if (info_a[3] && info_b[3])
			minmax_result = {1'b0, sv2v_cast_F2D56(1'sb1), sv2v_cast_14681(2 ** (MAN_BITS - 1))};
		else if (info_a[3])
			minmax_result = operand_b;
		else if (info_b[3])
			minmax_result = operand_a;
		else
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000: minmax_result = (operand_a_smaller ? operand_a : operand_b);
				3'b001: minmax_result = (operand_a_smaller ? operand_b : operand_a);
				default: minmax_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	assign minmax_extension_bit = 1'b1;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] cmp_result;
	reg [4:0] cmp_status;
	wire cmp_extension_bit;
	always @(*) begin : comparisons
		cmp_result = 1'sb0;
		cmp_status = 1'sb0;
		if (signalling_nan)
			cmp_status[4] = 1'b1;
		else
			case (inp_pipe_rnd_mode_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3])
				3'b000:
					if (any_operand_nan)
						cmp_status[4] = 1'b1;
					else
						cmp_result = (operand_a_smaller | operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b001:
					if (any_operand_nan)
						cmp_status[4] = 1'b1;
					else
						cmp_result = (operand_a_smaller & ~operands_equal) ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				3'b010:
					if (any_operand_nan)
						cmp_result = inp_pipe_op_mod_q[NUM_INP_REGS];
					else
						cmp_result = operands_equal ^ inp_pipe_op_mod_q[NUM_INP_REGS];
				default: cmp_result = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
			endcase
	end
	assign cmp_extension_bit = 1'b0;
	wire [4:0] class_status;
	wire class_extension_bit;
	reg [9:0] class_mask_d;
	always @(*) begin : classify
		if (info_a[7])
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000010 : 10'b0001000000);
		else if (info_a[6])
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000100 : 10'b0000100000);
		else if (info_a[5])
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000001000 : 10'b0000010000);
		else if (info_a[4])
			class_mask_d = (operand_a[1 + (EXP_BITS + (MAN_BITS - 1))] ? 10'b0000000001 : 10'b0010000000);
		else if (info_a[3])
			class_mask_d = (info_a[2] ? 10'b0100000000 : 10'b1000000000);
		else
			class_mask_d = 10'b1000000000;
	end
	assign class_status = 1'sb0;
	assign class_extension_bit = 1'b0;
	reg [((1 + EXP_BITS) + MAN_BITS) - 1:0] result_d;
	reg [4:0] status_d;
	reg extension_bit_d;
	wire is_class_d;
	always @(*) begin : select_result
		case (inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS])
			sv2v_cast_A53F3(6): begin
				result_d = sgnj_result;
				status_d = sgnj_status;
				extension_bit_d = sgnj_extension_bit;
			end
			sv2v_cast_A53F3(7): begin
				result_d = minmax_result;
				status_d = minmax_status;
				extension_bit_d = minmax_extension_bit;
			end
			sv2v_cast_A53F3(8): begin
				result_d = cmp_result;
				status_d = cmp_status;
				extension_bit_d = cmp_extension_bit;
			end
			sv2v_cast_A53F3(9): begin
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				status_d = class_status;
				extension_bit_d = class_extension_bit;
			end
			default: begin
				result_d = {fpnew_pkg_DONT_CARE, sv2v_cast_91364(fpnew_pkg_DONT_CARE), sv2v_cast_14681(fpnew_pkg_DONT_CARE)};
				status_d = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				extension_bit_d = fpnew_pkg_DONT_CARE;
			end
		endcase
	end
	assign is_class_d = inp_pipe_op_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * fpnew_pkg_OP_BITS+:fpnew_pkg_OP_BITS] == sv2v_cast_A53F3(9);
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)) + ((NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS)) - 1) : ((NUM_OUT_REGS + 1) * ((1 + EXP_BITS) + MAN_BITS)) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * ((1 + EXP_BITS) + MAN_BITS) : 0)] out_pipe_result_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 5) + ((NUM_OUT_REGS * 5) - 1) : ((NUM_OUT_REGS + 1) * 5) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 5 : 0)] out_pipe_status_q;
	reg [0:NUM_OUT_REGS] out_pipe_extension_bit_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 10) + ((NUM_OUT_REGS * 10) - 1) : ((NUM_OUT_REGS + 1) * 10) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 10 : 0)] out_pipe_class_mask_q;
	reg [0:NUM_OUT_REGS] out_pipe_is_class_q;
	reg [(0 >= NUM_OUT_REGS ? ((1 - NUM_OUT_REGS) * 3) + ((NUM_OUT_REGS * 3) - 1) : ((NUM_OUT_REGS + 1) * 3) - 1):(0 >= NUM_OUT_REGS ? NUM_OUT_REGS * 3 : 0)] out_pipe_tag_q;
	reg [0:NUM_OUT_REGS] out_pipe_aux_q;
	reg [0:NUM_OUT_REGS] out_pipe_valid_q;
	wire [0:NUM_OUT_REGS] out_pipe_ready;
	wire [((1 + EXP_BITS) + MAN_BITS) * 1:1] sv2v_tmp_07494;
	assign sv2v_tmp_07494 = result_d;
	always @(*) out_pipe_result_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] = sv2v_tmp_07494;
	wire [5:1] sv2v_tmp_CCE43;
	assign sv2v_tmp_CCE43 = status_d;
	always @(*) out_pipe_status_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 5+:5] = sv2v_tmp_CCE43;
	wire [1:1] sv2v_tmp_8E9A9;
	assign sv2v_tmp_8E9A9 = extension_bit_d;
	always @(*) out_pipe_extension_bit_q[0] = sv2v_tmp_8E9A9;
	wire [10:1] sv2v_tmp_94259;
	assign sv2v_tmp_94259 = class_mask_d;
	always @(*) out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 10+:10] = sv2v_tmp_94259;
	wire [1:1] sv2v_tmp_7DF01;
	assign sv2v_tmp_7DF01 = is_class_d;
	always @(*) out_pipe_is_class_q[0] = sv2v_tmp_7DF01;
	wire [3:1] sv2v_tmp_5F9BA;
	assign sv2v_tmp_5F9BA = inp_pipe_tag_q[(0 >= NUM_INP_REGS ? NUM_INP_REGS : NUM_INP_REGS - NUM_INP_REGS) * 3+:3];
	always @(*) out_pipe_tag_q[(0 >= NUM_OUT_REGS ? 0 : NUM_OUT_REGS) * 3+:3] = sv2v_tmp_5F9BA;
	wire [1:1] sv2v_tmp_FA930;
	assign sv2v_tmp_FA930 = inp_pipe_aux_q[NUM_INP_REGS];
	always @(*) out_pipe_aux_q[0] = sv2v_tmp_FA930;
	wire [1:1] sv2v_tmp_2CB8C;
	assign sv2v_tmp_2CB8C = inp_pipe_valid_q[NUM_INP_REGS];
	always @(*) out_pipe_valid_q[0] = sv2v_tmp_2CB8C;
	assign inp_pipe_ready[NUM_INP_REGS] = out_pipe_ready[0];
	generate
		for (i = 0; i < NUM_OUT_REGS; i = i + 1) begin : gen_output_pipeline
			wire reg_ena;
			assign out_pipe_ready[i] = out_pipe_ready[i + 1] | ~out_pipe_valid_q[i + 1];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_valid_q[i + 1] <= 1'b0;
				else
					out_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (out_pipe_ready[i] ? out_pipe_valid_q[i] : out_pipe_valid_q[i + 1]));
			assign reg_ena = out_pipe_ready[i] & out_pipe_valid_q[i];
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= 1'sb0;
				else
					out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] <= (reg_ena ? out_pipe_result_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS] : out_pipe_result_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= 1'sb0;
				else
					out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5] <= (reg_ena ? out_pipe_status_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 5+:5] : out_pipe_status_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 5+:5]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_extension_bit_q[i + 1] <= 1'sb0;
				else
					out_pipe_extension_bit_q[i + 1] <= (reg_ena ? out_pipe_extension_bit_q[i] : out_pipe_extension_bit_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= 10'b1000000000;
				else
					out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10] <= (reg_ena ? out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 10+:10] : out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 10+:10]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_is_class_q[i + 1] <= 1'sb0;
				else
					out_pipe_is_class_q[i + 1] <= (reg_ena ? out_pipe_is_class_q[i] : out_pipe_is_class_q[i + 1]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= 3'b000;
				else
					out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3] <= (reg_ena ? out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i : NUM_OUT_REGS - i) * 3+:3] : out_pipe_tag_q[(0 >= NUM_OUT_REGS ? i + 1 : NUM_OUT_REGS - (i + 1)) * 3+:3]);
			always @(posedge clk_i or negedge rst_ni)
				if (!rst_ni)
					out_pipe_aux_q[i + 1] <= 1'b0;
				else
					out_pipe_aux_q[i + 1] <= (reg_ena ? out_pipe_aux_q[i] : out_pipe_aux_q[i + 1]);
		end
	endgenerate
	assign out_pipe_ready[NUM_OUT_REGS] = out_ready_i;
	assign result_o = out_pipe_result_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * ((1 + EXP_BITS) + MAN_BITS)+:(1 + EXP_BITS) + MAN_BITS];
	assign status_o = out_pipe_status_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 5+:5];
	assign extension_bit_o = out_pipe_extension_bit_q[NUM_OUT_REGS];
	assign class_mask_o = out_pipe_class_mask_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 10+:10];
	assign is_class_o = out_pipe_is_class_q[NUM_OUT_REGS];
	assign tag_o = out_pipe_tag_q[(0 >= NUM_OUT_REGS ? NUM_OUT_REGS : NUM_OUT_REGS - NUM_OUT_REGS) * 3+:3];
	assign aux_o = out_pipe_aux_q[NUM_OUT_REGS];
	assign out_valid_o = out_pipe_valid_q[NUM_OUT_REGS];
	assign busy_o = |{inp_pipe_valid_q, out_pipe_valid_q};
endmodule
module fpnew_opgroup_block_AC56A (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [1:0] OpGroup = 2'd0;
	parameter [31:0] Width = 32;
	parameter [0:0] EnableVectors = 1'b1;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	parameter [0:4] FpFmtMask = 1'sb1;
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	parameter [0:3] IntFmtMask = 1'sb1;
	parameter [159:0] FmtPipeRegs = {fpnew_pkg_NUM_FP_FORMATS {32'd0}};
	parameter [9:0] FmtUnitTypes = {fpnew_pkg_NUM_FP_FORMATS {2'd1}};
	parameter [1:0] PipeConfig = 2'd0;
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	function automatic [31:0] fpnew_pkg_num_operands;
		input reg [1:0] grp;
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	input wire clk_i;
	input wire rst_ni;
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	input wire [2:0] src_fmt_i;
	input wire [2:0] dst_fmt_i;
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	input wire [1:0] int_fmt_i;
	input wire vectorial_op_i;
	input wire [2:0] tag_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [Width - 1:0] result_o;
	output wire [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	wire [4:0] fmt_in_ready;
	wire [4:0] fmt_out_valid;
	wire [4:0] fmt_out_ready;
	wire [4:0] fmt_busy;
	wire [((Width + 8) >= 0 ? (5 * (Width + 9)) - 1 : (5 * (1 - (Width + 8))) + (Width + 7)):((Width + 8) >= 0 ? 0 : Width + 8)] fmt_outputs;
	assign in_ready_o = in_valid_i & fmt_in_ready[dst_fmt_i];
	genvar fmt;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	function automatic fpnew_pkg_any_enabled_multi;
		input reg [9:0] types;
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				begin : sv2v_autoblock_2
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_any_enabled_multi = 1'b1;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_any_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [2:0] fpnew_pkg_get_first_enabled_multi;
		input reg [9:0] types;
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			begin : sv2v_autoblock_3
				reg [31:0] i;
				begin : sv2v_autoblock_4
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(i);
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_get_first_enabled_multi = sv2v_cast_0BC43(0);
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic fpnew_pkg_is_first_enabled_multi;
		input reg [2:0] fmt;
		input reg [9:0] types;
		input reg [0:4] cfg;
		reg [0:1] _sv2v_jump;
		begin
			_sv2v_jump = 2'b00;
			begin : sv2v_autoblock_5
				reg [31:0] i;
				begin : sv2v_autoblock_6
					reg [31:0] _sv2v_value_on_break;
					for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
						if (_sv2v_jump < 2'b10) begin
							_sv2v_jump = 2'b00;
							if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2)) begin
								fpnew_pkg_is_first_enabled_multi = sv2v_cast_0BC43(i) == fmt;
								_sv2v_jump = 2'b11;
							end
							_sv2v_value_on_break = i;
						end
					if (!(_sv2v_jump < 2'b10))
						i = _sv2v_value_on_break;
					if (_sv2v_jump != 2'b11)
						_sv2v_jump = 2'b00;
				end
			end
			if (_sv2v_jump == 2'b00) begin
				fpnew_pkg_is_first_enabled_multi = 1'b0;
				_sv2v_jump = 2'b11;
			end
		end
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	function automatic [2:0] sv2v_cast_3;
		input reg [2:0] inp;
		sv2v_cast_3 = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_parallel_slices
			localparam [0:0] ANY_MERGED = fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask);
			localparam [0:0] IS_FIRST_MERGED = fpnew_pkg_is_first_enabled_multi(sv2v_cast_0BC43(fmt), FmtUnitTypes, FpFmtMask);
			if (FpFmtMask[fmt] && (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd1)) begin : active_format
				wire in_valid;
				assign in_valid = in_valid_i & (dst_fmt_i == fmt);
				fpnew_opgroup_fmt_slice_BAB27 #(
					.OpGroup(OpGroup),
					.FpFormat(sv2v_cast_0BC43(fmt)),
					.Width(Width),
					.EnableVectors(EnableVectors),
					.NumPipeRegs(FmtPipeRegs[(4 - fmt) * 32+:32]),
					.PipeConfig(PipeConfig)
				) i_fmt_slice(
					.clk_i(clk_i),
					.rst_ni(rst_ni),
					.operands_i(operands_i),
					.is_boxed_i(is_boxed_i[fmt * NUM_OPERANDS+:NUM_OPERANDS]),
					.rnd_mode_i(rnd_mode_i),
					.op_i(op_i),
					.op_mod_i(op_mod_i),
					.vectorial_op_i(vectorial_op_i),
					.tag_i(tag_i),
					.in_valid_i(in_valid),
					.in_ready_o(fmt_in_ready[fmt]),
					.flush_i(flush_i),
					.result_o(fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8)) : (((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8))) + ((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))) - 1)-:((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))]),
					.status_o(fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0)) + 4)-:5]),
					.extension_bit_o(fmt_outputs[(fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 3 : Width + 5)]),
					.tag_o(fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6)) + 2)-:3]),
					.out_valid_o(fmt_out_valid[fmt]),
					.out_ready_i(fmt_out_ready[fmt]),
					.busy_o(fmt_busy[fmt])
				);
			end
			else if ((FpFmtMask[fmt] && ANY_MERGED) && !IS_FIRST_MERGED) begin : merged_unused
				assign fmt_in_ready[fmt] = fmt_in_ready[fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask)];
				assign fmt_out_valid[fmt] = 1'b0;
				assign fmt_busy[fmt] = 1'b0;
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8)) : (((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8))) + ((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))) - 1)-:((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))] = {Width {fpnew_pkg_DONT_CARE}};
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				assign fmt_outputs[(fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 3 : Width + 5)] = fpnew_pkg_DONT_CARE;
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6)) + 2)-:3] = sv2v_cast_3(fpnew_pkg_DONT_CARE);
			end
			else if (!FpFmtMask[fmt] || (FmtUnitTypes[(4 - fmt) * 2+:2] == 2'd0)) begin : disable_fmt
				assign fmt_in_ready[fmt] = 1'b0;
				assign fmt_out_valid[fmt] = 1'b0;
				assign fmt_busy[fmt] = 1'b0;
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8)) : (((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8))) + ((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))) - 1)-:((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))] = {Width {fpnew_pkg_DONT_CARE}};
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0)) + 4)-:5] = {fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE, fpnew_pkg_DONT_CARE};
				assign fmt_outputs[(fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 3 : Width + 5)] = fpnew_pkg_DONT_CARE;
				assign fmt_outputs[((Width + 8) >= 0 ? (fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6) : ((fmt * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6)) + 2)-:3] = sv2v_cast_3(fpnew_pkg_DONT_CARE);
			end
		end
	endgenerate
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_get_num_regs_multi;
		input reg [159:0] regs;
		input reg [9:0] types;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_7
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i] && (types[(4 - i) * 2+:2] == 2'd2))
						res = fpnew_pkg_maximum(res, regs[(4 - i) * 32+:32]);
			end
			fpnew_pkg_get_num_regs_multi = res;
		end
	endfunction
	generate
		if (fpnew_pkg_any_enabled_multi(FmtUnitTypes, FpFmtMask)) begin : gen_merged_slice
			localparam FMT = fpnew_pkg_get_first_enabled_multi(FmtUnitTypes, FpFmtMask);
			localparam REG = fpnew_pkg_get_num_regs_multi(FmtPipeRegs, FmtUnitTypes, FpFmtMask);
			wire in_valid;
			assign in_valid = in_valid_i & (FmtUnitTypes[(4 - dst_fmt_i) * 2+:2] == 2'd2);
			fpnew_opgroup_multifmt_slice_F1CBB #(
				.OpGroup(OpGroup),
				.Width(Width),
				.FpFmtConfig(FpFmtMask),
				.IntFmtConfig(IntFmtMask),
				.EnableVectors(EnableVectors),
				.NumPipeRegs(REG),
				.PipeConfig(PipeConfig)
			) i_multifmt_slice(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i),
				.is_boxed_i(is_boxed_i),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(fmt_in_ready[FMT]),
				.flush_i(flush_i),
				.result_o(fmt_outputs[((Width + 8) >= 0 ? (FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8)) : (((FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? Width + 8 : (Width + 8) - (Width + 8))) + ((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))) - 1)-:((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))]),
				.status_o(fmt_outputs[((Width + 8) >= 0 ? (FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0) : ((FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 8 : Width + 0)) + 4)-:5]),
				.extension_bit_o(fmt_outputs[(FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 3 : Width + 5)]),
				.tag_o(fmt_outputs[((Width + 8) >= 0 ? (FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6) : ((FMT * ((Width + 8) >= 0 ? Width + 9 : 1 - (Width + 8))) + ((Width + 8) >= 0 ? 2 : Width + 6)) + 2)-:3]),
				.out_valid_o(fmt_out_valid[FMT]),
				.out_ready_i(fmt_out_ready[FMT]),
				.busy_o(fmt_busy[FMT])
			);
		end
	endgenerate
	wire [Width + 8:0] arbiter_output;
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_FORMATS;
	localparam [2:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_36817_A990F #(
		.DataType_Width(Width),
		.NumIn(NUM_FORMATS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(fmt_out_valid),
		.gnt_o(fmt_out_ready),
		.data_i(fmt_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	assign result_o = arbiter_output[Width + 8-:((Width + 8) >= 9 ? Width + 0 : 10 - (Width + 8))];
	assign status_o = arbiter_output[8-:5];
	assign extension_bit_o = arbiter_output[3];
	assign tag_o = arbiter_output[2-:3];
	assign busy_o = |fmt_busy;
endmodule
module fpnew_opgroup_fmt_slice_BAB27 (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [1:0] OpGroup = 2'd0;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	parameter [2:0] FpFormat = sv2v_cast_0BC43(0);
	parameter [31:0] Width = 32;
	parameter [0:0] EnableVectors = 1'b1;
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	function automatic [31:0] fpnew_pkg_num_operands;
		input reg [1:0] grp;
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	input wire clk_i;
	input wire rst_ni;
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	input wire [NUM_OPERANDS - 1:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	input wire vectorial_op_i;
	input wire [2:0] tag_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [Width - 1:0] result_o;
	output reg [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(FpFormat);
	function automatic [31:0] fpnew_pkg_num_lanes;
		input reg [31:0] width;
		input reg [2:0] fmt;
		input reg vec;
		fpnew_pkg_num_lanes = (vec ? width / fpnew_pkg_fp_width(fmt) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_num_lanes(Width, FpFormat, EnableVectors);
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	wire vectorial_op;
	wire [(NUM_LANES * FP_WIDTH) - 1:0] slice_result;
	wire [Width - 1:0] slice_regular_result;
	wire [Width - 1:0] slice_class_result;
	wire [Width - 1:0] slice_vec_class_result;
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	wire [NUM_LANES - 1:0] lane_ext_bit;
	wire [(NUM_LANES * 10) - 1:0] lane_class_mask;
	wire [(NUM_LANES * 3) - 1:0] lane_tags;
	wire [NUM_LANES - 1:0] lane_vectorial;
	wire [NUM_LANES - 1:0] lane_busy;
	wire [NUM_LANES - 1:0] lane_is_class;
	wire result_is_vector;
	wire result_is_class;
	assign in_ready_o = lane_in_ready[0];
	assign vectorial_op = vectorial_op_i & EnableVectors;
	genvar lane;
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			wire [FP_WIDTH - 1:0] local_result;
			wire local_sign;
			if ((lane == 0) || EnableVectors) begin : active_lane
				wire in_valid;
				wire out_valid;
				wire out_ready;
				reg [(NUM_OPERANDS * FP_WIDTH) - 1:0] local_operands;
				wire [FP_WIDTH - 1:0] op_result;
				wire [4:0] op_status;
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				always @(*) begin : prepare_input
					begin : sv2v_autoblock_1
						reg signed [31:0] i;
						for (i = 0; i < sv2v_cast_32_signed(NUM_OPERANDS); i = i + 1)
							local_operands[i * FP_WIDTH+:FP_WIDTH] = operands_i[(i * Width) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (($unsigned(lane) + 1) * FP_WIDTH) - 1 : (((($unsigned(lane) + 1) * FP_WIDTH) - 1) + (((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:(((($unsigned(lane) + 1) * FP_WIDTH) - 1) >= ($unsigned(lane) * FP_WIDTH) ? (((($unsigned(lane) + 1) * FP_WIDTH) - 1) - ($unsigned(lane) * FP_WIDTH)) + 1 : (($unsigned(lane) * FP_WIDTH) - ((($unsigned(lane) + 1) * FP_WIDTH) - 1)) + 1)];
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					fpnew_fma_F8EAE #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fma(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane * 3+:3]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
					assign lane_is_class[lane] = 1'b0;
					assign lane_class_mask[lane * 10+:10] = 10'b0000000001;
				end
				// else if (OpGroup == 2'd1) begin
				// 	;
				// end
				else if (OpGroup == 2'd2) begin : lane_instance
					fpnew_noncomp_CF7FE #(
						.FpFormat(FpFormat),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_noncomp(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i[NUM_OPERANDS - 1:0]),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.tag_i(tag_i),
						.aux_i(vectorial_op),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.class_mask_o(lane_class_mask[lane * 10+:10]),
						.is_class_o(lane_is_class[lane]),
						.tag_o(lane_tags[lane * 3+:3]),
						.aux_o(lane_vectorial[lane]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				assign local_result = (lane_out_valid[lane] ? op_result : {FP_WIDTH {lane_ext_bit[0]}});
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : genblk1
				assign lane_out_valid[lane] = 1'b0;
				assign lane_in_ready[lane] = 1'b0;
				assign local_result = {FP_WIDTH {lane_ext_bit[0]}};
				assign lane_status[lane * 5+:5] = 1'sb0;
				assign lane_busy[lane] = 1'b0;
				assign lane_is_class[lane] = 1'b0;
			end
			assign slice_result[(($unsigned(lane) + 1) * FP_WIDTH) - 1:$unsigned(lane) * FP_WIDTH] = local_result;
			if (((lane + 1) * 8) <= Width) begin : vectorial_class
				assign local_sign = (((lane_class_mask[lane * 10+:10] == 10'b0000000001) || (lane_class_mask[lane * 10+:10] == 10'b0000000010)) || (lane_class_mask[lane * 10+:10] == 10'b0000000100)) || (lane_class_mask[lane * 10+:10] == 10'b0000001000);
				assign slice_vec_class_result[((lane + 1) * 8) - 1:lane * 8] = {local_sign, ~local_sign, lane_class_mask[lane * 10+:10] == 10'b1000000000, lane_class_mask[lane * 10+:10] == 10'b0100000000, (lane_class_mask[lane * 10+:10] == 10'b0000010000) || (lane_class_mask[lane * 10+:10] == 10'b0000001000), (lane_class_mask[lane * 10+:10] == 10'b0000100000) || (lane_class_mask[lane * 10+:10] == 10'b0000000100), (lane_class_mask[lane * 10+:10] == 10'b0001000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000010), (lane_class_mask[lane * 10+:10] == 10'b0010000000) || (lane_class_mask[lane * 10+:10] == 10'b0000000001)};
			end
		end
	endgenerate
	assign result_is_vector = lane_vectorial[0];
	assign result_is_class = lane_is_class[0];
	assign slice_regular_result = $signed({extension_bit_o, slice_result});
	localparam [31:0] CLASS_VEC_BITS = ((NUM_LANES * 8) > Width ? 8 * (Width / 8) : NUM_LANES * 8);
	generate
		if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
			assign slice_vec_class_result[Width - 1:CLASS_VEC_BITS] = 1'sb0;
		end
	endgenerate
	assign slice_class_result = (result_is_vector ? slice_vec_class_result : lane_class_mask[0+:10]);
	assign result_o = (result_is_class ? slice_class_result : slice_regular_result);
	assign extension_bit_o = lane_ext_bit[0];
	assign tag_o = lane_tags[0+:3];
	assign busy_o = |lane_busy;
	assign out_valid_o = lane_out_valid[0];
	always @(*) begin : output_processing
		reg [4:0] temp_status;
		temp_status = 1'sb0;
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				temp_status = temp_status | lane_status[i * 5+:5];
		end
		status_o = temp_status;
	end
endmodule
module fpnew_opgroup_multifmt_slice_F1CBB (
	clk_i,
	rst_ni,
	operands_i,
	is_boxed_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	extension_bit_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	parameter [1:0] OpGroup = 2'd3;
	parameter [31:0] Width = 64;
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	parameter [0:4] FpFmtConfig = 1'sb1;
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	parameter [0:3] IntFmtConfig = 1'sb1;
	parameter [0:0] EnableVectors = 1'b1;
	parameter [31:0] NumPipeRegs = 0;
	parameter [1:0] PipeConfig = 2'd0;
	function automatic [31:0] fpnew_pkg_num_operands;
		input reg [1:0] grp;
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	localparam [31:0] NUM_OPERANDS = fpnew_pkg_num_operands(OpGroup);
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	input wire clk_i;
	input wire rst_ni;
	input wire [(NUM_OPERANDS * Width) - 1:0] operands_i;
	input wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	input wire [2:0] src_fmt_i;
	input wire [2:0] dst_fmt_i;
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	input wire [1:0] int_fmt_i;
	input wire vectorial_op_i;
	input wire [2:0] tag_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [Width - 1:0] result_o;
	output reg [4:0] status_o;
	output wire extension_bit_o;
	output wire [2:0] tag_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic signed [31:0] fpnew_pkg_maximum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_maximum = (a > b ? a : b);
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_max_fp_width;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_1
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						res = $unsigned(fpnew_pkg_maximum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_max_fp_width = res;
		end
	endfunction
	localparam [31:0] MAX_FP_WIDTH = fpnew_pkg_max_fp_width(FpFmtConfig);
	function automatic [1:0] sv2v_cast_87CC5;
		input reg [1:0] inp;
		sv2v_cast_87CC5 = inp;
	endfunction
	function automatic [31:0] fpnew_pkg_int_width;
		input reg [1:0] ifmt;
		case (ifmt)
			sv2v_cast_87CC5(0): fpnew_pkg_int_width = 8;
			sv2v_cast_87CC5(1): fpnew_pkg_int_width = 16;
			sv2v_cast_87CC5(2): fpnew_pkg_int_width = 32;
			sv2v_cast_87CC5(3): fpnew_pkg_int_width = 64;
		endcase
	endfunction
	function automatic [31:0] fpnew_pkg_max_int_width;
		input reg [0:3] cfg;
		reg [31:0] res;
		begin
			res = 0;
			begin : sv2v_autoblock_2
				reg signed [31:0] ifmt;
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					if (cfg[ifmt])
						res = fpnew_pkg_maximum(res, fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)));
			end
			fpnew_pkg_max_int_width = res;
		end
	endfunction
	localparam [31:0] MAX_INT_WIDTH = fpnew_pkg_max_int_width(IntFmtConfig);
	function automatic signed [31:0] fpnew_pkg_minimum;
		input reg signed [31:0] a;
		input reg signed [31:0] b;
		fpnew_pkg_minimum = (a < b ? a : b);
	endfunction
	function automatic [31:0] fpnew_pkg_min_fp_width;
		input reg [0:4] cfg;
		reg [31:0] res;
		begin
			res = fpnew_pkg_max_fp_width(cfg);
			begin : sv2v_autoblock_3
				reg [31:0] i;
				for (i = 0; i < fpnew_pkg_NUM_FP_FORMATS; i = i + 1)
					if (cfg[i])
						res = $unsigned(fpnew_pkg_minimum(res, fpnew_pkg_fp_width(sv2v_cast_0BC43(i))));
			end
			fpnew_pkg_min_fp_width = res;
		end
	endfunction
	function automatic [31:0] fpnew_pkg_max_num_lanes;
		input reg [31:0] width;
		input reg [0:4] cfg;
		input reg vec;
		fpnew_pkg_max_num_lanes = (vec ? width / fpnew_pkg_min_fp_width(cfg) : 1);
	endfunction
	localparam [31:0] NUM_LANES = fpnew_pkg_max_num_lanes(Width, FpFmtConfig, 1'b1);
	localparam [31:0] NUM_INT_FORMATS = fpnew_pkg_NUM_INT_FORMATS;
	localparam [31:0] FMT_BITS = fpnew_pkg_maximum(3, 2);
	localparam [31:0] AUX_BITS = FMT_BITS + 2;
	wire [NUM_LANES - 1:0] lane_in_ready;
	wire [NUM_LANES - 1:0] lane_out_valid;
	wire vectorial_op;
	wire [FMT_BITS - 1:0] dst_fmt;
	wire [AUX_BITS - 1:0] aux_data;
	wire dst_fmt_is_int;
	wire dst_is_cpk;
	wire [1:0] dst_vec_op;
	wire [2:0] target_aux_d;
	wire [2:0] target_aux_q;
	wire is_up_cast;
	wire is_down_cast;
	wire [(NUM_FORMATS * Width) - 1:0] fmt_slice_result;
	wire [(NUM_INT_FORMATS * Width) - 1:0] ifmt_slice_result;
	wire [Width - 1:0] conv_slice_result;
	wire [Width - 1:0] conv_target_d;
	wire [Width - 1:0] conv_target_q;
	wire [(NUM_LANES * 5) - 1:0] lane_status;
	wire [NUM_LANES - 1:0] lane_ext_bit;
	wire [(NUM_LANES * 3) - 1:0] lane_tags;
	wire [(NUM_LANES * AUX_BITS) - 1:0] lane_aux;
	wire [NUM_LANES - 1:0] lane_busy;
	wire result_is_vector;
	wire [FMT_BITS - 1:0] result_fmt;
	wire result_fmt_is_int;
	wire result_is_cpk;
	wire [1:0] result_vec_op;
	assign in_ready_o = lane_in_ready[0];
	assign vectorial_op = vectorial_op_i & EnableVectors;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	assign dst_fmt_is_int = (OpGroup == 2'd3) & (op_i == sv2v_cast_A53F3(11));
	assign dst_is_cpk = (OpGroup == 2'd3) & ((op_i == sv2v_cast_A53F3(13)) || (op_i == sv2v_cast_A53F3(14)));
	assign dst_vec_op = (OpGroup == 2'd3) & {op_i == sv2v_cast_A53F3(14), op_mod_i};
	assign is_up_cast = fpnew_pkg_fp_width(dst_fmt_i) > fpnew_pkg_fp_width(src_fmt_i);
	assign is_down_cast = fpnew_pkg_fp_width(dst_fmt_i) < fpnew_pkg_fp_width(src_fmt_i);
	assign dst_fmt = (dst_fmt_is_int ? int_fmt_i : dst_fmt_i);
	assign aux_data = {dst_fmt_is_int, vectorial_op, dst_fmt};
	assign target_aux_d = {dst_vec_op, dst_is_cpk};
	generate
		if (OpGroup == 2'd3) begin : conv_target
			assign conv_target_d = (dst_is_cpk ? operands_i[2 * Width+:Width] : operands_i[Width+:Width]);
		end
	endgenerate
	reg [4:0] is_boxed_1op;
	reg [9:0] is_boxed_2op;
	always @(*) begin : boxed_2op
		begin : sv2v_autoblock_4
			reg signed [31:0] fmt;
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
				begin
					is_boxed_1op[fmt] = is_boxed_i[fmt * NUM_OPERANDS];
					is_boxed_2op[fmt * 2+:2] = is_boxed_i[(fmt * NUM_OPERANDS) + 1-:2];
				end
		end
	end
	genvar lane;
	localparam [0:4] fpnew_pkg_CPK_FORMATS = 5'b11000;
	function automatic [0:4] fpnew_pkg_get_conv_lane_formats;
		input reg [31:0] width;
		input reg [0:4] cfg;
		input reg [31:0] lane_no;
		reg [0:4] res;
		begin
			begin : sv2v_autoblock_5
				reg [31:0] fmt;
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					res[fmt] = cfg[fmt] && (((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no) || (fpnew_pkg_CPK_FORMATS[fmt] && (lane_no < 2)));
			end
			fpnew_pkg_get_conv_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_conv_lane_int_formats;
		input reg [31:0] width;
		input reg [0:4] cfg;
		input reg [0:3] icfg;
		input reg [31:0] lane_no;
		reg [0:3] res;
		reg [0:4] lanefmts;
		begin
			res = 1'sb0;
			lanefmts = fpnew_pkg_get_conv_lane_formats(width, cfg, lane_no);
			begin : sv2v_autoblock_6
				reg [31:0] ifmt;
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_7
						reg [31:0] fmt;
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							res[ifmt] = res[ifmt] | ((icfg[ifmt] && lanefmts[fmt]) && (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt))));
					end
			end
			fpnew_pkg_get_conv_lane_int_formats = res;
		end
	endfunction
	function automatic [0:4] fpnew_pkg_get_lane_formats;
		input reg [31:0] width;
		input reg [0:4] cfg;
		input reg [31:0] lane_no;
		reg [0:4] res;
		begin
			begin : sv2v_autoblock_8
				reg [31:0] fmt;
				for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
					res[fmt] = cfg[fmt] & ((width / fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt))) > lane_no);
			end
			fpnew_pkg_get_lane_formats = res;
		end
	endfunction
	function automatic [0:3] fpnew_pkg_get_lane_int_formats;
		input reg [31:0] width;
		input reg [0:4] cfg;
		input reg [0:3] icfg;
		input reg [31:0] lane_no;
		reg [0:3] res;
		reg [0:4] lanefmts;
		begin
			res = 1'sb0;
			lanefmts = fpnew_pkg_get_lane_formats(width, cfg, lane_no);
			begin : sv2v_autoblock_9
				reg [31:0] ifmt;
				for (ifmt = 0; ifmt < fpnew_pkg_NUM_INT_FORMATS; ifmt = ifmt + 1)
					begin : sv2v_autoblock_10
						reg [31:0] fmt;
						for (fmt = 0; fmt < fpnew_pkg_NUM_FP_FORMATS; fmt = fmt + 1)
							if (fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt)) == fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt)))
								res[ifmt] = res[ifmt] | (icfg[ifmt] && lanefmts[fmt]);
					end
			end
			fpnew_pkg_get_lane_int_formats = res;
		end
	endfunction
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [4:0] sv2v_cast_F8FCA;
		input reg [4:0] inp;
		sv2v_cast_F8FCA = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (lane = 0; lane < sv2v_cast_32_signed(NUM_LANES); lane = lane + 1) begin : gen_num_lanes
			localparam [31:0] LANE = $unsigned(lane);
			localparam [0:4] ACTIVE_FORMATS = fpnew_pkg_get_lane_formats(Width, FpFmtConfig, LANE);
			localparam [0:3] ACTIVE_INT_FORMATS = fpnew_pkg_get_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			localparam [31:0] MAX_WIDTH = fpnew_pkg_max_fp_width(ACTIVE_FORMATS);
			localparam [0:4] CONV_FORMATS = fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, LANE);
			localparam [0:3] CONV_INT_FORMATS = fpnew_pkg_get_conv_lane_int_formats(Width, FpFmtConfig, IntFmtConfig, LANE);
			localparam [31:0] CONV_WIDTH = fpnew_pkg_max_fp_width(CONV_FORMATS);
			localparam [0:4] LANE_FORMATS = (OpGroup == 2'd3 ? CONV_FORMATS : ACTIVE_FORMATS);
			localparam [31:0] LANE_WIDTH = (OpGroup == 2'd3 ? CONV_WIDTH : MAX_WIDTH);
			wire [LANE_WIDTH - 1:0] local_result;
			if ((lane == 0) || EnableVectors) begin : active_lane
				wire in_valid;
				wire out_valid;
				wire out_ready;
				reg [(NUM_OPERANDS * LANE_WIDTH) - 1:0] local_operands;
				wire [LANE_WIDTH - 1:0] op_result;
				wire [4:0] op_status;
				assign in_valid = in_valid_i & ((lane == 0) | vectorial_op);
				always @(*) begin : prepare_input
					begin : sv2v_autoblock_11
						reg [31:0] i;
						for (i = 0; i < NUM_OPERANDS; i = i + 1)
							local_operands[i * (OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[i * Width+:Width] >> (LANE * fpnew_pkg_fp_width(src_fmt_i));
					end
					if (OpGroup == 2'd3) begin
						if (op_i == sv2v_cast_A53F3(12))
							local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> (LANE * fpnew_pkg_int_width(int_fmt_i));
						else if (op_i == sv2v_cast_A53F3(10)) begin
							if ((vectorial_op && op_mod_i) && is_up_cast)
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[0+:Width] >> ((LANE * fpnew_pkg_fp_width(src_fmt_i)) + (MAX_FP_WIDTH / 2));
						end
						else if (dst_is_cpk) begin
							if (lane == 1)
								local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))] = operands_i[Width + (LANE_WIDTH - 1)-:LANE_WIDTH];
						end
					end
				end
				if (OpGroup == 2'd0) begin : lane_instance
					fpnew_fma_multi_FF0B0_361DB #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_fma_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands),
						.is_boxed_i(is_boxed_i),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane * 3+:3]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				else if (OpGroup == 2'd1) begin : lane_instance
					fpnew_divsqrt_multi_C04AD_31CA4 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_divsqrt_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) * 2]),
						.is_boxed_i(is_boxed_2op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.dst_fmt_i(dst_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane * 3+:3]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				// else if (OpGroup == 2'd2) begin
				// 	;
				// end
				else if (OpGroup == 2'd3) begin : lane_instance
					fpnew_cast_multi_5BCFE_D3186 #(
						.AuxType_AUX_BITS(AUX_BITS),
						.FpFmtConfig(LANE_FORMATS),
						.IntFmtConfig(CONV_INT_FORMATS),
						.NumPipeRegs(NumPipeRegs),
						.PipeConfig(PipeConfig)
					) i_fpnew_cast_multi(
						.clk_i(clk_i),
						.rst_ni(rst_ni),
						.operands_i(local_operands[0+:(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))) : fpnew_pkg_max_fp_width(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))]),
						.is_boxed_i(is_boxed_1op),
						.rnd_mode_i(rnd_mode_i),
						.op_i(op_i),
						.op_mod_i(op_mod_i),
						.src_fmt_i(src_fmt_i),
						.dst_fmt_i(dst_fmt_i),
						.int_fmt_i(int_fmt_i),
						.tag_i(tag_i),
						.aux_i(aux_data),
						.in_valid_i(in_valid),
						.in_ready_o(lane_in_ready[lane]),
						.flush_i(flush_i),
						.result_o(op_result),
						.status_o(op_status),
						.extension_bit_o(lane_ext_bit[lane]),
						.tag_o(lane_tags[lane * 3+:3]),
						.aux_o(lane_aux[lane * AUX_BITS+:AUX_BITS]),
						.out_valid_o(out_valid),
						.out_ready_i(out_ready),
						.busy_o(lane_busy[lane])
					);
				end
				assign out_ready = out_ready_i & ((lane == 0) | result_is_vector);
				assign lane_out_valid[lane] = out_valid & ((lane == 0) | result_is_vector);
				assign local_result = (lane_out_valid[lane] ? op_result : {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}});
				assign lane_status[lane * 5+:5] = (lane_out_valid[lane] ? op_status : {5 {1'sb0}});
			end
			else begin : inactive_lane
				assign lane_out_valid[lane] = 1'b0;
				assign lane_in_ready[lane] = 1'b0;
				assign local_result = {(OpGroup == 2'd3 ? fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_conv_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane))))) : fpnew_pkg_max_fp_width(sv2v_cast_F8FCA(fpnew_pkg_get_lane_formats(Width, FpFmtConfig, sv2v_cast_32($unsigned(lane)))))) {lane_ext_bit[0]}};
				assign lane_status[lane * 5+:5] = 1'sb0;
				assign lane_busy[lane] = 1'b0;
			end
			genvar fmt;
			for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : pack_fp_result
				localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
				if (ACTIVE_FORMATS[fmt]) begin : genblk1
					assign fmt_slice_result[(fmt * Width) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((LANE + 1) * FP_WIDTH) - 1 : ((((LANE + 1) * FP_WIDTH) - 1) + ((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * FP_WIDTH) - 1) >= (LANE * FP_WIDTH) ? ((((LANE + 1) * FP_WIDTH) - 1) - (LANE * FP_WIDTH)) + 1 : ((LANE * FP_WIDTH) - (((LANE + 1) * FP_WIDTH) - 1)) + 1)] = local_result[FP_WIDTH - 1:0];
				end
			end
			if (OpGroup == 2'd3) begin : int_results_enabled
				genvar ifmt;
				for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : pack_int_result
					localparam [31:0] INT_WIDTH = fpnew_pkg_int_width(sv2v_cast_87CC5(ifmt));
					if (ACTIVE_INT_FORMATS[ifmt]) begin : genblk1
						assign ifmt_slice_result[(ifmt * Width) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((LANE + 1) * INT_WIDTH) - 1 : ((((LANE + 1) * INT_WIDTH) - 1) + ((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)) - 1)-:((((LANE + 1) * INT_WIDTH) - 1) >= (LANE * INT_WIDTH) ? ((((LANE + 1) * INT_WIDTH) - 1) - (LANE * INT_WIDTH)) + 1 : ((LANE * INT_WIDTH) - (((LANE + 1) * INT_WIDTH) - 1)) + 1)] = local_result[INT_WIDTH - 1:0];
					end
				end
			end
		end
	endgenerate
	genvar fmt;
	generate
		for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1) begin : extend_fp_result
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if ((NUM_LANES * FP_WIDTH) < Width) begin : genblk1
				assign fmt_slice_result[(fmt * Width) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? Width - 1 : ((Width - 1) + ((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)) - 1)-:((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1)] = {((Width - 1) >= (NUM_LANES * FP_WIDTH) ? ((Width - 1) - (NUM_LANES * FP_WIDTH)) + 1 : ((NUM_LANES * FP_WIDTH) - (Width - 1)) + 1) {lane_ext_bit[0]}};
			end
		end
	endgenerate
	genvar ifmt;
	generate
		for (ifmt = 0; ifmt < NUM_INT_FORMATS; ifmt = ifmt + 1) begin : int_results_disabled
			if (OpGroup != 2'd3) begin : mute_int_result
				assign ifmt_slice_result[ifmt * Width+:Width] = 1'sb0;
			end
		end
		if (OpGroup == 2'd3) begin : target_regs
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * Width) + ((NumPipeRegs * Width) - 1) : ((NumPipeRegs + 1) * Width) - 1):(0 >= NumPipeRegs ? NumPipeRegs * Width : 0)] byp_pipe_target_q;
			reg [(0 >= NumPipeRegs ? ((1 - NumPipeRegs) * 3) + ((NumPipeRegs * 3) - 1) : ((NumPipeRegs + 1) * 3) - 1):(0 >= NumPipeRegs ? NumPipeRegs * 3 : 0)] byp_pipe_aux_q;
			reg [0:NumPipeRegs] byp_pipe_valid_q;
			wire [0:NumPipeRegs] byp_pipe_ready;
			wire [Width * 1:1] sv2v_tmp_FBD8C;
			assign sv2v_tmp_FBD8C = conv_target_d;
			always @(*) byp_pipe_target_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * Width+:Width] = sv2v_tmp_FBD8C;
			wire [3:1] sv2v_tmp_A0A5D;
			assign sv2v_tmp_A0A5D = target_aux_d;
			always @(*) byp_pipe_aux_q[(0 >= NumPipeRegs ? 0 : NumPipeRegs) * 3+:3] = sv2v_tmp_A0A5D;
			wire [1:1] sv2v_tmp_49222;
			assign sv2v_tmp_49222 = in_valid_i & vectorial_op;
			always @(*) byp_pipe_valid_q[0] = sv2v_tmp_49222;
			genvar i;
			for (i = 0; i < NumPipeRegs; i = i + 1) begin : gen_bypass_pipeline
				wire reg_ena;
				assign byp_pipe_ready[i] = byp_pipe_ready[i + 1] | ~byp_pipe_valid_q[i + 1];
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						byp_pipe_valid_q[i + 1] <= 1'b0;
					else
						byp_pipe_valid_q[i + 1] <= (flush_i ? 1'b0 : (byp_pipe_ready[i] ? byp_pipe_valid_q[i] : byp_pipe_valid_q[i + 1]));
				assign reg_ena = byp_pipe_ready[i] & byp_pipe_valid_q[i];
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= 1'sb0;
					else
						byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width] <= (reg_ena ? byp_pipe_target_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * Width+:Width] : byp_pipe_target_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * Width+:Width]);
				always @(posedge clk_i or negedge rst_ni)
					if (!rst_ni)
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= 1'sb0;
					else
						byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3] <= (reg_ena ? byp_pipe_aux_q[(0 >= NumPipeRegs ? i : NumPipeRegs - i) * 3+:3] : byp_pipe_aux_q[(0 >= NumPipeRegs ? i + 1 : NumPipeRegs - (i + 1)) * 3+:3]);
			end
			assign byp_pipe_ready[NumPipeRegs] = out_ready_i & result_is_vector;
			assign conv_target_q = byp_pipe_target_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * Width+:Width];
			assign {result_vec_op, result_is_cpk} = byp_pipe_aux_q[(0 >= NumPipeRegs ? NumPipeRegs : NumPipeRegs - NumPipeRegs) * 3+:3];
		end
		else begin : no_conv
			assign {result_vec_op, result_is_cpk} = 1'sb0;
		end
	endgenerate
	assign {result_fmt_is_int, result_is_vector, result_fmt} = lane_aux[0+:AUX_BITS];
	assign result_o = (result_fmt_is_int ? ifmt_slice_result[result_fmt * Width+:Width] : fmt_slice_result[result_fmt * Width+:Width]);
	assign extension_bit_o = lane_ext_bit[0];
	assign tag_o = lane_tags[0+:3];
	assign busy_o = |lane_busy;
	assign out_valid_o = lane_out_valid[0];
	always @(*) begin : output_processing
		reg [4:0] temp_status;
		temp_status = 1'sb0;
		begin : sv2v_autoblock_12
			reg signed [31:0] i;
			for (i = 0; i < sv2v_cast_32_signed(NUM_LANES); i = i + 1)
				temp_status = temp_status | lane_status[i * 5+:5];
		end
		status_o = temp_status;
	end
endmodule
module fpnew_rounding (
	abs_value_i,
	sign_i,
	round_sticky_bits_i,
	rnd_mode_i,
	effective_subtraction_i,
	abs_rounded_o,
	sign_o,
	exact_zero_o
);
	parameter [31:0] AbsWidth = 2;
	input wire [AbsWidth - 1:0] abs_value_i;
	input wire sign_i;
	input wire [1:0] round_sticky_bits_i;
	input wire [2:0] rnd_mode_i;
	input wire effective_subtraction_i;
	output wire [AbsWidth - 1:0] abs_rounded_o;
	output wire sign_o;
	output wire exact_zero_o;
	reg round_up;
	localparam [0:0] fpnew_pkg_DONT_CARE = 1'b1;
	always @(*) begin : rounding_decision
		case (rnd_mode_i)
			3'b000:
				case (round_sticky_bits_i)
					2'b00, 2'b01: round_up = 1'b0;
					2'b10: round_up = abs_value_i[0];
					2'b11: round_up = 1'b1;
					default: round_up = fpnew_pkg_DONT_CARE;
				endcase
			3'b001: round_up = 1'b0;
			3'b010: round_up = (|round_sticky_bits_i ? sign_i : 1'b0);
			3'b011: round_up = (|round_sticky_bits_i ? ~sign_i : 1'b0);
			3'b100: round_up = round_sticky_bits_i[1];
			default: round_up = fpnew_pkg_DONT_CARE;
		endcase
	end
	assign abs_rounded_o = abs_value_i + round_up;
	assign exact_zero_o = (abs_value_i == {AbsWidth {1'sb0}}) && (round_sticky_bits_i == {2 {1'sb0}});
	assign sign_o = (exact_zero_o && effective_subtraction_i ? rnd_mode_i == 3'b010 : sign_i);
endmodule
module fpnew_top_60D59 (
	clk_i,
	rst_ni,
	operands_i,
	rnd_mode_i,
	op_i,
	op_mod_i,
	src_fmt_i,
	dst_fmt_i,
	int_fmt_i,
	vectorial_op_i,
	tag_i,
	in_valid_i,
	in_ready_o,
	flush_i,
	result_o,
	status_o,
	tag_o,
	out_valid_o,
	out_ready_i,
	busy_o
);
	localparam [31:0] fpnew_pkg_NUM_FP_FORMATS = 5;
	localparam [31:0] fpnew_pkg_NUM_INT_FORMATS = 4;
	localparam [42:0] fpnew_pkg_RV64D_Xsflt = 43'h000000207ff;
	parameter [42:0] Features = fpnew_pkg_RV64D_Xsflt;
	localparam [31:0] fpnew_pkg_NUM_OPGROUPS = 4;
	function automatic [159:0] sv2v_cast_B9240;
		input reg [159:0] inp;
		sv2v_cast_B9240 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 32) - 1:0] sv2v_cast_CDC93;
		input reg [((32'd4 * 32'd5) * 32) - 1:0] inp;
		sv2v_cast_CDC93 = inp;
	endfunction
	function automatic [((32'd4 * 32'd5) * 2) - 1:0] sv2v_cast_15FEF;
		input reg [((32'd4 * 32'd5) * 2) - 1:0] inp;
		sv2v_cast_15FEF = inp;
	endfunction
	localparam [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] fpnew_pkg_DEFAULT_NOREGS = {sv2v_cast_CDC93({fpnew_pkg_NUM_OPGROUPS {sv2v_cast_B9240(0)}}), sv2v_cast_15FEF({{fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}, {fpnew_pkg_NUM_FP_FORMATS {2'd1}}, {fpnew_pkg_NUM_FP_FORMATS {2'd2}}}), 2'd0};
	parameter [(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + ((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2)) + 1:0] Implementation = fpnew_pkg_DEFAULT_NOREGS;
	localparam [31:0] WIDTH = Features[42-:32];
	localparam [31:0] NUM_OPERANDS = 3;
	input wire clk_i;
	input wire rst_ni;
	input wire [(NUM_OPERANDS * WIDTH) - 1:0] operands_i;
	input wire [2:0] rnd_mode_i;
	localparam [31:0] fpnew_pkg_OP_BITS = 4;
	input wire [3:0] op_i;
	input wire op_mod_i;
	localparam [31:0] fpnew_pkg_FP_FORMAT_BITS = 3;
	input wire [2:0] src_fmt_i;
	input wire [2:0] dst_fmt_i;
	localparam [31:0] fpnew_pkg_INT_FORMAT_BITS = 2;
	input wire [1:0] int_fmt_i;
	input wire vectorial_op_i;
	input wire [2:0] tag_i;
	input wire in_valid_i;
	output wire in_ready_o;
	input wire flush_i;
	output wire [WIDTH - 1:0] result_o;
	output wire [4:0] status_o;
	output wire [2:0] tag_o;
	output wire out_valid_o;
	input wire out_ready_i;
	output wire busy_o;
	localparam [31:0] NUM_OPGROUPS = fpnew_pkg_NUM_OPGROUPS;
	localparam [31:0] NUM_FORMATS = fpnew_pkg_NUM_FP_FORMATS;
	wire [3:0] opgrp_in_ready;
	wire [3:0] opgrp_out_valid;
	wire [3:0] opgrp_out_ready;
	wire [3:0] opgrp_ext;
	wire [3:0] opgrp_busy;
	wire [((WIDTH + 7) >= 0 ? (4 * (WIDTH + 8)) - 1 : (4 * (1 - (WIDTH + 7))) + (WIDTH + 6)):((WIDTH + 7) >= 0 ? 0 : WIDTH + 7)] opgrp_outputs;
	wire [(NUM_FORMATS * NUM_OPERANDS) - 1:0] is_boxed;
	function automatic [3:0] sv2v_cast_A53F3;
		input reg [3:0] inp;
		sv2v_cast_A53F3 = inp;
	endfunction
	function automatic [1:0] fpnew_pkg_get_opgroup;
		input reg [3:0] op;
		case (op)
			sv2v_cast_A53F3(0), sv2v_cast_A53F3(1), sv2v_cast_A53F3(2), sv2v_cast_A53F3(3): fpnew_pkg_get_opgroup = 2'd0;
			sv2v_cast_A53F3(4), sv2v_cast_A53F3(5): fpnew_pkg_get_opgroup = 2'd1;
			sv2v_cast_A53F3(6), sv2v_cast_A53F3(7), sv2v_cast_A53F3(8), sv2v_cast_A53F3(9): fpnew_pkg_get_opgroup = 2'd2;
			sv2v_cast_A53F3(10), sv2v_cast_A53F3(11), sv2v_cast_A53F3(12), sv2v_cast_A53F3(13), sv2v_cast_A53F3(14): fpnew_pkg_get_opgroup = 2'd3;
			default: fpnew_pkg_get_opgroup = 2'd2;
		endcase
	endfunction
	assign in_ready_o = in_valid_i & opgrp_in_ready[fpnew_pkg_get_opgroup(op_i)];
	genvar fmt;
	localparam [319:0] fpnew_pkg_FP_ENCODINGS = 320'h8000000170000000b00000034000000050000000a00000005000000020000000800000007;
	function automatic [31:0] fpnew_pkg_fp_width;
		input reg [2:0] fmt;
		fpnew_pkg_fp_width = (fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 63-:32] + fpnew_pkg_FP_ENCODINGS[((4 - fmt) * 64) + 31-:32]) + 1;
	endfunction
	function automatic [2:0] sv2v_cast_0BC43;
		input reg [2:0] inp;
		sv2v_cast_0BC43 = inp;
	endfunction
	function automatic signed [31:0] sv2v_cast_32_signed;
		input reg signed [31:0] inp;
		sv2v_cast_32_signed = inp;
	endfunction
	generate
		for (fmt = 0; fmt < sv2v_cast_32_signed(NUM_FORMATS); fmt = fmt + 1) begin : gen_nanbox_check
			localparam [31:0] FP_WIDTH = fpnew_pkg_fp_width(sv2v_cast_0BC43(fmt));
			if (Features[9] && (FP_WIDTH < WIDTH)) begin : check
				genvar op;
				for (op = 0; op < sv2v_cast_32_signed(NUM_OPERANDS); op = op + 1) begin : operands
					assign is_boxed[(fmt * NUM_OPERANDS) + op] = (!vectorial_op_i ? operands_i[(op * WIDTH) + ((WIDTH - 1) >= FP_WIDTH ? WIDTH - 1 : ((WIDTH - 1) + ((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)) - 1)-:((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1)] == {((WIDTH - 1) >= FP_WIDTH ? ((WIDTH - 1) - FP_WIDTH) + 1 : (FP_WIDTH - (WIDTH - 1)) + 1) * 1 {1'sb1}} : 1'b1);
				end
			end
			else begin : no_check
				assign is_boxed[fmt * NUM_OPERANDS+:NUM_OPERANDS] = 1'sb1;
			end
		end
	endgenerate
	genvar opgrp;
	function automatic [31:0] fpnew_pkg_num_operands;
		input reg [1:0] grp;
		case (grp)
			2'd0: fpnew_pkg_num_operands = 3;
			2'd1: fpnew_pkg_num_operands = 2;
			2'd2: fpnew_pkg_num_operands = 2;
			2'd3: fpnew_pkg_num_operands = 3;
			default: fpnew_pkg_num_operands = 0;
		endcase
	endfunction
	function automatic [1:0] sv2v_cast_2;
		input reg [1:0] inp;
		sv2v_cast_2 = inp;
	endfunction
	generate
		for (opgrp = 0; opgrp < sv2v_cast_32_signed(NUM_OPGROUPS); opgrp = opgrp + 1) begin : gen_operation_groups
			localparam [31:0] NUM_OPS = fpnew_pkg_num_operands(sv2v_cast_2(opgrp));
			wire in_valid;
			reg [(NUM_FORMATS * NUM_OPS) - 1:0] input_boxed;
			assign in_valid = in_valid_i & (fpnew_pkg_get_opgroup(op_i) == sv2v_cast_2(opgrp));
			always @(*) begin : slice_inputs
				begin : sv2v_autoblock_1
					reg [31:0] fmt;
					for (fmt = 0; fmt < NUM_FORMATS; fmt = fmt + 1)
						input_boxed[fmt * fpnew_pkg_num_operands(sv2v_cast_2(opgrp))+:fpnew_pkg_num_operands(sv2v_cast_2(opgrp))] = is_boxed[(fmt * NUM_OPERANDS) + (NUM_OPS - 1)-:NUM_OPS];
				end
			end
			fpnew_opgroup_block_AC56A #(
				.OpGroup(sv2v_cast_2(opgrp)),
				.Width(WIDTH),
				.EnableVectors(Features[10]),
				.FpFmtMask(Features[8-:5]),
				.IntFmtMask(Features[3-:fpnew_pkg_NUM_INT_FORMATS]),
				.FmtPipeRegs(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) + (((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1)) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 32) - 1) - (32 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:160]),
				.FmtUnitTypes(Implementation[(((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) + 1) - ((((fpnew_pkg_NUM_OPGROUPS * fpnew_pkg_NUM_FP_FORMATS) * 2) - 1) - (2 * ((3 - opgrp) * fpnew_pkg_NUM_FP_FORMATS)))+:10]),
				.PipeConfig(Implementation[1-:2])
			) i_opgroup_block(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.operands_i(operands_i[WIDTH * ((NUM_OPS - 1) - (NUM_OPS - 1))+:WIDTH * NUM_OPS]),
				.is_boxed_i(input_boxed),
				.rnd_mode_i(rnd_mode_i),
				.op_i(op_i),
				.op_mod_i(op_mod_i),
				.src_fmt_i(src_fmt_i),
				.dst_fmt_i(dst_fmt_i),
				.int_fmt_i(int_fmt_i),
				.vectorial_op_i(vectorial_op_i),
				.tag_i(tag_i),
				.in_valid_i(in_valid),
				.in_ready_o(opgrp_in_ready[opgrp]),
				.flush_i(flush_i),
				.result_o(opgrp_outputs[((WIDTH + 7) >= 0 ? (opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? WIDTH + 7 : (WIDTH + 7) - (WIDTH + 7)) : (((opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? WIDTH + 7 : (WIDTH + 7) - (WIDTH + 7))) + ((WIDTH + 7) >= 8 ? WIDTH + 0 : 9 - (WIDTH + 7))) - 1)-:((WIDTH + 7) >= 8 ? WIDTH + 0 : 9 - (WIDTH + 7))]),
				.status_o(opgrp_outputs[((WIDTH + 7) >= 0 ? (opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? 7 : WIDTH + 0) : ((opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? 7 : WIDTH + 0)) + 4)-:5]),
				.extension_bit_o(opgrp_ext[opgrp]),
				.tag_o(opgrp_outputs[((WIDTH + 7) >= 0 ? (opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? 2 : WIDTH + 5) : ((opgrp * ((WIDTH + 7) >= 0 ? WIDTH + 8 : 1 - (WIDTH + 7))) + ((WIDTH + 7) >= 0 ? 2 : WIDTH + 5)) + 2)-:3]),
				.out_valid_o(opgrp_out_valid[opgrp]),
				.out_ready_i(opgrp_out_ready[opgrp]),
				.busy_o(opgrp_busy[opgrp])
			);
		end
	endgenerate
	wire [WIDTH + 7:0] arbiter_output;
	localparam [31:0] sv2v_uu_i_arbiter_NumIn = NUM_OPGROUPS;
	localparam [1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_79FBE_62ECB #(
		.DataType_WIDTH(WIDTH),
		.NumIn(NUM_OPGROUPS),
		.AxiVldRdy(1'b1)
	) i_arbiter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
		.req_i(opgrp_out_valid),
		.gnt_o(opgrp_out_ready),
		.data_i(opgrp_outputs),
		.gnt_i(out_ready_i),
		.req_o(out_valid_o),
		.data_o(arbiter_output),
		.idx_o()
	);
	assign result_o = arbiter_output[WIDTH + 7-:((WIDTH + 7) >= 8 ? WIDTH + 0 : 9 - (WIDTH + 7))];
	assign status_o = arbiter_output[7-:5];
	assign tag_o = arbiter_output[2-:3];
	assign busy_o = |opgrp_busy;
endmodule
module control_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Numerator_DI,
	Exp_num_DI,
	Denominator_DI,
	Exp_den_DI,
	Div_start_dly_SO,
	Sqrt_start_dly_SO,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_result_prenorm_DO,
	Exp_result_prenorm_DO
);
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire Div_start_SI;
	input wire Sqrt_start_SI;
	input wire Start_SI;
	input wire Kill_SI;
	input wire Special_case_SBI;
	input wire Special_case_dly_SBI;
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	input wire [1:0] Format_sel_SI;
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Numerator_DI;
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_num_DI;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Denominator_DI;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_den_DI;
	output wire Div_start_dly_SO;
	output wire Sqrt_start_dly_SO;
	output reg Div_enable_SO;
	output reg Sqrt_enable_SO;
	output wire Full_precision_SO;
	output wire FP32_SO;
	output wire FP64_SO;
	output wire FP16_SO;
	output wire FP16ALT_SO;
	output reg Ready_SO;
	output reg Done_SO;
	output reg [56:0] Mant_result_prenorm_DO;
	output wire [12:0] Exp_result_prenorm_DO;
	reg [57:0] Partial_remainder_DN;
	reg [57:0] Partial_remainder_DP;
	reg [56:0] Quotient_DP;
	wire [53:0] Numerator_se_D;
	wire [53:0] Denominator_se_D;
	reg [53:0] Denominator_se_DB;
	assign Numerator_se_D = {1'b0, Numerator_DI};
	assign Denominator_se_D = {1'b0, Denominator_DI};
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	always @(*)
		if (FP32_SO)
			Denominator_se_DB = {~Denominator_se_D[53:29], {29 {1'b0}}};
		else if (FP64_SO)
			Denominator_se_DB = ~Denominator_se_D;
		else if (FP16_SO)
			Denominator_se_DB = {~Denominator_se_D[53:42], {42 {1'b0}}};
		else
			Denominator_se_DB = {~Denominator_se_D[53:45], {45 {1'b0}}};
	wire [53:0] Mant_D_sqrt_Norm;
	assign Mant_D_sqrt_Norm = (Exp_num_DI[0] ? {1'b0, Numerator_DI} : {Numerator_DI, 1'b0});
	reg [1:0] Format_sel_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Format_sel_S <= 'b0;
		else if (Start_SI && Ready_SO)
			Format_sel_S <= Format_sel_SI;
		else
			Format_sel_S <= Format_sel_S;
	assign FP32_SO = Format_sel_S == 2'b00;
	assign FP64_SO = Format_sel_S == 2'b01;
	assign FP16_SO = Format_sel_S == 2'b10;
	assign FP16ALT_SO = Format_sel_S == 2'b11;
	reg [5:0] Precision_ctl_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Precision_ctl_S <= 'b0;
		else if (Start_SI && Ready_SO)
			Precision_ctl_S <= Precision_ctl_SI;
		else
			Precision_ctl_S <= Precision_ctl_S;
	assign Full_precision_SO = Precision_ctl_S == 6'h00;
	reg [5:0] State_ctl_S;
	wire [5:0] State_Two_iteration_unit_S;
	wire [5:0] State_Four_iteration_unit_S;
	assign State_Two_iteration_unit_S = Precision_ctl_S[5:1];
	assign State_Four_iteration_unit_S = Precision_ctl_S[5:2];
	localparam defs_div_sqrt_mvp_Iteration_unit_num_S = 2'b10;
	always @(*)
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				case (Format_sel_S)
					2'b00:
						if (Full_precision_SO)
							State_ctl_S = 6'h1b;
						else
							State_ctl_S = Precision_ctl_S;
					2'b01:
						if (Full_precision_SO)
							State_ctl_S = 6'h38;
						else
							State_ctl_S = Precision_ctl_S;
					2'b10:
						if (Full_precision_SO)
							State_ctl_S = 6'h0e;
						else
							State_ctl_S = Precision_ctl_S;
					2'b11:
						if (Full_precision_SO)
							State_ctl_S = 6'h0b;
						else
							State_ctl_S = Precision_ctl_S;
				endcase
			2'b01:
				case (Format_sel_S)
					2'b00:
						if (Full_precision_SO)
							State_ctl_S = 6'h0d;
						else
							State_ctl_S = State_Two_iteration_unit_S;
					2'b01:
						if (Full_precision_SO)
							State_ctl_S = 6'h1b;
						else
							State_ctl_S = State_Two_iteration_unit_S;
					2'b10:
						if (Full_precision_SO)
							State_ctl_S = 6'h06;
						else
							State_ctl_S = State_Two_iteration_unit_S;
					2'b11:
						if (Full_precision_SO)
							State_ctl_S = 6'h05;
						else
							State_ctl_S = State_Two_iteration_unit_S;
				endcase
			2'b10:
				case (Format_sel_S)
					2'b00:
						case (Precision_ctl_S)
							6'h00: State_ctl_S = 6'h08;
							6'h06, 6'h07, 6'h08: State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b: State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e: State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11: State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14: State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17: State_ctl_S = 6'h07;
							default: State_ctl_S = 6'h08;
						endcase
					2'b01:
						case (Precision_ctl_S)
							6'h00: State_ctl_S = 6'h12;
							6'h06, 6'h07, 6'h08: State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b: State_ctl_S = 6'h03;
							6'h0c, 6'h0d, 6'h0e: State_ctl_S = 6'h04;
							6'h0f, 6'h10, 6'h11: State_ctl_S = 6'h05;
							6'h12, 6'h13, 6'h14: State_ctl_S = 6'h06;
							6'h15, 6'h16, 6'h17: State_ctl_S = 6'h07;
							6'h18, 6'h19, 6'h1a: State_ctl_S = 6'h08;
							6'h1b, 6'h1c, 6'h1d: State_ctl_S = 6'h09;
							6'h1e, 6'h1f, 6'h20: State_ctl_S = 6'h0a;
							6'h21, 6'h22, 6'h23: State_ctl_S = 6'h0b;
							6'h24, 6'h25, 6'h26: State_ctl_S = 6'h0c;
							6'h27, 6'h28, 6'h29: State_ctl_S = 6'h0d;
							6'h2a, 6'h2b, 6'h2c: State_ctl_S = 6'h0e;
							6'h2d, 6'h2e, 6'h2f: State_ctl_S = 6'h0f;
							6'h30, 6'h31, 6'h32: State_ctl_S = 6'h10;
							6'h33, 6'h34, 6'h35: State_ctl_S = 6'h11;
							default: State_ctl_S = 6'h12;
						endcase
					2'b10:
						case (Precision_ctl_S)
							6'h00: State_ctl_S = 6'h04;
							6'h06, 6'h07, 6'h08: State_ctl_S = 6'h02;
							6'h09, 6'h0a, 6'h0b: State_ctl_S = 6'h03;
							default: State_ctl_S = 6'h04;
						endcase
					2'b11:
						case (Precision_ctl_S)
							6'h00: State_ctl_S = 6'h03;
							6'h06, 6'h07, 6'h08: State_ctl_S = 6'h02;
							default: State_ctl_S = 6'h03;
						endcase
				endcase
			2'b11:
				case (Format_sel_S)
					2'b00:
						if (Full_precision_SO)
							State_ctl_S = 6'h06;
						else
							State_ctl_S = State_Four_iteration_unit_S;
					2'b01:
						if (Full_precision_SO)
							State_ctl_S = 6'h0d;
						else
							State_ctl_S = State_Four_iteration_unit_S;
					2'b10:
						if (Full_precision_SO)
							State_ctl_S = 6'h03;
						else
							State_ctl_S = State_Four_iteration_unit_S;
					2'b11:
						if (Full_precision_SO)
							State_ctl_S = 6'h02;
						else
							State_ctl_S = State_Four_iteration_unit_S;
				endcase
		endcase
	reg Div_start_dly_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Div_start_dly_S <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			Div_start_dly_S <= 1'b1;
		else
			Div_start_dly_S <= 1'b0;
	assign Div_start_dly_SO = Div_start_dly_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Div_enable_SO <= 1'b0;
		else if (Kill_SI)
			Div_enable_SO <= 1'b0;
		else if (Div_start_SI && Ready_SO)
			Div_enable_SO <= 1'b1;
		else if (Done_SO)
			Div_enable_SO <= 1'b0;
		else
			Div_enable_SO <= Div_enable_SO;
	reg Sqrt_start_dly_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Sqrt_start_dly_S <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			Sqrt_start_dly_S <= 1'b1;
		else
			Sqrt_start_dly_S <= 1'b0;
	assign Sqrt_start_dly_SO = Sqrt_start_dly_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Sqrt_enable_SO <= 1'b0;
		else if (Kill_SI)
			Sqrt_enable_SO <= 1'b0;
		else if (Sqrt_start_SI && Ready_SO)
			Sqrt_enable_SO <= 1'b1;
		else if (Done_SO)
			Sqrt_enable_SO <= 1'b0;
		else
			Sqrt_enable_SO <= Sqrt_enable_SO;
	reg [5:0] Crtl_cnt_S;
	wire Start_dly_S;
	assign Start_dly_S = Div_start_dly_S | Sqrt_start_dly_S;
	wire Fsm_enable_S;
	assign Fsm_enable_S = ((Start_dly_S | |Crtl_cnt_S) && ~Kill_SI) && Special_case_dly_SBI;
	wire Final_state_S;
	assign Final_state_S = Crtl_cnt_S == State_ctl_S;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Crtl_cnt_S <= 1'sb0;
		else if (Final_state_S | Kill_SI)
			Crtl_cnt_S <= 1'sb0;
		else if (Fsm_enable_S)
			Crtl_cnt_S <= Crtl_cnt_S + 1;
		else
			Crtl_cnt_S <= 1'sb0;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Done_SO <= 1'b0;
		else if (Start_SI && Ready_SO) begin
			if (~Special_case_SBI)
				Done_SO <= 1'b1;
			else
				Done_SO <= 1'b0;
		end
		else if (Final_state_S)
			Done_SO <= 1'b1;
		else
			Done_SO <= 1'b0;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Ready_SO <= 1'b1;
		else if (Start_SI && Ready_SO) begin
			if (~Special_case_SBI)
				Ready_SO <= 1'b1;
			else
				Ready_SO <= 1'b0;
		end
		else if (Final_state_S | Kill_SI)
			Ready_SO <= 1'b1;
		else
			Ready_SO <= Ready_SO;
	wire Qcnt_one_0;
	wire Qcnt_one_1;
	wire [1:0] Qcnt_one_2;
	wire [2:0] Qcnt_one_3;
	wire [3:0] Qcnt_one_4;
	wire [4:0] Qcnt_one_5;
	wire [5:0] Qcnt_one_6;
	wire [6:0] Qcnt_one_7;
	wire [7:0] Qcnt_one_8;
	wire [8:0] Qcnt_one_9;
	wire [9:0] Qcnt_one_10;
	wire [10:0] Qcnt_one_11;
	wire [11:0] Qcnt_one_12;
	wire [12:0] Qcnt_one_13;
	wire [13:0] Qcnt_one_14;
	wire [14:0] Qcnt_one_15;
	wire [15:0] Qcnt_one_16;
	wire [16:0] Qcnt_one_17;
	wire [17:0] Qcnt_one_18;
	wire [18:0] Qcnt_one_19;
	wire [19:0] Qcnt_one_20;
	wire [20:0] Qcnt_one_21;
	wire [21:0] Qcnt_one_22;
	wire [22:0] Qcnt_one_23;
	wire [23:0] Qcnt_one_24;
	wire [24:0] Qcnt_one_25;
	wire [25:0] Qcnt_one_26;
	wire [26:0] Qcnt_one_27;
	wire [27:0] Qcnt_one_28;
	wire [28:0] Qcnt_one_29;
	wire [29:0] Qcnt_one_30;
	wire [30:0] Qcnt_one_31;
	wire [31:0] Qcnt_one_32;
	wire [32:0] Qcnt_one_33;
	wire [33:0] Qcnt_one_34;
	wire [34:0] Qcnt_one_35;
	wire [35:0] Qcnt_one_36;
	wire [36:0] Qcnt_one_37;
	wire [37:0] Qcnt_one_38;
	wire [38:0] Qcnt_one_39;
	wire [39:0] Qcnt_one_40;
	wire [40:0] Qcnt_one_41;
	wire [41:0] Qcnt_one_42;
	wire [42:0] Qcnt_one_43;
	wire [43:0] Qcnt_one_44;
	wire [44:0] Qcnt_one_45;
	wire [45:0] Qcnt_one_46;
	wire [46:0] Qcnt_one_47;
	wire [47:0] Qcnt_one_48;
	wire [48:0] Qcnt_one_49;
	wire [49:0] Qcnt_one_50;
	wire [50:0] Qcnt_one_51;
	wire [51:0] Qcnt_one_52;
	wire [52:0] Qcnt_one_53;
	wire [53:0] Qcnt_one_54;
	wire [54:0] Qcnt_one_55;
	wire [55:0] Qcnt_one_56;
	wire [56:0] Qcnt_one_57;
	wire [57:0] Qcnt_one_58;
	wire [58:0] Qcnt_one_59;
	wire [59:0] Qcnt_one_60;
	wire [1:0] Qcnt_two_0;
	wire [2:0] Qcnt_two_1;
	wire [4:0] Qcnt_two_2;
	wire [6:0] Qcnt_two_3;
	wire [8:0] Qcnt_two_4;
	wire [10:0] Qcnt_two_5;
	wire [12:0] Qcnt_two_6;
	wire [14:0] Qcnt_two_7;
	wire [16:0] Qcnt_two_8;
	wire [18:0] Qcnt_two_9;
	wire [20:0] Qcnt_two_10;
	wire [22:0] Qcnt_two_11;
	wire [24:0] Qcnt_two_12;
	wire [26:0] Qcnt_two_13;
	wire [28:0] Qcnt_two_14;
	wire [30:0] Qcnt_two_15;
	wire [32:0] Qcnt_two_16;
	wire [34:0] Qcnt_two_17;
	wire [36:0] Qcnt_two_18;
	wire [38:0] Qcnt_two_19;
	wire [40:0] Qcnt_two_20;
	wire [42:0] Qcnt_two_21;
	wire [44:0] Qcnt_two_22;
	wire [46:0] Qcnt_two_23;
	wire [48:0] Qcnt_two_24;
	wire [50:0] Qcnt_two_25;
	wire [52:0] Qcnt_two_26;
	wire [54:0] Qcnt_two_27;
	wire [56:0] Qcnt_two_28;
	wire [2:0] Qcnt_three_0;
	wire [4:0] Qcnt_three_1;
	wire [7:0] Qcnt_three_2;
	wire [10:0] Qcnt_three_3;
	wire [13:0] Qcnt_three_4;
	wire [16:0] Qcnt_three_5;
	wire [19:0] Qcnt_three_6;
	wire [22:0] Qcnt_three_7;
	wire [25:0] Qcnt_three_8;
	wire [28:0] Qcnt_three_9;
	wire [31:0] Qcnt_three_10;
	wire [34:0] Qcnt_three_11;
	wire [37:0] Qcnt_three_12;
	wire [40:0] Qcnt_three_13;
	wire [43:0] Qcnt_three_14;
	wire [46:0] Qcnt_three_15;
	wire [49:0] Qcnt_three_16;
	wire [52:0] Qcnt_three_17;
	wire [55:0] Qcnt_three_18;
	wire [58:0] Qcnt_three_19;
	wire [61:0] Qcnt_three_20;
	wire [3:0] Qcnt_four_0;
	wire [6:0] Qcnt_four_1;
	wire [10:0] Qcnt_four_2;
	wire [14:0] Qcnt_four_3;
	wire [18:0] Qcnt_four_4;
	wire [22:0] Qcnt_four_5;
	wire [26:0] Qcnt_four_6;
	wire [30:0] Qcnt_four_7;
	wire [34:0] Qcnt_four_8;
	wire [38:0] Qcnt_four_9;
	wire [42:0] Qcnt_four_10;
	wire [46:0] Qcnt_four_11;
	wire [50:0] Qcnt_four_12;
	wire [54:0] Qcnt_four_13;
	wire [58:0] Qcnt_four_14;
	wire [57:0] Sqrt_R0;
	reg [57:0] Sqrt_Q0;
	reg [57:0] Q_sqrt0;
	reg [57:0] Q_sqrt_com_0;
	wire [57:0] Sqrt_R1;
	reg [57:0] Sqrt_Q1;
	reg [57:0] Q_sqrt1;
	reg [57:0] Q_sqrt_com_1;
	wire [57:0] Sqrt_R2;
	reg [57:0] Sqrt_Q2;
	reg [57:0] Q_sqrt2;
	reg [57:0] Q_sqrt_com_2;
	wire [57:0] Sqrt_R3;
	reg [57:0] Sqrt_Q3;
	reg [57:0] Q_sqrt3;
	reg [57:0] Q_sqrt_com_3;
	wire [57:0] Sqrt_R4;
	reg [1:0] Sqrt_DI [3:0];
	wire [1:0] Sqrt_DO [3:0];
	wire Sqrt_carry_DO;
	wire [57:0] Iteration_cell_a_D [3:0];
	wire [57:0] Iteration_cell_b_D [3:0];
	wire [57:0] Iteration_cell_a_BMASK_D [3:0];
	wire [57:0] Iteration_cell_b_BMASK_D [3:0];
	wire Iteration_cell_carry_D [3:0];
	wire [57:0] Iteration_cell_sum_D [3:0];
	wire [57:0] Iteration_cell_sum_AMASK_D [3:0];
	reg [3:0] Sqrt_quotinent_S;
	always @(*)
		case (Format_sel_S)
			2'b00: begin
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][28], ~Iteration_cell_sum_AMASK_D[1][28], ~Iteration_cell_sum_AMASK_D[2][28], ~Iteration_cell_sum_AMASK_D[3][28]};
				Q_sqrt_com_0 = {{29 {1'b0}}, ~Q_sqrt0[28:0]};
				Q_sqrt_com_1 = {{29 {1'b0}}, ~Q_sqrt1[28:0]};
				Q_sqrt_com_2 = {{29 {1'b0}}, ~Q_sqrt2[28:0]};
				Q_sqrt_com_3 = {{29 {1'b0}}, ~Q_sqrt3[28:0]};
			end
			2'b01: begin
				Sqrt_quotinent_S = {Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]};
				Q_sqrt_com_0 = ~Q_sqrt0;
				Q_sqrt_com_1 = ~Q_sqrt1;
				Q_sqrt_com_2 = ~Q_sqrt2;
				Q_sqrt_com_3 = ~Q_sqrt3;
			end
			2'b10: begin
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][15], ~Iteration_cell_sum_AMASK_D[1][15], ~Iteration_cell_sum_AMASK_D[2][15], ~Iteration_cell_sum_AMASK_D[3][15]};
				Q_sqrt_com_0 = {{42 {1'b0}}, ~Q_sqrt0[15:0]};
				Q_sqrt_com_1 = {{42 {1'b0}}, ~Q_sqrt1[15:0]};
				Q_sqrt_com_2 = {{42 {1'b0}}, ~Q_sqrt2[15:0]};
				Q_sqrt_com_3 = {{42 {1'b0}}, ~Q_sqrt3[15:0]};
			end
			2'b11: begin
				Sqrt_quotinent_S = {~Iteration_cell_sum_AMASK_D[0][12], ~Iteration_cell_sum_AMASK_D[1][12], ~Iteration_cell_sum_AMASK_D[2][12], ~Iteration_cell_sum_AMASK_D[3][12]};
				Q_sqrt_com_0 = {{45 {1'b0}}, ~Q_sqrt0[12:0]};
				Q_sqrt_com_1 = {{45 {1'b0}}, ~Q_sqrt1[12:0]};
				Q_sqrt_com_2 = {{45 {1'b0}}, ~Q_sqrt2[12:0]};
				Q_sqrt_com_3 = {{45 {1'b0}}, ~Q_sqrt3[12:0]};
			end
		endcase
	assign Qcnt_one_0 = 1'b0;
	assign Qcnt_one_1 = {Quotient_DP[0]};
	assign Qcnt_one_2 = {Quotient_DP[1:0]};
	assign Qcnt_one_3 = {Quotient_DP[2:0]};
	assign Qcnt_one_4 = {Quotient_DP[3:0]};
	assign Qcnt_one_5 = {Quotient_DP[4:0]};
	assign Qcnt_one_6 = {Quotient_DP[5:0]};
	assign Qcnt_one_7 = {Quotient_DP[6:0]};
	assign Qcnt_one_8 = {Quotient_DP[7:0]};
	assign Qcnt_one_9 = {Quotient_DP[8:0]};
	assign Qcnt_one_10 = {Quotient_DP[9:0]};
	assign Qcnt_one_11 = {Quotient_DP[10:0]};
	assign Qcnt_one_12 = {Quotient_DP[11:0]};
	assign Qcnt_one_13 = {Quotient_DP[12:0]};
	assign Qcnt_one_14 = {Quotient_DP[13:0]};
	assign Qcnt_one_15 = {Quotient_DP[14:0]};
	assign Qcnt_one_16 = {Quotient_DP[15:0]};
	assign Qcnt_one_17 = {Quotient_DP[16:0]};
	assign Qcnt_one_18 = {Quotient_DP[17:0]};
	assign Qcnt_one_19 = {Quotient_DP[18:0]};
	assign Qcnt_one_20 = {Quotient_DP[19:0]};
	assign Qcnt_one_21 = {Quotient_DP[20:0]};
	assign Qcnt_one_22 = {Quotient_DP[21:0]};
	assign Qcnt_one_23 = {Quotient_DP[22:0]};
	assign Qcnt_one_24 = {Quotient_DP[23:0]};
	assign Qcnt_one_25 = {Quotient_DP[24:0]};
	assign Qcnt_one_26 = {Quotient_DP[25:0]};
	assign Qcnt_one_27 = {Quotient_DP[26:0]};
	assign Qcnt_one_28 = {Quotient_DP[27:0]};
	assign Qcnt_one_29 = {Quotient_DP[28:0]};
	assign Qcnt_one_30 = {Quotient_DP[29:0]};
	assign Qcnt_one_31 = {Quotient_DP[30:0]};
	assign Qcnt_one_32 = {Quotient_DP[31:0]};
	assign Qcnt_one_33 = {Quotient_DP[32:0]};
	assign Qcnt_one_34 = {Quotient_DP[33:0]};
	assign Qcnt_one_35 = {Quotient_DP[34:0]};
	assign Qcnt_one_36 = {Quotient_DP[35:0]};
	assign Qcnt_one_37 = {Quotient_DP[36:0]};
	assign Qcnt_one_38 = {Quotient_DP[37:0]};
	assign Qcnt_one_39 = {Quotient_DP[38:0]};
	assign Qcnt_one_40 = {Quotient_DP[39:0]};
	assign Qcnt_one_41 = {Quotient_DP[40:0]};
	assign Qcnt_one_42 = {Quotient_DP[41:0]};
	assign Qcnt_one_43 = {Quotient_DP[42:0]};
	assign Qcnt_one_44 = {Quotient_DP[43:0]};
	assign Qcnt_one_45 = {Quotient_DP[44:0]};
	assign Qcnt_one_46 = {Quotient_DP[45:0]};
	assign Qcnt_one_47 = {Quotient_DP[46:0]};
	assign Qcnt_one_48 = {Quotient_DP[47:0]};
	assign Qcnt_one_49 = {Quotient_DP[48:0]};
	assign Qcnt_one_50 = {Quotient_DP[49:0]};
	assign Qcnt_one_51 = {Quotient_DP[50:0]};
	assign Qcnt_one_52 = {Quotient_DP[51:0]};
	assign Qcnt_one_53 = {Quotient_DP[52:0]};
	assign Qcnt_one_54 = {Quotient_DP[53:0]};
	assign Qcnt_one_55 = {Quotient_DP[54:0]};
	assign Qcnt_one_56 = {Quotient_DP[55:0]};
	assign Qcnt_one_57 = {Quotient_DP[56:0]};
	assign Qcnt_two_0 = {1'b0, Sqrt_quotinent_S[3]};
	assign Qcnt_two_1 = {Quotient_DP[1:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_2 = {Quotient_DP[3:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_3 = {Quotient_DP[5:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_4 = {Quotient_DP[7:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_5 = {Quotient_DP[9:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_6 = {Quotient_DP[11:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_7 = {Quotient_DP[13:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_8 = {Quotient_DP[15:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_9 = {Quotient_DP[17:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_10 = {Quotient_DP[19:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_11 = {Quotient_DP[21:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_12 = {Quotient_DP[23:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_13 = {Quotient_DP[25:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_14 = {Quotient_DP[27:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_15 = {Quotient_DP[29:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_16 = {Quotient_DP[31:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_17 = {Quotient_DP[33:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_18 = {Quotient_DP[35:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_19 = {Quotient_DP[37:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_20 = {Quotient_DP[39:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_21 = {Quotient_DP[41:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_22 = {Quotient_DP[43:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_23 = {Quotient_DP[45:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_24 = {Quotient_DP[47:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_25 = {Quotient_DP[49:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_26 = {Quotient_DP[51:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_27 = {Quotient_DP[53:0], Sqrt_quotinent_S[3]};
	assign Qcnt_two_28 = {Quotient_DP[55:0], Sqrt_quotinent_S[3]};
	assign Qcnt_three_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_1 = {Quotient_DP[2:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_2 = {Quotient_DP[5:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_3 = {Quotient_DP[8:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_4 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_5 = {Quotient_DP[14:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_6 = {Quotient_DP[17:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_7 = {Quotient_DP[20:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_8 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_9 = {Quotient_DP[26:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_10 = {Quotient_DP[29:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_11 = {Quotient_DP[32:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_12 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_13 = {Quotient_DP[38:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_14 = {Quotient_DP[41:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_15 = {Quotient_DP[44:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_16 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_17 = {Quotient_DP[50:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_18 = {Quotient_DP[53:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_three_19 = {Quotient_DP[56:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2]};
	assign Qcnt_four_0 = {1'b0, Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_1 = {Quotient_DP[3:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_2 = {Quotient_DP[7:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_3 = {Quotient_DP[11:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_4 = {Quotient_DP[15:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_5 = {Quotient_DP[19:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_6 = {Quotient_DP[23:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_7 = {Quotient_DP[27:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_8 = {Quotient_DP[31:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_9 = {Quotient_DP[35:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_10 = {Quotient_DP[39:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_11 = {Quotient_DP[43:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_12 = {Quotient_DP[47:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_13 = {Quotient_DP[51:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	assign Qcnt_four_14 = {Quotient_DP[55:0], Sqrt_quotinent_S[3], Sqrt_quotinent_S[2], Sqrt_quotinent_S[1]};
	always @(*)
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				case (Crtl_cnt_S)
					6'b000000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_0};
						Sqrt_Q0 = Q_sqrt_com_0;
					end
					6'b000001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_one_1};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_one_2};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						Q_sqrt0 = {{55 {1'b0}}, Qcnt_one_3};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_one_4};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[43:42];
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_one_5};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_one_6};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b000111: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[39:38];
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_one_7};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_one_8};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_one_9};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_one_10};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[31:30];
						Q_sqrt0 = {{47 {1'b0}}, Qcnt_one_11};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_one_12};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[27:26];
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_one_13};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_one_14};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b001111: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						Q_sqrt0 = {{43 {1'b0}}, Qcnt_one_15};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_one_16};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[19:18];
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_one_17};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_one_18};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[15:14];
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_one_19};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_one_20};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_one_21};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_one_22};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b010111: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[7:6];
						Q_sqrt0 = {{35 {1'b0}}, Qcnt_one_23};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_one_24};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[3:2];
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_one_25};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_one_26};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{31 {1'b0}}, Qcnt_one_27};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_one_28};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_one_29};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_one_30};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b011111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_one_31};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_one_32};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_one_33};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_one_34};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{23 {1'b0}}, Qcnt_one_35};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_one_36};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_one_37};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_one_38};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b100111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{19 {1'b0}}, Qcnt_one_39};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_one_40};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_one_41};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_one_42};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_one_43};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_one_44};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_one_45};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_one_46};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b101111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{11 {1'b0}}, Qcnt_one_47};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_one_48};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_one_49};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_one_50};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{7 {1'b0}}, Qcnt_one_51};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_one_52};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_one_53};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_one_54};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b110111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_one_55};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					6'b111000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_one_56};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
					end
					default: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = 1'sb0;
						Sqrt_Q0 = 1'sb0;
					end
				endcase
			2'b01:
				case (Crtl_cnt_S)
					6'b000000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt0 = {{56 {1'b0}}, Qcnt_two_1[2:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[47:46];
						Q_sqrt1 = {{55 {1'b0}}, Qcnt_two_1[2:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_two_2[4:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_two_2[4:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						Q_sqrt0 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_two_3[6:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						Q_sqrt1 = {{51 {1'b0}}, Qcnt_two_3[6:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						Q_sqrt0 = {{50 {1'b0}}, Qcnt_two_4[8:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						Q_sqrt1 = {{49 {1'b0}}, Qcnt_two_4[8:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[33:32];
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_two_5[10:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[31:30];
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_two_5[10:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						Q_sqrt0 = {{46 {1'b0}}, Qcnt_two_6[12:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						Q_sqrt1 = {{45 {1'b0}}, Qcnt_two_6[12:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b000111: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[25:24];
						Q_sqrt0 = {{44 {1'b0}}, Qcnt_two_7[14:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[23:22];
						Q_sqrt1 = {{43 {1'b0}}, Qcnt_two_7[14:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_two_8[16:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_two_8[16:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						Q_sqrt0 = {{40 {1'b0}}, Qcnt_two_9[18:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						Q_sqrt1 = {{39 {1'b0}}, Qcnt_two_9[18:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						Q_sqrt0 = {{38 {1'b0}}, Qcnt_two_10[20:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						Q_sqrt1 = {{37 {1'b0}}, Qcnt_two_10[20:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[9:8];
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_two_11[22:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[7:6];
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_two_11[22:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						Q_sqrt0 = {{34 {1'b0}}, Qcnt_two_12[24:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						Q_sqrt1 = {{33 {1'b0}}, Qcnt_two_12[24:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[1:0];
						Q_sqrt0 = {{32 {1'b0}}, Qcnt_two_13[26:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{31 {1'b0}}, Qcnt_two_13[26:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_two_14[28:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_two_14[28:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b001111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{28 {1'b0}}, Qcnt_two_15[30:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{27 {1'b0}}, Qcnt_two_15[30:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{26 {1'b0}}, Qcnt_two_16[32:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{25 {1'b0}}, Qcnt_two_16[32:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_two_17[34:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_two_17[34:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{22 {1'b0}}, Qcnt_two_18[36:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{21 {1'b0}}, Qcnt_two_18[36:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{20 {1'b0}}, Qcnt_two_19[38:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{19 {1'b0}}, Qcnt_two_19[38:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_two_20[40:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_two_20[40:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{16 {1'b0}}, Qcnt_two_21[42:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{15 {1'b0}}, Qcnt_two_21[42:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{14 {1'b0}}, Qcnt_two_22[44:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{13 {1'b0}}, Qcnt_two_22[44:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b010111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_two_23[46:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_two_23[46:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{10 {1'b0}}, Qcnt_two_24[48:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{9 {1'b0}}, Qcnt_two_24[48:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{8 {1'b0}}, Qcnt_two_25[50:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{7 {1'b0}}, Qcnt_two_25[50:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_two_26[52:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_two_26[52:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{4 {1'b0}}, Qcnt_two_27[54:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{3 {1'b0}}, Qcnt_two_27[54:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					6'b011100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{2 {1'b0}}, Qcnt_two_28[56:1]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {1'b0, Qcnt_two_28[56:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
					default: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_two_0[1]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_two_0[1:0]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
					end
				endcase
			2'b10:
				case (Crtl_cnt_S)
					6'b000000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[47:46];
						Q_sqrt0 = {{54 {1'b0}}, Qcnt_three_1[4:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[45:44];
						Q_sqrt1 = {{53 {1'b0}}, Qcnt_three_1[4:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[43:42];
						Q_sqrt2 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_three_1[4:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[41:40];
						Q_sqrt0 = {{51 {1'b0}}, Qcnt_three_2[7:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[39:38];
						Q_sqrt1 = {{50 {1'b0}}, Qcnt_three_2[7:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[37:36];
						Q_sqrt2 = {{49 {1'b0}}, Qcnt_three_2[7:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[35:34];
						Q_sqrt0 = {{48 {1'b0}}, Qcnt_three_3[10:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[33:32];
						Q_sqrt1 = {{47 {1'b0}}, Qcnt_three_3[10:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[31:30];
						Q_sqrt2 = {{46 {1'b0}}, Qcnt_three_3[10:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_three_4[13:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_three_4[13:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_three_4[13:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[23:22];
						Q_sqrt0 = {{42 {1'b0}}, Qcnt_three_5[16:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[21:20];
						Q_sqrt1 = {{41 {1'b0}}, Qcnt_three_5[16:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[19:18];
						Q_sqrt2 = {{40 {1'b0}}, Qcnt_three_5[16:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[17:16];
						Q_sqrt0 = {{39 {1'b0}}, Qcnt_three_6[19:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[15:14];
						Q_sqrt1 = {{38 {1'b0}}, Qcnt_three_6[19:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[13:12];
						Q_sqrt2 = {{37 {1'b0}}, Qcnt_three_6[19:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b000111: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[11:10];
						Q_sqrt0 = {{36 {1'b0}}, Qcnt_three_7[22:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[9:8];
						Q_sqrt1 = {{35 {1'b0}}, Qcnt_three_7[22:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[7:6];
						Q_sqrt2 = {{34 {1'b0}}, Qcnt_three_7[22:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_three_8[25:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_three_8[25:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_three_8[25:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{30 {1'b0}}, Qcnt_three_9[28:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{29 {1'b0}}, Qcnt_three_9[28:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{28 {1'b0}}, Qcnt_three_9[28:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{27 {1'b0}}, Qcnt_three_10[31:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{26 {1'b0}}, Qcnt_three_10[31:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{25 {1'b0}}, Qcnt_three_10[31:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{24 {1'b0}}, Qcnt_three_11[34:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{23 {1'b0}}, Qcnt_three_11[34:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{22 {1'b0}}, Qcnt_three_11[34:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_three_12[37:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_three_12[37:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_three_12[37:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{18 {1'b0}}, Qcnt_three_13[40:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{17 {1'b0}}, Qcnt_three_13[40:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{16 {1'b0}}, Qcnt_three_13[40:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001110: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{15 {1'b0}}, Qcnt_three_14[43:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{14 {1'b0}}, Qcnt_three_14[43:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{13 {1'b0}}, Qcnt_three_14[43:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b001111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{12 {1'b0}}, Qcnt_three_15[46:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{11 {1'b0}}, Qcnt_three_15[46:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{10 {1'b0}}, Qcnt_three_15[46:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_three_16[49:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_three_16[49:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_three_16[49:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{6 {1'b0}}, Qcnt_three_17[52:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{5 {1'b0}}, Qcnt_three_17[52:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{4 {1'b0}}, Qcnt_three_17[52:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					6'b010010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{3 {1'b0}}, Qcnt_three_18[55:2]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{2 {1'b0}}, Qcnt_three_18[55:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {1'b0, Qcnt_three_18[55:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
					default: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_three_0[2]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_three_0[2:1]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_three_0[2:0]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
					end
				endcase
			2'b11:
				case (Crtl_cnt_S)
					6'b000000: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000001: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[45:44];
						Q_sqrt0 = {{53 {1'b0}}, Qcnt_four_1[6:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[43:42];
						Q_sqrt1 = {{defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}, Qcnt_four_1[6:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[41:40];
						Q_sqrt2 = {{51 {1'b0}}, Qcnt_four_1[6:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[39:38];
						Q_sqrt3 = {{50 {1'b0}}, Qcnt_four_1[6:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000010: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[37:36];
						Q_sqrt0 = {{49 {1'b0}}, Qcnt_four_2[10:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[35:34];
						Q_sqrt1 = {{48 {1'b0}}, Qcnt_four_2[10:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[33:32];
						Q_sqrt2 = {{47 {1'b0}}, Qcnt_four_2[10:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[31:30];
						Q_sqrt3 = {{46 {1'b0}}, Qcnt_four_2[10:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000011: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[29:28];
						Q_sqrt0 = {{45 {1'b0}}, Qcnt_four_3[14:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[27:26];
						Q_sqrt1 = {{44 {1'b0}}, Qcnt_four_3[14:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[25:24];
						Q_sqrt2 = {{43 {1'b0}}, Qcnt_four_3[14:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[23:22];
						Q_sqrt3 = {{42 {1'b0}}, Qcnt_four_3[14:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000100: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[21:20];
						Q_sqrt0 = {{41 {1'b0}}, Qcnt_four_4[18:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[19:18];
						Q_sqrt1 = {{40 {1'b0}}, Qcnt_four_4[18:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[17:16];
						Q_sqrt2 = {{39 {1'b0}}, Qcnt_four_4[18:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[15:14];
						Q_sqrt3 = {{38 {1'b0}}, Qcnt_four_4[18:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000101: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[13:12];
						Q_sqrt0 = {{37 {1'b0}}, Qcnt_four_5[22:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[11:10];
						Q_sqrt1 = {{36 {1'b0}}, Qcnt_four_5[22:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[9:8];
						Q_sqrt2 = {{35 {1'b0}}, Qcnt_four_5[22:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[7:6];
						Q_sqrt3 = {{34 {1'b0}}, Qcnt_four_5[22:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000110: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[5:4];
						Q_sqrt0 = {{33 {1'b0}}, Qcnt_four_6[26:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = Mant_D_sqrt_Norm[3:2];
						Q_sqrt1 = {{32 {1'b0}}, Qcnt_four_6[26:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[1:0];
						Q_sqrt2 = {{31 {1'b0}}, Qcnt_four_6[26:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{30 {1'b0}}, Qcnt_four_6[26:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b000111: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{29 {1'b0}}, Qcnt_four_7[30:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{28 {1'b0}}, Qcnt_four_7[30:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{27 {1'b0}}, Qcnt_four_7[30:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{26 {1'b0}}, Qcnt_four_7[30:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001000: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{25 {1'b0}}, Qcnt_four_8[34:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{24 {1'b0}}, Qcnt_four_8[34:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{23 {1'b0}}, Qcnt_four_8[34:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{22 {1'b0}}, Qcnt_four_8[34:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001001: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{21 {1'b0}}, Qcnt_four_9[38:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{20 {1'b0}}, Qcnt_four_9[38:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{19 {1'b0}}, Qcnt_four_9[38:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{18 {1'b0}}, Qcnt_four_9[38:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001010: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{17 {1'b0}}, Qcnt_four_10[42:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{16 {1'b0}}, Qcnt_four_10[42:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{15 {1'b0}}, Qcnt_four_10[42:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{14 {1'b0}}, Qcnt_four_10[42:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001011: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{13 {1'b0}}, Qcnt_four_11[46:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{12 {1'b0}}, Qcnt_four_11[46:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{11 {1'b0}}, Qcnt_four_11[46:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{10 {1'b0}}, Qcnt_four_11[46:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001100: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{9 {1'b0}}, Qcnt_four_12[50:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{8 {1'b0}}, Qcnt_four_12[50:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{7 {1'b0}}, Qcnt_four_12[50:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{6 {1'b0}}, Qcnt_four_12[50:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					6'b001101: begin
						Sqrt_DI[0] = 2'b00;
						Q_sqrt0 = {{5 {1'b0}}, Qcnt_four_13[54:3]};
						Sqrt_Q0 = (Quotient_DP[0] ? Q_sqrt_com_0 : Q_sqrt0);
						Sqrt_DI[1] = 2'b00;
						Q_sqrt1 = {{4 {1'b0}}, Qcnt_four_13[54:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = 2'b00;
						Q_sqrt2 = {{3 {1'b0}}, Qcnt_four_13[54:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = 2'b00;
						Q_sqrt3 = {{2 {1'b0}}, Qcnt_four_13[54:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
					default: begin
						Sqrt_DI[0] = Mant_D_sqrt_Norm[53:defs_div_sqrt_mvp_C_MANT_FP64];
						Q_sqrt0 = {{57 {1'b0}}, Qcnt_four_0[3]};
						Sqrt_Q0 = Q_sqrt_com_0;
						Sqrt_DI[1] = Mant_D_sqrt_Norm[51:50];
						Q_sqrt1 = {{56 {1'b0}}, Qcnt_four_0[3:2]};
						Sqrt_Q1 = (Sqrt_quotinent_S[3] ? Q_sqrt_com_1 : Q_sqrt1);
						Sqrt_DI[2] = Mant_D_sqrt_Norm[49:48];
						Q_sqrt2 = {{55 {1'b0}}, Qcnt_four_0[3:1]};
						Sqrt_Q2 = (Sqrt_quotinent_S[2] ? Q_sqrt_com_2 : Q_sqrt2);
						Sqrt_DI[3] = Mant_D_sqrt_Norm[47:46];
						Q_sqrt3 = {{54 {1'b0}}, Qcnt_four_0[3:0]};
						Sqrt_Q3 = (Sqrt_quotinent_S[1] ? Q_sqrt_com_3 : Q_sqrt3);
					end
				endcase
		endcase
	assign Sqrt_R0 = (Sqrt_start_dly_S ? {58 {1'sb0}} : {Partial_remainder_DP[57:0]});
	assign Sqrt_R1 = {Iteration_cell_sum_AMASK_D[0][57], Iteration_cell_sum_AMASK_D[0][54:0], Sqrt_DO[0]};
	assign Sqrt_R2 = {Iteration_cell_sum_AMASK_D[1][57], Iteration_cell_sum_AMASK_D[1][54:0], Sqrt_DO[1]};
	assign Sqrt_R3 = {Iteration_cell_sum_AMASK_D[2][57], Iteration_cell_sum_AMASK_D[2][54:0], Sqrt_DO[2]};
	assign Sqrt_R4 = {Iteration_cell_sum_AMASK_D[3][57], Iteration_cell_sum_AMASK_D[3][54:0], Sqrt_DO[3]};
	wire [57:0] Denominator_se_format_DB;
	assign Denominator_se_format_DB = {Denominator_se_DB[53:45], (FP16ALT_SO ? FP16ALT_SO : Denominator_se_DB[44]), Denominator_se_DB[43:42], (FP16_SO ? FP16_SO : Denominator_se_DB[41]), Denominator_se_DB[40:29], (FP32_SO ? FP32_SO : Denominator_se_DB[28]), Denominator_se_DB[27:0], FP64_SO, 3'b000};
	wire [57:0] First_iteration_cell_div_a_D;
	wire [57:0] First_iteration_cell_div_b_D;
	wire Sel_b_for_first_S;
	assign First_iteration_cell_div_a_D = (Div_start_dly_S ? {Numerator_se_D[53:45], (FP16ALT_SO ? FP16ALT_SO : Numerator_se_D[44]), Numerator_se_D[43:42], (FP16_SO ? FP16_SO : Numerator_se_D[41]), Numerator_se_D[40:29], (FP32_SO ? FP32_SO : Numerator_se_D[28]), Numerator_se_D[27:0], FP64_SO, 3'b000} : {Partial_remainder_DP[56:48], (FP16ALT_SO ? Quotient_DP[0] : Partial_remainder_DP[47]), Partial_remainder_DP[46:45], (FP16_SO ? Quotient_DP[0] : Partial_remainder_DP[44]), Partial_remainder_DP[43:32], (FP32_SO ? Quotient_DP[0] : Partial_remainder_DP[31]), Partial_remainder_DP[30:3], FP64_SO && Quotient_DP[0], 3'b000});
	assign Sel_b_for_first_S = (Div_start_dly_S ? 1 : Quotient_DP[0]);
	assign First_iteration_cell_div_b_D = (Sel_b_for_first_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
	assign Iteration_cell_a_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_R0 : {First_iteration_cell_div_a_D});
	assign Iteration_cell_b_BMASK_D[0] = (Sqrt_enable_SO ? Sqrt_Q0 : {First_iteration_cell_div_b_D});
	wire [57:0] Sec_iteration_cell_div_a_D;
	wire [57:0] Sec_iteration_cell_div_b_D;
	wire Sel_b_for_sec_S;
	generate
		if (|defs_div_sqrt_mvp_Iteration_unit_num_S) begin : genblk1
			assign Sel_b_for_sec_S = ~Iteration_cell_sum_AMASK_D[0][57];
			assign Sec_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[0][56:48], (FP16ALT_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][47]), Iteration_cell_sum_AMASK_D[0][46:45], (FP16_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][44]), Iteration_cell_sum_AMASK_D[0][43:32], (FP32_SO ? Sel_b_for_sec_S : Iteration_cell_sum_AMASK_D[0][31]), Iteration_cell_sum_AMASK_D[0][30:3], FP64_SO && Sel_b_for_sec_S, 3'b000};
			assign Sec_iteration_cell_div_b_D = (Sel_b_for_sec_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			assign Iteration_cell_a_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_R1 : {Sec_iteration_cell_div_a_D});
			assign Iteration_cell_b_BMASK_D[1] = (Sqrt_enable_SO ? Sqrt_Q1 : {Sec_iteration_cell_div_b_D});
		end
	endgenerate
	wire [57:0] Thi_iteration_cell_div_a_D;
	wire [57:0] Thi_iteration_cell_div_b_D;
	wire Sel_b_for_thi_S;
	generate
		if (1'd1 | 1'd0) begin : genblk2
			assign Sel_b_for_thi_S = ~Iteration_cell_sum_AMASK_D[1][57];
			assign Thi_iteration_cell_div_a_D = {Iteration_cell_sum_AMASK_D[1][56:48], (FP16ALT_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][47]), Iteration_cell_sum_AMASK_D[1][46:45], (FP16_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][44]), Iteration_cell_sum_AMASK_D[1][43:32], (FP32_SO ? Sel_b_for_thi_S : Iteration_cell_sum_AMASK_D[1][31]), Iteration_cell_sum_AMASK_D[1][30:3], FP64_SO && Sel_b_for_thi_S, 3'b000};
			assign Thi_iteration_cell_div_b_D = (Sel_b_for_thi_S ? Denominator_se_format_DB : {Denominator_se_D, 4'b0000});
			assign Iteration_cell_a_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_R2 : {Thi_iteration_cell_div_a_D});
			assign Iteration_cell_b_BMASK_D[2] = (Sqrt_enable_SO ? Sqrt_Q2 : {Thi_iteration_cell_div_b_D});
		end
	endgenerate
	wire [57:0] Fou_iteration_cell_div_a_D;
	wire [57:0] Fou_iteration_cell_div_b_D;
	wire Sel_b_for_fou_S;
	wire [57:0] Mask_bits_ctl_S;
	assign Mask_bits_ctl_S = 58'h3ffffffffffffff;
	wire Div_enable_SI [3:0];
	wire Div_start_dly_SI [3:0];
	wire Sqrt_enable_SI [3:0];
	genvar i;
	genvar j;
	generate
		for (i = 0; i <= defs_div_sqrt_mvp_Iteration_unit_num_S; i = i + 1) begin : genblk4
			for (j = 0; j <= 57; j = j + 1) begin : genblk1
				assign Iteration_cell_a_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_a_BMASK_D[i][j];
				assign Iteration_cell_b_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_b_BMASK_D[i][j];
				assign Iteration_cell_sum_AMASK_D[i][j] = Mask_bits_ctl_S[j] && Iteration_cell_sum_D[i][j];
			end
			assign Div_enable_SI[i] = Div_enable_SO;
			assign Div_start_dly_SI[i] = Div_start_dly_S;
			assign Sqrt_enable_SI[i] = Sqrt_enable_SO;
			iteration_div_sqrt_mvp #(.WIDTH(58)) iteration_div_sqrt(
				.A_DI(Iteration_cell_a_D[i]),
				.B_DI(Iteration_cell_b_D[i]),
				.Div_enable_SI(Div_enable_SI[i]),
				.Div_start_dly_SI(Div_start_dly_SI[i]),
				.Sqrt_enable_SI(Sqrt_enable_SI[i]),
				.D_DI(Sqrt_DI[i]),
				.D_DO(Sqrt_DO[i]),
				.Sum_DO(Iteration_cell_sum_D[i]),
				.Carry_out_DO(Iteration_cell_carry_D[i])
			);
		end
	endgenerate
	always @(*)
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				if (Fsm_enable_S)
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R1 : Iteration_cell_sum_AMASK_D[0]);
				else
					Partial_remainder_DN = Partial_remainder_DP;
			2'b01:
				if (Fsm_enable_S)
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R2 : Iteration_cell_sum_AMASK_D[1]);
				else
					Partial_remainder_DN = Partial_remainder_DP;
			2'b10:
				if (Fsm_enable_S)
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R3 : Iteration_cell_sum_AMASK_D[2]);
				else
					Partial_remainder_DN = Partial_remainder_DP;
			2'b11:
				if (Fsm_enable_S)
					Partial_remainder_DN = (Sqrt_enable_SO ? Sqrt_R4 : Iteration_cell_sum_AMASK_D[3]);
				else
					Partial_remainder_DN = Partial_remainder_DP;
		endcase
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Partial_remainder_DP <= 1'sb0;
		else
			Partial_remainder_DP <= Partial_remainder_DN;
	reg [56:0] Quotient_DN;
	always @(*)
		case (defs_div_sqrt_mvp_Iteration_unit_num_S)
			2'b00:
				if (Fsm_enable_S)
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[55:0], Sqrt_quotinent_S[3]} : {Quotient_DP[55:0], Iteration_cell_carry_D[0]});
				else
					Quotient_DN = Quotient_DP;
			2'b01:
				if (Fsm_enable_S)
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[54:0], Sqrt_quotinent_S[3:2]} : {Quotient_DP[54:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1]});
				else
					Quotient_DN = Quotient_DP;
			2'b10:
				if (Fsm_enable_S)
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[53:0], Sqrt_quotinent_S[3:1]} : {Quotient_DP[53:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2]});
				else
					Quotient_DN = Quotient_DP;
			2'b11:
				if (Fsm_enable_S)
					Quotient_DN = (Sqrt_enable_SO ? {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Sqrt_quotinent_S} : {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP64:0], Iteration_cell_carry_D[0], Iteration_cell_carry_D[1], Iteration_cell_carry_D[2], Iteration_cell_carry_D[3]});
				else
					Quotient_DN = Quotient_DP;
		endcase
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Quotient_DP <= 1'sb0;
		else
			Quotient_DP <= Quotient_DN;
	generate
		if (1) begin : genblk7
			always @(*)
				case (Format_sel_S)
					2'b00:
						case (Precision_ctl_S)
							6'h00: Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15: Mant_result_prenorm_DO = {Quotient_DP[defs_div_sqrt_mvp_C_MANT_FP32:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12: Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f: Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c: Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09: Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06: Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default: Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
						endcase
					2'b01:
						case (Precision_ctl_S)
							6'h00: Mant_result_prenorm_DO = Quotient_DP[56:0];
							6'h34, 6'h33: Mant_result_prenorm_DO = {Quotient_DP[53:1], {4 {1'b0}}};
							6'h32, 6'h31, 6'h30: Mant_result_prenorm_DO = {Quotient_DP[50:0], {6 {1'b0}}};
							6'h2f, 6'h2e, 6'h2d: Mant_result_prenorm_DO = {Quotient_DP[47:0], {9 {1'b0}}};
							6'h2c, 6'h2b, 6'h2a: Mant_result_prenorm_DO = {Quotient_DP[44:0], {12 {1'b0}}};
							6'h29, 6'h28, 6'h27: Mant_result_prenorm_DO = {Quotient_DP[41:0], {15 {1'b0}}};
							6'h26, 6'h25, 6'h24: Mant_result_prenorm_DO = {Quotient_DP[38:0], {18 {1'b0}}};
							6'h23, 6'h22, 6'h21: Mant_result_prenorm_DO = {Quotient_DP[35:0], {21 {1'b0}}};
							6'h20, 6'h1f, 6'h1e: Mant_result_prenorm_DO = {Quotient_DP[32:0], {24 {1'b0}}};
							6'h1d, 6'h1c, 6'h1b: Mant_result_prenorm_DO = {Quotient_DP[29:0], {27 {1'b0}}};
							6'h1a, 6'h19, 6'h18: Mant_result_prenorm_DO = {Quotient_DP[26:0], {30 {1'b0}}};
							6'h17, 6'h16, 6'h15: Mant_result_prenorm_DO = {Quotient_DP[23:0], {33 {1'b0}}};
							6'h14, 6'h13, 6'h12: Mant_result_prenorm_DO = {Quotient_DP[20:0], {36 {1'b0}}};
							6'h11, 6'h10, 6'h0f: Mant_result_prenorm_DO = {Quotient_DP[17:0], {39 {1'b0}}};
							6'h0e, 6'h0d, 6'h0c: Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0b, 6'h0a, 6'h09: Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h08, 6'h07, 6'h06: Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default: Mant_result_prenorm_DO = Quotient_DP[56:0];
						endcase
					2'b10:
						case (Precision_ctl_S)
							6'b000000: Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
							6'h0a, 6'h09: Mant_result_prenorm_DO = {Quotient_DP[11:1], {46 {1'b0}}};
							6'h08, 6'h07, 6'h06: Mant_result_prenorm_DO = {Quotient_DP[8:0], {48 {1'b0}}};
							default: Mant_result_prenorm_DO = {Quotient_DP[14:0], {42 {1'b0}}};
						endcase
					2'b11:
						case (Precision_ctl_S)
							6'b000000: Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
							6'h07, 6'h06: Mant_result_prenorm_DO = {Quotient_DP[8:1], {49 {1'b0}}};
							default: Mant_result_prenorm_DO = {Quotient_DP[11:0], {45 {1'b0}}};
						endcase
				endcase
		end
	endgenerate
	wire [12:0] Exp_result_prenorm_DN;
	reg [12:0] Exp_result_prenorm_DP;
	wire [12:0] Exp_add_a_D;
	wire [12:0] Exp_add_b_D;
	wire [12:0] Exp_add_c_D;
	integer C_BIAS_AONE;
	integer C_HALF_BIAS;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16 = 5'h10;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP32 = 8'h80;
	localparam defs_div_sqrt_mvp_C_BIAS_AONE_FP64 = 11'h400;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16 = 7;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP32 = 63;
	localparam defs_div_sqrt_mvp_C_HALF_BIAS_FP64 = 511;
	always @(*)
		case (Format_sel_S)
			2'b00: begin
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP32;
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP32;
			end
			2'b01: begin
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP64;
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP64;
			end
			2'b10: begin
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16;
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16;
			end
			2'b11: begin
				C_BIAS_AONE = defs_div_sqrt_mvp_C_BIAS_AONE_FP16ALT;
				C_HALF_BIAS = defs_div_sqrt_mvp_C_HALF_BIAS_FP16ALT;
			end
		endcase
	assign Exp_add_a_D = {(Sqrt_start_dly_S ? {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64:1]} : {Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI[defs_div_sqrt_mvp_C_EXP_FP64], Exp_num_DI})};
	localparam defs_div_sqrt_mvp_C_EXP_ZERO_FP64 = 11'h000;
	assign Exp_add_b_D = {(Sqrt_start_dly_S ? {1'b0, defs_div_sqrt_mvp_C_EXP_ZERO_FP64, Exp_num_DI[0]} : {~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI[defs_div_sqrt_mvp_C_EXP_FP64], ~Exp_den_DI})};
	assign Exp_add_c_D = {(Div_start_dly_S ? {C_BIAS_AONE} : {C_HALF_BIAS})};
	assign Exp_result_prenorm_DN = (Start_dly_S ? {(Exp_add_a_D + Exp_add_b_D) + Exp_add_c_D} : Exp_result_prenorm_DP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Exp_result_prenorm_DP <= 1'sb0;
		else
			Exp_result_prenorm_DP <= Exp_result_prenorm_DN;
	assign Exp_result_prenorm_DO = Exp_result_prenorm_DP;
endmodule
module div_sqrt_top_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Precision_ctl_SI,
	Format_sel_SI,
	Kill_SI,
	Result_DO,
	Fflags_SO,
	Ready_SO,
	Done_SO
);
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire Div_start_SI;
	input wire Sqrt_start_SI;
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	input wire [63:0] Operand_b_DI;
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	input wire Kill_SI;
	output wire [63:0] Result_DO;
	output wire [4:0] Fflags_SO;
	output wire Ready_SO;
	output wire Done_SO;
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_D;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_D;
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	wire [12:0] Exp_z_D;
	wire [56:0] Mant_z_D;
	wire Sign_z_D;
	wire Start_S;
	wire [2:0] RM_dly_S;
	wire Div_enable_S;
	wire Sqrt_enable_S;
	wire Inf_a_S;
	wire Inf_b_S;
	wire Zero_a_S;
	wire Zero_b_S;
	wire NaN_a_S;
	wire NaN_b_S;
	wire SNaN_S;
	wire Special_case_SB;
	wire Special_case_dly_SB;
	wire Full_precision_S;
	wire FP32_S;
	wire FP64_S;
	wire FP16_S;
	wire FP16ALT_S;
	preprocess_mvp preprocess_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Ready_SI(Ready_SO),
		.Operand_a_DI(Operand_a_DI),
		.Operand_b_DI(Operand_b_DI),
		.RM_SI(RM_SI),
		.Format_sel_SI(Format_sel_SI),
		.Start_SO(Start_S),
		.Exp_a_DO_norm(Exp_a_D),
		.Exp_b_DO_norm(Exp_b_D),
		.Mant_a_DO_norm(Mant_a_D),
		.Mant_b_DO_norm(Mant_b_D),
		.RM_dly_SO(RM_dly_S),
		.Sign_z_DO(Sign_z_D),
		.Inf_a_SO(Inf_a_S),
		.Inf_b_SO(Inf_b_S),
		.Zero_a_SO(Zero_a_S),
		.Zero_b_SO(Zero_b_S),
		.NaN_a_SO(NaN_a_S),
		.NaN_b_SO(NaN_b_S),
		.SNaN_SO(SNaN_S),
		.Special_case_SBO(Special_case_SB),
		.Special_case_dly_SBO(Special_case_dly_SB)
	);
	nrbd_nrsc_mvp nrbd_nrsc_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_S),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SB),
		.Special_case_dly_SBI(Special_case_dly_SB),
		.Div_enable_SO(Div_enable_S),
		.Sqrt_enable_SO(Sqrt_enable_S),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Exp_a_DI(Exp_a_D),
		.Exp_b_DI(Exp_b_D),
		.Mant_a_DI(Mant_a_D),
		.Mant_b_DI(Mant_b_D),
		.Full_precision_SO(Full_precision_S),
		.FP32_SO(FP32_S),
		.FP64_SO(FP64_S),
		.FP16_SO(FP16_S),
		.FP16ALT_SO(FP16ALT_S),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Exp_z_DO(Exp_z_D),
		.Mant_z_DO(Mant_z_D)
	);
	norm_div_sqrt_mvp fpu_norm_U0(
		.Mant_in_DI(Mant_z_D),
		.Exp_in_DI(Exp_z_D),
		.Sign_in_DI(Sign_z_D),
		.Div_enable_SI(Div_enable_S),
		.Sqrt_enable_SI(Sqrt_enable_S),
		.Inf_a_SI(Inf_a_S),
		.Inf_b_SI(Inf_b_S),
		.Zero_a_SI(Zero_a_S),
		.Zero_b_SI(Zero_b_S),
		.NaN_a_SI(NaN_a_S),
		.NaN_b_SI(NaN_b_S),
		.SNaN_SI(SNaN_S),
		.RM_SI(RM_dly_S),
		.Full_precision_SI(Full_precision_S),
		.FP32_SI(FP32_S),
		.FP64_SI(FP64_S),
		.FP16_SI(FP16_S),
		.FP16ALT_SI(FP16ALT_S),
		.Result_DO(Result_DO),
		.Fflags_SO(Fflags_SO)
	);
endmodule
module iteration_div_sqrt_mvp (
	A_DI,
	B_DI,
	Div_enable_SI,
	Div_start_dly_SI,
	Sqrt_enable_SI,
	D_DI,
	D_DO,
	Sum_DO,
	Carry_out_DO
);
	parameter WIDTH = 25;
	input wire [WIDTH - 1:0] A_DI;
	input wire [WIDTH - 1:0] B_DI;
	input wire Div_enable_SI;
	input wire Div_start_dly_SI;
	input wire Sqrt_enable_SI;
	input wire [1:0] D_DI;
	output wire [1:0] D_DO;
	output wire [WIDTH - 1:0] Sum_DO;
	output wire Carry_out_DO;
	wire D_carry_D;
	wire Sqrt_cin_D;
	wire Cin_D;
	assign D_DO[0] = ~D_DI[0];
	assign D_DO[1] = ~(D_DI[1] ^ D_DI[0]);
	assign D_carry_D = D_DI[1] | D_DI[0];
	assign Sqrt_cin_D = Sqrt_enable_SI && D_carry_D;
	assign Cin_D = (Div_enable_SI ? 1'b0 : Sqrt_cin_D);
	assign {Carry_out_DO, Sum_DO} = (A_DI + B_DI) + Cin_D;
endmodule
module norm_div_sqrt_mvp (
	Mant_in_DI,
	Exp_in_DI,
	Sign_in_DI,
	Div_enable_SI,
	Sqrt_enable_SI,
	Inf_a_SI,
	Inf_b_SI,
	Zero_a_SI,
	Zero_b_SI,
	NaN_a_SI,
	NaN_b_SI,
	SNaN_SI,
	RM_SI,
	Full_precision_SI,
	FP32_SI,
	FP64_SI,
	FP16_SI,
	FP16ALT_SI,
	Result_DO,
	Fflags_SO
);
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [56:0] Mant_in_DI;
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire signed [12:0] Exp_in_DI;
	input wire Sign_in_DI;
	input wire Div_enable_SI;
	input wire Sqrt_enable_SI;
	input wire Inf_a_SI;
	input wire Inf_b_SI;
	input wire Zero_a_SI;
	input wire Zero_b_SI;
	input wire NaN_a_SI;
	input wire NaN_b_SI;
	input wire SNaN_SI;
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	input wire Full_precision_SI;
	input wire FP32_SI;
	input wire FP64_SI;
	input wire FP16_SI;
	input wire FP16ALT_SI;
	output reg [63:0] Result_DO;
	output wire [4:0] Fflags_SO;
	reg Sign_res_D;
	reg NV_OP_S;
	reg Exp_OF_S;
	reg Exp_UF_S;
	reg Div_Zero_S;
	wire In_Exact_S;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_res_norm_D;
	reg [10:0] Exp_res_norm_D;
	wire [12:0] Exp_Max_RS_FP64_D;
	localparam defs_div_sqrt_mvp_C_EXP_FP32 = 8;
	wire [9:0] Exp_Max_RS_FP32_D;
	localparam defs_div_sqrt_mvp_C_EXP_FP16 = 5;
	wire [6:0] Exp_Max_RS_FP16_D;
	localparam defs_div_sqrt_mvp_C_EXP_FP16ALT = 8;
	wire [9:0] Exp_Max_RS_FP16ALT_D;
	assign Exp_Max_RS_FP64_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] + defs_div_sqrt_mvp_C_MANT_FP64) + 1;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	assign Exp_Max_RS_FP32_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32:0] + defs_div_sqrt_mvp_C_MANT_FP32) + 1;
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	assign Exp_Max_RS_FP16_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16:0] + defs_div_sqrt_mvp_C_MANT_FP16) + 1;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	assign Exp_Max_RS_FP16ALT_D = (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT:0] + defs_div_sqrt_mvp_C_MANT_FP16ALT) + 1;
	wire [12:0] Num_RS_D;
	assign Num_RS_D = ~Exp_in_DI + 2;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_RS_D;
	wire [56:0] Mant_forsticky_D;
	assign {Mant_RS_D, Mant_forsticky_D} = {Mant_in_DI, {53 {1'b0}}} >> Num_RS_D;
	wire [12:0] Exp_subOne_D;
	assign Exp_subOne_D = Exp_in_DI - 1;
	reg [1:0] Mant_lower_D;
	reg Mant_sticky_bit_D;
	reg [56:0] Mant_forround_D;
	localparam defs_div_sqrt_mvp_C_EXP_ONE_FP64 = 13'h0001;
	localparam defs_div_sqrt_mvp_C_MANT_NAN_FP64 = 52'h8000000000000;
	always @(*)
		if (NaN_a_SI) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			Exp_res_norm_D = 1'sb1;
			Mant_forround_D = 1'sb0;
			Sign_res_D = 1'b0;
			NV_OP_S = SNaN_SI;
		end
		else if (NaN_b_SI) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			Exp_res_norm_D = 1'sb1;
			Mant_forround_D = 1'sb0;
			Sign_res_D = 1'b0;
			NV_OP_S = SNaN_SI;
		end
		else if (Inf_a_SI) begin
			if (Div_enable_SI && Inf_b_SI) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = 1'b0;
				NV_OP_S = 1'b1;
			end
			else if (Sqrt_enable_SI && Sign_in_DI) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = 1'b0;
				NV_OP_S = 1'b1;
			end
			else begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b1;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
		end
		else if (Div_enable_SI && Inf_b_SI) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b1;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = 1'sb0;
			Exp_res_norm_D = 1'sb0;
			Mant_forround_D = 1'sb0;
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
		else if (Zero_a_SI) begin
			if (Div_enable_SI && Zero_b_SI) begin
				Div_Zero_S = 1'b1;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = 1'b0;
				NV_OP_S = 1'b1;
			end
			else begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb0;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
		end
		else if (Div_enable_SI && Zero_b_SI) begin
			Div_Zero_S = 1'b1;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = 1'sb0;
			Exp_res_norm_D = 1'sb1;
			Mant_forround_D = 1'sb0;
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
		else if (Sign_in_DI && Sqrt_enable_SI) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = {1'b0, defs_div_sqrt_mvp_C_MANT_NAN_FP64};
			Exp_res_norm_D = 1'sb1;
			Mant_forround_D = 1'sb0;
			Sign_res_D = 1'b0;
			NV_OP_S = 1'b1;
		end
		else if (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == {12 {1'sb0}}) begin
			if (Mant_in_DI != {57 {1'sb0}}) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b1;
				Mant_res_norm_D = {1'b0, Mant_in_DI[56:5]};
				Exp_res_norm_D = 1'sb0;
				Mant_forround_D = {Mant_in_DI[4:0], {defs_div_sqrt_mvp_C_MANT_FP64 {1'b0}}};
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
			else begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb0;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
		end
		else if ((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64:0] == defs_div_sqrt_mvp_C_EXP_ONE_FP64) && ~Mant_in_DI[56]) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b1;
			Mant_res_norm_D = Mant_in_DI[56:4];
			Exp_res_norm_D = 1'sb0;
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
		else if (Exp_in_DI[12]) begin
			if ((((~Exp_Max_RS_FP32_D[9] && FP32_SI) | (~Exp_Max_RS_FP64_D[12] && FP64_SI)) | (~Exp_Max_RS_FP16_D[6] && FP16_SI)) | (~Exp_Max_RS_FP16ALT_D[9] && FP16ALT_SI)) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b1;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb0;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
			else begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b1;
				Mant_res_norm_D = {Mant_RS_D[defs_div_sqrt_mvp_C_MANT_FP64:0]};
				Exp_res_norm_D = 1'sb0;
				Mant_forround_D = {Mant_forsticky_D[56:0]};
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
		end
		else if ((((Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP32] && FP32_SI) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP64] && FP64_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16] && FP16_SI)) | (Exp_in_DI[defs_div_sqrt_mvp_C_EXP_FP16ALT] && FP16ALT_SI)) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b1;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = 1'sb0;
			Exp_res_norm_D = 1'sb1;
			Mant_forround_D = 1'sb0;
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
		else if (((((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP32_SI) | ((Exp_in_DI[10:0] == {11 {1'sb1}}) && FP64_SI)) | ((Exp_in_DI[4:0] == {5 {1'sb1}}) && FP16_SI)) | ((Exp_in_DI[7:0] == {8 {1'sb1}}) && FP16ALT_SI)) begin
			if (~Mant_in_DI[56]) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b0;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = Mant_in_DI[55:3];
				Exp_res_norm_D = Exp_subOne_D;
				Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
			else if (Mant_in_DI != {57 {1'sb0}}) begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b1;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
			else begin
				Div_Zero_S = 1'b0;
				Exp_OF_S = 1'b1;
				Exp_UF_S = 1'b0;
				Mant_res_norm_D = 1'sb0;
				Exp_res_norm_D = 1'sb1;
				Mant_forround_D = 1'sb0;
				Sign_res_D = Sign_in_DI;
				NV_OP_S = 1'b0;
			end
		end
		else if (Mant_in_DI[56]) begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = Mant_in_DI[56:4];
			Exp_res_norm_D = Exp_in_DI[10:0];
			Mant_forround_D = {Mant_in_DI[3:0], {53 {1'b0}}};
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
		else begin
			Div_Zero_S = 1'b0;
			Exp_OF_S = 1'b0;
			Exp_UF_S = 1'b0;
			Mant_res_norm_D = Mant_in_DI[55:3];
			Exp_res_norm_D = Exp_subOne_D;
			Mant_forround_D = {Mant_in_DI[2:0], {54 {1'b0}}};
			Sign_res_D = Sign_in_DI;
			NV_OP_S = 1'b0;
		end
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_upper_D;
	wire [53:0] Mant_upperRounded_D;
	reg Mant_roundUp_S;
	wire Mant_rounded_S;
	always @(*)
		if (FP32_SI) begin
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:29], {29 {1'b0}}};
			Mant_lower_D = Mant_res_norm_D[28:27];
			Mant_sticky_bit_D = |Mant_res_norm_D[26:0];
		end
		else if (FP64_SI) begin
			Mant_upper_D = Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:0];
			Mant_lower_D = Mant_forround_D[56:55];
			Mant_sticky_bit_D = |Mant_forround_D[55:0];
		end
		else if (FP16_SI) begin
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:42], {42 {1'b0}}};
			Mant_lower_D = Mant_res_norm_D[41:40];
			Mant_sticky_bit_D = |Mant_res_norm_D[39:30];
		end
		else begin
			Mant_upper_D = {Mant_res_norm_D[defs_div_sqrt_mvp_C_MANT_FP64:45], {45 {1'b0}}};
			Mant_lower_D = Mant_res_norm_D[44:43];
			Mant_sticky_bit_D = |Mant_res_norm_D[42:30];
		end
	assign Mant_rounded_S = |Mant_lower_D | Mant_sticky_bit_D;
	localparam defs_div_sqrt_mvp_C_RM_MINUSINF = 3'h3;
	localparam defs_div_sqrt_mvp_C_RM_NEAREST = 3'h0;
	localparam defs_div_sqrt_mvp_C_RM_PLUSINF = 3'h2;
	localparam defs_div_sqrt_mvp_C_RM_TRUNC = 3'h1;
	always @(*) begin
		Mant_roundUp_S = 1'b0;
		case (RM_SI)
			defs_div_sqrt_mvp_C_RM_NEAREST: Mant_roundUp_S = Mant_lower_D[1] && ((Mant_lower_D[0] | Mant_sticky_bit_D) | ((((FP32_SI && Mant_upper_D[29]) | (FP64_SI && Mant_upper_D[0])) | (FP16_SI && Mant_upper_D[42])) | (FP16ALT_SI && Mant_upper_D[45])));
			defs_div_sqrt_mvp_C_RM_TRUNC: Mant_roundUp_S = 0;
			defs_div_sqrt_mvp_C_RM_PLUSINF: Mant_roundUp_S = Mant_rounded_S & ~Sign_in_DI;
			defs_div_sqrt_mvp_C_RM_MINUSINF: Mant_roundUp_S = Mant_rounded_S & Sign_in_DI;
			default: Mant_roundUp_S = 0;
		endcase
	end
	wire Mant_renorm_S;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_roundUp_Vector_S;
	assign Mant_roundUp_Vector_S = {7'h00, FP16ALT_SI && Mant_roundUp_S, 2'h0, FP16_SI && Mant_roundUp_S, 12'h000, FP32_SI && Mant_roundUp_S, 28'h0000000, FP64_SI && Mant_roundUp_S};
	assign Mant_upperRounded_D = Mant_upper_D + Mant_roundUp_Vector_S;
	assign Mant_renorm_S = Mant_upperRounded_D[53];
	wire [51:0] Mant_res_round_D;
	wire [10:0] Exp_res_round_D;
	assign Mant_res_round_D = (Mant_renorm_S ? Mant_upperRounded_D[defs_div_sqrt_mvp_C_MANT_FP64:1] : Mant_upperRounded_D[51:0]);
	assign Exp_res_round_D = Exp_res_norm_D + Mant_renorm_S;
	wire [51:0] Mant_before_format_ctl_D;
	wire [10:0] Exp_before_format_ctl_D;
	assign Mant_before_format_ctl_D = (Full_precision_SI ? Mant_res_round_D : Mant_res_norm_D);
	assign Exp_before_format_ctl_D = (Full_precision_SI ? Exp_res_round_D : Exp_res_norm_D);
	always @(*)
		if (FP32_SI)
			Result_DO = {32'hffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:29]};
		else if (FP64_SI)
			Result_DO = {Sign_res_D, Exp_before_format_ctl_D[10:0], Mant_before_format_ctl_D[51:0]};
		else if (FP16_SI)
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[4:0], Mant_before_format_ctl_D[51:42]};
		else
			Result_DO = {48'hffffffffffff, Sign_res_D, Exp_before_format_ctl_D[7:0], Mant_before_format_ctl_D[51:45]};
	assign In_Exact_S = ~Full_precision_SI | Mant_rounded_S;
	assign Fflags_SO = {NV_OP_S, Div_Zero_S, Exp_OF_S, Exp_UF_S, In_Exact_S};
endmodule
module nrbd_nrsc_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Start_SI,
	Kill_SI,
	Special_case_SBI,
	Special_case_dly_SBI,
	Precision_ctl_SI,
	Format_sel_SI,
	Mant_a_DI,
	Mant_b_DI,
	Exp_a_DI,
	Exp_b_DI,
	Div_enable_SO,
	Sqrt_enable_SO,
	Full_precision_SO,
	FP32_SO,
	FP64_SO,
	FP16_SO,
	FP16ALT_SO,
	Ready_SO,
	Done_SO,
	Mant_z_DO,
	Exp_z_DO
);
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire Div_start_SI;
	input wire Sqrt_start_SI;
	input wire Start_SI;
	input wire Kill_SI;
	input wire Special_case_SBI;
	input wire Special_case_dly_SBI;
	localparam defs_div_sqrt_mvp_C_PC = 6;
	input wire [5:0] Precision_ctl_SI;
	input wire [1:0] Format_sel_SI;
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DI;
	input wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DI;
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DI;
	input wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DI;
	output wire Div_enable_SO;
	output wire Sqrt_enable_SO;
	output wire Full_precision_SO;
	output wire FP32_SO;
	output wire FP64_SO;
	output wire FP16_SO;
	output wire FP16ALT_SO;
	output wire Ready_SO;
	output wire Done_SO;
	output wire [56:0] Mant_z_DO;
	output wire [12:0] Exp_z_DO;
	wire Div_start_dly_S;
	wire Sqrt_start_dly_S;
	control_mvp control_U0(
		.Clk_CI(Clk_CI),
		.Rst_RBI(Rst_RBI),
		.Div_start_SI(Div_start_SI),
		.Sqrt_start_SI(Sqrt_start_SI),
		.Start_SI(Start_SI),
		.Kill_SI(Kill_SI),
		.Special_case_SBI(Special_case_SBI),
		.Special_case_dly_SBI(Special_case_dly_SBI),
		.Precision_ctl_SI(Precision_ctl_SI),
		.Format_sel_SI(Format_sel_SI),
		.Numerator_DI(Mant_a_DI),
		.Exp_num_DI(Exp_a_DI),
		.Denominator_DI(Mant_b_DI),
		.Exp_den_DI(Exp_b_DI),
		.Div_start_dly_SO(Div_start_dly_S),
		.Sqrt_start_dly_SO(Sqrt_start_dly_S),
		.Div_enable_SO(Div_enable_SO),
		.Sqrt_enable_SO(Sqrt_enable_SO),
		.Full_precision_SO(Full_precision_SO),
		.FP32_SO(FP32_SO),
		.FP64_SO(FP64_SO),
		.FP16_SO(FP16_SO),
		.FP16ALT_SO(FP16ALT_SO),
		.Ready_SO(Ready_SO),
		.Done_SO(Done_SO),
		.Mant_result_prenorm_DO(Mant_z_DO),
		.Exp_result_prenorm_DO(Exp_z_DO)
	);
endmodule
module preprocess_mvp (
	Clk_CI,
	Rst_RBI,
	Div_start_SI,
	Sqrt_start_SI,
	Ready_SI,
	Operand_a_DI,
	Operand_b_DI,
	RM_SI,
	Format_sel_SI,
	Start_SO,
	Exp_a_DO_norm,
	Exp_b_DO_norm,
	Mant_a_DO_norm,
	Mant_b_DO_norm,
	RM_dly_SO,
	Sign_z_DO,
	Inf_a_SO,
	Inf_b_SO,
	Zero_a_SO,
	Zero_b_SO,
	NaN_a_SO,
	NaN_b_SO,
	SNaN_SO,
	Special_case_SBO,
	Special_case_dly_SBO
);
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire Div_start_SI;
	input wire Sqrt_start_SI;
	input wire Ready_SI;
	localparam defs_div_sqrt_mvp_C_OP_FP64 = 64;
	input wire [63:0] Operand_a_DI;
	input wire [63:0] Operand_b_DI;
	localparam defs_div_sqrt_mvp_C_RM = 3;
	input wire [2:0] RM_SI;
	localparam defs_div_sqrt_mvp_C_FS = 2;
	input wire [1:0] Format_sel_SI;
	output wire Start_SO;
	localparam defs_div_sqrt_mvp_C_EXP_FP64 = 11;
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_DO_norm;
	output wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_DO_norm;
	localparam defs_div_sqrt_mvp_C_MANT_FP64 = 52;
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_DO_norm;
	output wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_DO_norm;
	output wire [2:0] RM_dly_SO;
	output wire Sign_z_DO;
	output wire Inf_a_SO;
	output wire Inf_b_SO;
	output wire Zero_a_SO;
	output wire Zero_b_SO;
	output wire NaN_a_SO;
	output wire NaN_b_SO;
	output wire SNaN_SO;
	output wire Special_case_SBO;
	output reg Special_case_dly_SBO;
	wire Hb_a_D;
	wire Hb_b_D;
	reg [10:0] Exp_a_D;
	reg [10:0] Exp_b_D;
	reg [51:0] Mant_a_NonH_D;
	reg [51:0] Mant_b_NonH_D;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_D;
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_D;
	reg Sign_a_D;
	reg Sign_b_D;
	wire Start_S;
	localparam defs_div_sqrt_mvp_C_MANT_FP16 = 10;
	localparam defs_div_sqrt_mvp_C_MANT_FP16ALT = 7;
	localparam defs_div_sqrt_mvp_C_MANT_FP32 = 23;
	localparam defs_div_sqrt_mvp_C_OP_FP16 = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP16ALT = 16;
	localparam defs_div_sqrt_mvp_C_OP_FP32 = 32;
	always @(*)
		case (Format_sel_SI)
			2'b00: begin
				Sign_a_D = Operand_a_DI[31];
				Sign_b_D = Operand_b_DI[31];
				Exp_a_D = {3'h0, Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				Exp_b_D = {3'h0, Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32]};
				Mant_a_NonH_D = {Operand_a_DI[22:0], 29'h00000000};
				Mant_b_NonH_D = {Operand_b_DI[22:0], 29'h00000000};
			end
			2'b01: begin
				Sign_a_D = Operand_a_DI[63];
				Sign_b_D = Operand_b_DI[63];
				Exp_a_D = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				Exp_b_D = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64];
				Mant_a_NonH_D = Operand_a_DI[51:0];
				Mant_b_NonH_D = Operand_b_DI[51:0];
			end
			2'b10: begin
				Sign_a_D = Operand_a_DI[15];
				Sign_b_D = Operand_b_DI[15];
				Exp_a_D = {6'h00, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				Exp_b_D = {6'h00, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16]};
				Mant_a_NonH_D = {Operand_a_DI[9:0], 42'h00000000000};
				Mant_b_NonH_D = {Operand_b_DI[9:0], 42'h00000000000};
			end
			2'b11: begin
				Sign_a_D = Operand_a_DI[15];
				Sign_b_D = Operand_b_DI[15];
				Exp_a_D = {3'h0, Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				Exp_b_D = {3'h0, Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT]};
				Mant_a_NonH_D = {Operand_a_DI[6:0], 45'h000000000000};
				Mant_b_NonH_D = {Operand_b_DI[6:0], 45'h000000000000};
			end
		endcase
	assign Mant_a_D = {Hb_a_D, Mant_a_NonH_D};
	assign Mant_b_D = {Hb_b_D, Mant_b_NonH_D};
	assign Hb_a_D = |Exp_a_D;
	assign Hb_b_D = |Exp_b_D;
	assign Start_S = Div_start_SI | Sqrt_start_SI;
	reg Mant_a_prenorm_zero_S;
	reg Mant_b_prenorm_zero_S;
	wire Exp_a_prenorm_zero_S;
	wire Exp_b_prenorm_zero_S;
	assign Exp_a_prenorm_zero_S = ~Hb_a_D;
	assign Exp_b_prenorm_zero_S = ~Hb_b_D;
	reg Exp_a_prenorm_Inf_NaN_S;
	reg Exp_b_prenorm_Inf_NaN_S;
	wire Mant_a_prenorm_QNaN_S;
	wire Mant_a_prenorm_SNaN_S;
	wire Mant_b_prenorm_QNaN_S;
	wire Mant_b_prenorm_SNaN_S;
	assign Mant_a_prenorm_QNaN_S = Mant_a_NonH_D[51] && ~(|Mant_a_NonH_D[50:0]);
	assign Mant_a_prenorm_SNaN_S = ~Mant_a_NonH_D[51] && |Mant_a_NonH_D[50:0];
	assign Mant_b_prenorm_QNaN_S = Mant_b_NonH_D[51] && ~(|Mant_b_NonH_D[50:0]);
	assign Mant_b_prenorm_SNaN_S = ~Mant_b_NonH_D[51] && |Mant_b_NonH_D[50:0];
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16 = 5'h1f;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP16ALT = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP32 = 8'hff;
	localparam defs_div_sqrt_mvp_C_EXP_INF_FP64 = 11'h7ff;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16 = 10'h000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT = 7'h00;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP32 = 23'h000000;
	localparam defs_div_sqrt_mvp_C_MANT_ZERO_FP64 = 52'h0000000000000;
	always @(*)
		case (Format_sel_SI)
			2'b00: begin
				Mant_a_prenorm_zero_S = Operand_a_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				Mant_b_prenorm_zero_S = Operand_b_DI[22:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP32;
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[30:defs_div_sqrt_mvp_C_MANT_FP32] == defs_div_sqrt_mvp_C_EXP_INF_FP32;
			end
			2'b01: begin
				Mant_a_prenorm_zero_S = Operand_a_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				Mant_b_prenorm_zero_S = Operand_b_DI[51:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP64;
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[62:defs_div_sqrt_mvp_C_MANT_FP64] == defs_div_sqrt_mvp_C_EXP_INF_FP64;
			end
			2'b10: begin
				Mant_a_prenorm_zero_S = Operand_a_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				Mant_b_prenorm_zero_S = Operand_b_DI[9:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16;
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16] == defs_div_sqrt_mvp_C_EXP_INF_FP16;
			end
			2'b11: begin
				Mant_a_prenorm_zero_S = Operand_a_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				Mant_b_prenorm_zero_S = Operand_b_DI[6:0] == defs_div_sqrt_mvp_C_MANT_ZERO_FP16ALT;
				Exp_a_prenorm_Inf_NaN_S = Operand_a_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
				Exp_b_prenorm_Inf_NaN_S = Operand_b_DI[14:defs_div_sqrt_mvp_C_MANT_FP16ALT] == defs_div_sqrt_mvp_C_EXP_INF_FP16ALT;
			end
		endcase
	wire Zero_a_SN;
	reg Zero_a_SP;
	wire Zero_b_SN;
	reg Zero_b_SP;
	wire Inf_a_SN;
	reg Inf_a_SP;
	wire Inf_b_SN;
	reg Inf_b_SP;
	wire NaN_a_SN;
	reg NaN_a_SP;
	wire NaN_b_SN;
	reg NaN_b_SP;
	wire SNaN_SN;
	reg SNaN_SP;
	assign Zero_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_zero_S && Mant_a_prenorm_zero_S : Zero_a_SP);
	assign Zero_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_zero_S && Mant_b_prenorm_zero_S : Zero_b_SP);
	assign Inf_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && Mant_a_prenorm_zero_S : Inf_a_SP);
	assign Inf_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && Mant_b_prenorm_zero_S : Inf_b_SP);
	assign NaN_a_SN = (Start_S && Ready_SI ? Exp_a_prenorm_Inf_NaN_S && ~Mant_a_prenorm_zero_S : NaN_a_SP);
	assign NaN_b_SN = (Start_S && Ready_SI ? Exp_b_prenorm_Inf_NaN_S && ~Mant_b_prenorm_zero_S : NaN_b_SP);
	assign SNaN_SN = (Start_S && Ready_SI ? (Mant_a_prenorm_SNaN_S && NaN_a_SN) | (Mant_b_prenorm_SNaN_S && NaN_b_SN) : SNaN_SP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI) begin
			Zero_a_SP <= 1'sb0;
			Zero_b_SP <= 1'sb0;
			Inf_a_SP <= 1'sb0;
			Inf_b_SP <= 1'sb0;
			NaN_a_SP <= 1'sb0;
			NaN_b_SP <= 1'sb0;
			SNaN_SP <= 1'sb0;
		end
		else begin
			Inf_a_SP <= Inf_a_SN;
			Inf_b_SP <= Inf_b_SN;
			Zero_a_SP <= Zero_a_SN;
			Zero_b_SP <= Zero_b_SN;
			NaN_a_SP <= NaN_a_SN;
			NaN_b_SP <= NaN_b_SN;
			SNaN_SP <= SNaN_SN;
		end
	assign Special_case_SBO = ~{(Div_start_SI ? ((((Zero_a_SN | Zero_b_SN) | Inf_a_SN) | Inf_b_SN) | NaN_a_SN) | NaN_b_SN : ((Zero_a_SN | Inf_a_SN) | NaN_a_SN) | Sign_a_D)} && (Start_S && Ready_SI);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Special_case_dly_SBO <= 1'sb0;
		else if (Start_S && Ready_SI)
			Special_case_dly_SBO <= Special_case_SBO;
		else if (Special_case_dly_SBO)
			Special_case_dly_SBO <= 1'b1;
		else
			Special_case_dly_SBO <= 1'sb0;
	reg Sign_z_DN;
	reg Sign_z_DP;
	always @(*)
		if (Div_start_SI && Ready_SI)
			Sign_z_DN = Sign_a_D ^ Sign_b_D;
		else if (Sqrt_start_SI && Ready_SI)
			Sign_z_DN = Sign_a_D;
		else
			Sign_z_DN = Sign_z_DP;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Sign_z_DP <= 1'sb0;
		else
			Sign_z_DP <= Sign_z_DN;
	reg [2:0] RM_DN;
	reg [2:0] RM_DP;
	always @(*)
		if (Start_S && Ready_SI)
			RM_DN = RM_SI;
		else
			RM_DN = RM_DP;
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			RM_DP <= 1'sb0;
		else
			RM_DP <= RM_DN;
	assign RM_dly_SO = RM_DP;
	wire [5:0] Mant_leadingOne_a;
	wire [5:0] Mant_leadingOne_b;
	wire Mant_zero_S_a;
	wire Mant_zero_S_b;
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ua(
		.in_i(Mant_a_D),
		.cnt_o(Mant_leadingOne_a),
		.empty_o(Mant_zero_S_a)
	);
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_a_norm_DP;
	assign Mant_a_norm_DN = (Start_S && Ready_SI ? Mant_a_D << Mant_leadingOne_a : Mant_a_norm_DP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Mant_a_norm_DP <= 1'sb0;
		else
			Mant_a_norm_DP <= Mant_a_norm_DN;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_a_norm_DP;
	assign Exp_a_norm_DN = (Start_S && Ready_SI ? (Exp_a_D - Mant_leadingOne_a) + |Mant_leadingOne_a : Exp_a_norm_DP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Exp_a_norm_DP <= 1'sb0;
		else
			Exp_a_norm_DP <= Exp_a_norm_DN;
	lzc #(
		.WIDTH(53),
		.MODE(1)
	) LOD_Ub(
		.in_i(Mant_b_D),
		.cnt_o(Mant_leadingOne_b),
		.empty_o(Mant_zero_S_b)
	);
	wire [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_MANT_FP64:0] Mant_b_norm_DP;
	assign Mant_b_norm_DN = (Start_S && Ready_SI ? Mant_b_D << Mant_leadingOne_b : Mant_b_norm_DP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Mant_b_norm_DP <= 1'sb0;
		else
			Mant_b_norm_DP <= Mant_b_norm_DN;
	wire [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DN;
	reg [defs_div_sqrt_mvp_C_EXP_FP64:0] Exp_b_norm_DP;
	assign Exp_b_norm_DN = (Start_S && Ready_SI ? (Exp_b_D - Mant_leadingOne_b) + |Mant_leadingOne_b : Exp_b_norm_DP);
	always @(posedge Clk_CI or negedge Rst_RBI)
		if (~Rst_RBI)
			Exp_b_norm_DP <= 1'sb0;
		else
			Exp_b_norm_DP <= Exp_b_norm_DN;
	assign Start_SO = Start_S;
	assign Exp_a_DO_norm = Exp_a_norm_DP;
	assign Exp_b_DO_norm = Exp_b_norm_DP;
	assign Mant_a_DO_norm = Mant_a_norm_DP;
	assign Mant_b_DO_norm = Mant_b_norm_DP;
	assign Sign_z_DO = Sign_z_DP;
	assign Inf_a_SO = Inf_a_SP;
	assign Inf_b_SO = Inf_b_SP;
	assign Zero_a_SO = Zero_a_SP;
	assign Zero_b_SO = Zero_b_SP;
	assign NaN_a_SO = NaN_a_SP;
	assign NaN_b_SO = NaN_b_SP;
	assign SNaN_SO = SNaN_SP;
endmodule
module bht (
	clk_i,
	rst_ni,
	flush_i,
	debug_mode_i,
	vpc_i,
	bht_update_i,
	bht_prediction_o
);
	parameter [31:0] NR_ENTRIES = 1024;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire debug_mode_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] vpc_i;
	input wire [65:0] bht_update_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	localparam [31:0] ariane_pkg_INSTR_PER_FETCH = 2;
	output wire [3:0] bht_prediction_o;
	localparam OFFSET = 1;
	localparam NR_ROWS = NR_ENTRIES / ariane_pkg_INSTR_PER_FETCH;
	localparam ROW_ADDR_BITS = 1;
	localparam PREDICTION_BITS = ($clog2(NR_ROWS) + OFFSET) + ROW_ADDR_BITS;
	unread i_unread(.d_i(|vpc_i));
	reg [((NR_ROWS * ariane_pkg_INSTR_PER_FETCH) * 3) - 1:0] bht_d;
	reg [((NR_ROWS * ariane_pkg_INSTR_PER_FETCH) * 3) - 1:0] bht_q;
	wire [$clog2(NR_ROWS) - 1:0] index;
	wire [$clog2(NR_ROWS) - 1:0] update_pc;
	wire [0:0] update_row_index;
	reg [1:0] saturation_counter;
	assign index = vpc_i[PREDICTION_BITS - 1:2];
	assign update_pc = bht_update_i[0 + PREDICTION_BITS:3];
	assign update_row_index = bht_update_i[2:2];
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_bht_output
			assign bht_prediction_o[(i * 2) + 1] = bht_q[(((index * ariane_pkg_INSTR_PER_FETCH) + i) * 3) + 2];
			assign bht_prediction_o[i * 2] = bht_q[(((index * ariane_pkg_INSTR_PER_FETCH) + i) * 3) + 1] == 1'b1;
		end
	endgenerate
	always @(*) begin : update_bht
		bht_d = bht_q;
		saturation_counter = bht_q[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 1-:2];
		if (bht_update_i[65] && !debug_mode_i) begin
			bht_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 2] = 1'b1;
			if (saturation_counter == 2'b11) begin
				if (!bht_update_i[0])
					bht_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 1-:2] = saturation_counter - 1;
			end
			else if (saturation_counter == 2'b00) begin
				if (bht_update_i[0])
					bht_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 1-:2] = saturation_counter + 1;
			end
			else if (bht_update_i[0])
				bht_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 1-:2] = saturation_counter + 1;
			else
				bht_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 3) + 1-:2] = saturation_counter - 1;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < NR_ROWS; i = i + 1)
				begin : sv2v_autoblock_2
					reg signed [31:0] j;
					for (j = 0; j < ariane_pkg_INSTR_PER_FETCH; j = j + 1)
						bht_q[((i * ariane_pkg_INSTR_PER_FETCH) + j) * 3+:3] <= 1'sb0;
				end
		end
		else if (flush_i) begin : sv2v_autoblock_3
			reg signed [31:0] i;
			for (i = 0; i < NR_ROWS; i = i + 1)
				begin : sv2v_autoblock_4
					reg signed [31:0] j;
					for (j = 0; j < ariane_pkg_INSTR_PER_FETCH; j = j + 1)
						begin
							bht_q[(((i * ariane_pkg_INSTR_PER_FETCH) + j) * 3) + 2] <= 1'b0;
							bht_q[(((i * ariane_pkg_INSTR_PER_FETCH) + j) * 3) + 1-:2] <= 2'b10;
						end
				end
		end
		else
			bht_q <= bht_d;
endmodule
module btb (
	clk_i,
	rst_ni,
	flush_i,
	debug_mode_i,
	vpc_i,
	btb_update_i,
	btb_prediction_o
);
	parameter signed [31:0] NR_ENTRIES = 8;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire debug_mode_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] vpc_i;
	input wire [128:0] btb_update_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	localparam [31:0] ariane_pkg_INSTR_PER_FETCH = 2;
	output wire [129:0] btb_prediction_o;
	localparam OFFSET = 1;
	localparam NR_ROWS = NR_ENTRIES / ariane_pkg_INSTR_PER_FETCH;
	localparam ROW_ADDR_BITS = 1;
	localparam PREDICTION_BITS = ($clog2(NR_ROWS) + OFFSET) + ROW_ADDR_BITS;
	localparam ANTIALIAS_BITS = 8;
	unread i_unread(.d_i(|vpc_i));
	reg [((NR_ROWS * ariane_pkg_INSTR_PER_FETCH) * 65) - 1:0] btb_d;
	reg [((NR_ROWS * ariane_pkg_INSTR_PER_FETCH) * 65) - 1:0] btb_q;
	wire [$clog2(NR_ROWS) - 1:0] index;
	wire [$clog2(NR_ROWS) - 1:0] update_pc;
	wire [0:0] update_row_index;
	assign index = vpc_i[PREDICTION_BITS - 1:2];
	assign update_pc = btb_update_i[63 + PREDICTION_BITS:66];
	assign update_row_index = btb_update_i[65:65];
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_btb_output
			assign btb_prediction_o[i * 65+:65] = btb_q[((index * ariane_pkg_INSTR_PER_FETCH) + i) * 65+:65];
		end
	endgenerate
	always @(*) begin : update_branch_predict
		btb_d = btb_q;
		if (btb_update_i[128] && !debug_mode_i) begin
			btb_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 65) + 64] = 1'b1;
			btb_d[(((update_pc * ariane_pkg_INSTR_PER_FETCH) + update_row_index) * 65) + 63-:riscv_VLEN] = btb_update_i[63-:riscv_VLEN];
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < NR_ROWS; i = i + 1)
				btb_q[65 * (i * ariane_pkg_INSTR_PER_FETCH)+:130] <= {ariane_pkg_INSTR_PER_FETCH {65'd0}};
		end
		else if (flush_i) begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < NR_ROWS; i = i + 1)
				begin : sv2v_autoblock_3
					reg signed [31:0] j;
					for (j = 0; j < ariane_pkg_INSTR_PER_FETCH; j = j + 1)
						btb_q[(((i * ariane_pkg_INSTR_PER_FETCH) + j) * 65) + 64] <= 1'b0;
				end
		end
		else
			btb_q <= btb_d;
endmodule
module frontend (
	clk_i,
	rst_ni,
	flush_i,
	flush_bp_i,
	debug_mode_i,
	boot_addr_i,
	resolved_branch_i,
	set_pc_commit_i,
	pc_commit_i,
	epc_i,
	eret_i,
	trap_vector_base_i,
	ex_valid_i,
	set_debug_pc_i,
	icache_dreq_o,
	icache_dreq_i,
	fetch_entry_o,
	fetch_entry_valid_o,
	fetch_entry_ready_i
);
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire flush_bp_i;
	input wire debug_mode_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] boot_addr_i;
	input wire [133:0] resolved_branch_i;
	input wire set_pc_commit_i;
	input wire [63:0] pc_commit_i;
	input wire [63:0] epc_i;
	input wire eret_i;
	input wire [63:0] trap_vector_base_i;
	input wire ex_valid_i;
	input wire set_debug_pc_i;
	output reg [67:0] icache_dreq_o;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	input wire [226:0] icache_dreq_i;
	output wire [291:0] fetch_entry_o;
	output wire fetch_entry_valid_o;
	input wire fetch_entry_ready_i;
	reg [31:0] icache_data_q;
	reg icache_valid_q;
	reg [1:0] icache_ex_valid_q;
	reg [63:0] icache_vaddr_q;
	wire instr_queue_ready;
	localparam [31:0] ariane_pkg_INSTR_PER_FETCH = 2;
	wire [1:0] instr_queue_consumed;
	reg [64:0] btb_q;
	reg [1:0] bht_q;
	wire if_ready;
	reg [63:0] npc_d;
	reg [63:0] npc_q;
	reg npc_rst_load_q;
	wire replay;
	wire [63:0] replay_addr;
	wire [0:0] shamt;
	assign shamt = icache_dreq_i[130:130];
	wire [1:0] rvi_return;
	wire [1:0] rvi_call;
	wire [1:0] rvi_branch;
	wire [1:0] rvi_jalr;
	wire [1:0] rvi_jump;
	wire [127:0] rvi_imm;
	wire [1:0] rvc_branch;
	wire [1:0] rvc_jump;
	wire [1:0] rvc_jr;
	wire [1:0] rvc_return;
	wire [1:0] rvc_jalr;
	wire [1:0] rvc_call;
	wire [127:0] rvc_imm;
	wire [63:0] instr;
	wire [127:0] addr;
	wire [1:0] instruction_valid;
	wire [3:0] bht_prediction;
	wire [129:0] btb_prediction;
	wire [3:0] bht_prediction_shifted;
	wire [129:0] btb_prediction_shifted;
	wire [64:0] ras_predict;
	wire is_mispredict;
	reg ras_push;
	reg ras_pop;
	reg [63:0] ras_update;
	reg [63:0] predict_address;
	reg [5:0] cf_type;
	reg [1:0] taken_rvi_cf;
	reg [1:0] taken_rvc_cf;
	wire serving_unaligned;
	instr_realign i_instr_realign(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(icache_dreq_o[65]),
		.valid_i(icache_valid_q),
		.serving_unaligned_o(serving_unaligned),
		.address_i(icache_vaddr_q),
		.data_i(icache_data_q),
		.valid_o(instruction_valid),
		.addr_o(addr),
		.instr_o(instr)
	);
	assign bht_prediction_shifted[0+:2] = (serving_unaligned ? bht_q : bht_prediction[0+:2]);
	assign btb_prediction_shifted[0+:65] = (serving_unaligned ? btb_q : btb_prediction[0+:65]);
	genvar i;
	generate
		for (i = 1; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_prediction_address
			assign bht_prediction_shifted[i * 2+:2] = bht_prediction[addr[(i * 64) + 1-:1] * 2+:2];
			assign btb_prediction_shifted[i * 65+:65] = btb_prediction[addr[(i * 64) + 1-:1] * 65+:65];
		end
	endgenerate
	reg bp_valid;
	wire [1:0] is_branch;
	wire [1:0] is_call;
	wire [1:0] is_jump;
	wire [1:0] is_return;
	wire [1:0] is_jalr;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : genblk2
			assign is_branch[i] = instruction_valid[i] & (rvi_branch[i] | rvc_branch[i]);
			assign is_call[i] = instruction_valid[i] & (rvi_call[i] | rvc_call[i]);
			assign is_return[i] = instruction_valid[i] & (rvi_return[i] | rvc_return[i]);
			assign is_jump[i] = instruction_valid[i] & (rvi_jump[i] | rvc_jump[i]);
			assign is_jalr[i] = ((instruction_valid[i] & ~is_return[i]) & ~is_call[i]) & ((rvi_jalr[i] | rvc_jalr[i]) | rvc_jr[i]);
		end
	endgenerate
	always @(*) begin
		taken_rvi_cf = 1'sb0;
		taken_rvc_cf = 1'sb0;
		predict_address = 1'sb0;
		begin : sv2v_autoblock_1
			reg signed [31:0] i;
			for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1)
				cf_type[i * 3+:3] = 3'd0;
		end
		ras_push = 1'b0;
		ras_pop = 1'b0;
		ras_update = 1'sb0;
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 1; i >= 0; i = i - 1)
				begin
					case ({is_branch[i], is_return[i], is_jump[i], is_jalr[i]})
						4'b0000:
							;
						4'b0001: begin
							ras_pop = 1'b0;
							ras_push = 1'b0;
							if (btb_prediction_shifted[(i * 65) + 64]) begin
								predict_address = btb_prediction_shifted[(i * 65) + 63-:riscv_VLEN];
								cf_type[i * 3+:3] = 3'd3;
							end
						end
						4'b0010: begin
							ras_pop = 1'b0;
							ras_push = 1'b0;
							taken_rvi_cf[i] = rvi_jump[i];
							taken_rvc_cf[i] = rvc_jump[i];
							cf_type[i * 3+:3] = 3'd2;
						end
						4'b0100: begin
							ras_pop = ras_predict[64] & instr_queue_consumed[i];
							ras_push = 1'b0;
							predict_address = ras_predict[63-:riscv_VLEN];
							cf_type[i * 3+:3] = 3'd4;
						end
						4'b1000: begin
							ras_pop = 1'b0;
							ras_push = 1'b0;
							if (bht_prediction_shifted[(i * 2) + 1]) begin
								taken_rvi_cf[i] = rvi_branch[i] & bht_prediction_shifted[i * 2];
								taken_rvc_cf[i] = rvc_branch[i] & bht_prediction_shifted[i * 2];
							end
							else begin
								taken_rvi_cf[i] = rvi_branch[i] & rvi_imm[(i * 64) + 63];
								taken_rvc_cf[i] = rvc_branch[i] & rvc_imm[(i * 64) + 63];
							end
							if (taken_rvi_cf[i] || taken_rvc_cf[i])
								cf_type[i * 3+:3] = 3'd1;
						end
						default:
							;
					endcase
					if (is_call[i]) begin
						ras_push = instr_queue_consumed[i];
						ras_update = addr[i * 64+:64] + (rvc_call[i] ? 2 : 4);
					end
					if (taken_rvc_cf[i] || taken_rvi_cf[i])
						predict_address = addr[i * 64+:64] + (taken_rvc_cf[i] ? rvc_imm[i * 64+:64] : rvi_imm[i * 64+:64]);
				end
		end
	end
	always @(*) begin
		bp_valid = 1'b0;
		begin : sv2v_autoblock_3
			reg signed [31:0] i;
			for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1)
				bp_valid = bp_valid | (((cf_type[i * 3+:3] != 3'd0) & (cf_type[i * 3+:3] != 3'd4)) | ((cf_type[i * 3+:3] == 3'd4) & ras_predict[64]));
		end
	end
	assign is_mispredict = resolved_branch_i[133] & resolved_branch_i[4];
	wire [1:1] sv2v_tmp_A26B3;
	assign sv2v_tmp_A26B3 = instr_queue_ready;
	always @(*) icache_dreq_o[67] = sv2v_tmp_A26B3;
	assign if_ready = icache_dreq_i[226] & instr_queue_ready;
	wire [1:1] sv2v_tmp_45F60;
	assign sv2v_tmp_45F60 = (is_mispredict | flush_i) | replay;
	always @(*) icache_dreq_o[66] = sv2v_tmp_45F60;
	wire [1:1] sv2v_tmp_E2C77;
	assign sv2v_tmp_E2C77 = icache_dreq_o[66] | bp_valid;
	always @(*) icache_dreq_o[65] = sv2v_tmp_E2C77;
	wire [65:0] bht_update;
	wire [128:0] btb_update;
	reg speculative_q;
	wire speculative_d;
	assign speculative_d = ((((speculative_q && !resolved_branch_i[133]) || |is_branch) || |is_return) || |is_jalr) && !flush_i;
	wire [1:1] sv2v_tmp_E032C;
	assign sv2v_tmp_E032C = speculative_d;
	always @(*) icache_dreq_o[64] = sv2v_tmp_E032C;
	assign bht_update[65] = resolved_branch_i[133] & (resolved_branch_i[2-:3] == 3'd1);
	assign bht_update[64-:64] = resolved_branch_i[132-:64];
	assign bht_update[0] = resolved_branch_i[3];
	assign btb_update[128] = (resolved_branch_i[133] & resolved_branch_i[4]) & (resolved_branch_i[2-:3] == 3'd3);
	assign btb_update[127-:64] = resolved_branch_i[132-:64];
	assign btb_update[63-:riscv_VLEN] = resolved_branch_i[68-:64];
	localparam [63:0] dm_HaltAddress = 64'h0000000000000800;
	always @(*) begin : npc_select
		reg [63:0] fetch_address;
		if (npc_rst_load_q) begin
			npc_d = boot_addr_i;
			fetch_address = boot_addr_i;
		end
		else begin
			fetch_address = npc_q;
			npc_d = npc_q;
		end
		if (bp_valid) begin
			fetch_address = predict_address;
			npc_d = predict_address;
		end
		if (if_ready)
			npc_d = {fetch_address[63:2], 2'b00} + 'h4;
		if (replay)
			npc_d = replay_addr;
		if (is_mispredict)
			npc_d = resolved_branch_i[68-:64];
		if (eret_i)
			npc_d = epc_i;
		if (ex_valid_i)
			npc_d = trap_vector_base_i;
		if (set_pc_commit_i)
			npc_d = pc_commit_i + {{61 {1'b0}}, 3'b100};
		if (set_debug_pc_i)
			npc_d = ArianeCfg[95:32] + dm_HaltAddress[63:0];
		icache_dreq_o[63-:riscv_VLEN] = fetch_address;
	end
	wire [31:0] icache_data;
	assign icache_data = icache_dreq_i[224-:32] >> {shamt, 4'b0000};
	localparam [63:0] riscv_INSTR_ACCESS_FAULT = 1;
	localparam [63:0] riscv_INSTR_PAGE_FAULT = 12;
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			npc_rst_load_q <= 1'b1;
			npc_q <= 1'sb0;
			speculative_q <= 1'sb0;
			icache_data_q <= 1'sb0;
			icache_valid_q <= 1'b0;
			icache_vaddr_q <= 'b0;
			icache_ex_valid_q <= 2'd0;
			btb_q <= 1'sb0;
			bht_q <= 1'sb0;
		end
		else begin
			npc_rst_load_q <= 1'b0;
			npc_q <= npc_d;
			speculative_q <= speculative_d;
			icache_valid_q <= icache_dreq_i[225];
			if (icache_dreq_i[225]) begin
				icache_data_q <= icache_data;
				icache_vaddr_q <= icache_dreq_i[192-:64];
				if (icache_dreq_i[128-:64] == riscv_INSTR_PAGE_FAULT)
					icache_ex_valid_q <= 2'd2;
				else if (icache_dreq_i[128-:64] == riscv_INSTR_ACCESS_FAULT)
					icache_ex_valid_q <= 2'd1;
				else
					icache_ex_valid_q <= 2'd0;
				btb_q <= btb_prediction[65+:65];
				bht_q <= bht_prediction[2+:2];
			end
		end
	ras #(.DEPTH($signed(ArianeCfg[6433-:32]))) i_ras(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_bp_i),
		.push_i(ras_push),
		.pop_i(ras_pop),
		.data_i(ras_update),
		.data_o(ras_predict)
	);
	btb #(.NR_ENTRIES($signed(ArianeCfg[6401-:32]))) i_btb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_bp_i),
		.debug_mode_i(debug_mode_i),
		.vpc_i(icache_vaddr_q),
		.btb_update_i(btb_update),
		.btb_prediction_o(btb_prediction)
	);
	bht #(.NR_ENTRIES($signed(ArianeCfg[6369-:32]))) i_bht(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_bp_i),
		.debug_mode_i(debug_mode_i),
		.vpc_i(icache_vaddr_q),
		.bht_update_i(bht_update),
		.bht_prediction_o(bht_prediction)
	);
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_instr_scan
			instr_scan i_instr_scan(
				.instr_i(instr[i * 32+:32]),
				.rvi_return_o(rvi_return[i]),
				.rvi_call_o(rvi_call[i]),
				.rvi_branch_o(rvi_branch[i]),
				.rvi_jalr_o(rvi_jalr[i]),
				.rvi_jump_o(rvi_jump[i]),
				.rvi_imm_o(rvi_imm[i * 64+:64]),
				.rvc_branch_o(rvc_branch[i]),
				.rvc_jump_o(rvc_jump[i]),
				.rvc_jr_o(rvc_jr[i]),
				.rvc_return_o(rvc_return[i]),
				.rvc_jalr_o(rvc_jalr[i]),
				.rvc_call_o(rvc_call[i]),
				.rvc_imm_o(rvc_imm[i * 64+:64])
			);
		end
	endgenerate
	instr_queue i_instr_queue(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.instr_i(instr),
		.addr_i(addr),
		.exception_i(icache_ex_valid_q),
		.exception_addr_i(icache_vaddr_q),
		.predict_address_i(predict_address),
		.cf_type_i(cf_type),
		.valid_i(instruction_valid),
		.consumed_o(instr_queue_consumed),
		.ready_o(instr_queue_ready),
		.replay_o(replay),
		.replay_addr_o(replay_addr),
		.fetch_entry_o(fetch_entry_o),
		.fetch_entry_valid_o(fetch_entry_valid_o),
		.fetch_entry_ready_i(fetch_entry_ready_i)
	);
endmodule
module instr_queue (
	clk_i,
	rst_ni,
	flush_i,
	instr_i,
	addr_i,
	valid_i,
	ready_o,
	consumed_o,
	exception_i,
	exception_addr_i,
	predict_address_i,
	cf_type_i,
	replay_o,
	replay_addr_o,
	fetch_entry_o,
	fetch_entry_valid_o,
	fetch_entry_ready_i
);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	localparam [31:0] ariane_pkg_INSTR_PER_FETCH = 2;
	input wire [63:0] instr_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [127:0] addr_i;
	input wire [1:0] valid_i;
	output wire ready_o;
	output wire [1:0] consumed_o;
	input wire [1:0] exception_i;
	input wire [63:0] exception_addr_i;
	input wire [63:0] predict_address_i;
	input wire [5:0] cf_type_i;
	output wire replay_o;
	output wire [63:0] replay_addr_o;
	output reg [291:0] fetch_entry_o;
	output wire fetch_entry_valid_o;
	input wire fetch_entry_ready_i;
	wire [0:0] branch_index;
	localparam [31:0] ariane_pkg_FETCH_FIFO_DEPTH = 4;
	wire [3:0] instr_queue_usage;
	wire [201:0] instr_data_in;
	wire [201:0] instr_data_out;
	wire [1:0] push_instr;
	wire [1:0] push_instr_fifo;
	reg [1:0] pop_instr;
	wire [1:0] instr_queue_full;
	wire [1:0] instr_queue_empty;
	wire instr_overflow;
	wire [1:0] address_queue_usage;
	wire [63:0] address_out;
	wire pop_address;
	reg push_address;
	wire full_address;
	wire empty_address;
	wire address_overflow;
	wire [0:0] idx_is_d;
	reg [0:0] idx_is_q;
	reg [1:0] idx_ds_d;
	reg [1:0] idx_ds_q;
	reg [63:0] pc_d;
	reg [63:0] pc_q;
	reg reset_address_d;
	reg reset_address_q;
	wire [2:0] branch_mask_extended;
	wire [1:0] branch_mask;
	wire branch_empty;
	wire [1:0] taken;
	wire [1:0] popcount;
	wire [0:0] shamt;
	wire [1:0] valid;
	wire [3:0] consumed_extended;
	wire [3:0] fifo_pos_extended;
	wire [1:0] fifo_pos;
	wire [127:0] instr;
	wire [11:0] cf;
	wire [1:0] instr_overflow_fifo;
	assign ready_o = ~(|instr_queue_full) & ~full_address;
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_unpack_taken
			assign taken[i] = cf_type_i[i * 3+:3] != 3'd0;
		end
	endgenerate
	lzc #(
		.WIDTH(ariane_pkg_INSTR_PER_FETCH),
		.MODE(0)
	) i_lzc_branch_index(
		.in_i(taken),
		.cnt_o(branch_index),
		.empty_o(branch_empty)
	);
	assign branch_mask_extended = {1'b0, {{ariane_pkg_INSTR_PER_FETCH} {1'b1}}} << branch_index;
	assign branch_mask = branch_mask_extended[2:1];
	assign valid = valid_i & branch_mask;
	assign consumed_extended = {push_instr_fifo, push_instr_fifo} >> idx_is_q;
	assign consumed_o = consumed_extended[1:0];
	popcount #(.INPUT_WIDTH(ariane_pkg_INSTR_PER_FETCH)) i_popcount(
		.data_i(push_instr_fifo),
		.popcount_o(popcount)
	);
	assign shamt = popcount[0:0];
	assign idx_is_d = idx_is_q + shamt;
	assign fifo_pos_extended = {valid, valid} << idx_is_q;
	assign fifo_pos = fifo_pos_extended[3:ariane_pkg_INSTR_PER_FETCH];
	assign push_instr = fifo_pos & ~instr_queue_full;
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_duplicate_instr_input
			assign instr[i * 32+:32] = instr_i[i * 32+:32];
			assign instr[(i + ariane_pkg_INSTR_PER_FETCH) * 32+:32] = instr_i[i * 32+:32];
			assign cf[i * 3+:3] = cf_type_i[i * 3+:3];
			assign cf[(i + ariane_pkg_INSTR_PER_FETCH) * 3+:3] = cf_type_i[i * 3+:3];
		end
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_fifo_input_select
			assign instr_data_in[(i * 101) + 100-:32] = instr[(i + idx_is_q) * 32+:32];
			assign instr_data_in[(i * 101) + 68-:3] = cf[(i + idx_is_q) * 3+:3];
			assign instr_data_in[(i * 101) + 65-:2] = exception_i;
			assign instr_data_in[(i * 101) + 63-:riscv_VLEN] = exception_addr_i;
		end
	endgenerate
	assign instr_overflow_fifo = instr_queue_full & fifo_pos;
	assign instr_overflow = |instr_overflow_fifo;
	assign address_overflow = full_address & push_address;
	assign replay_o = instr_overflow | address_overflow;
	assign replay_addr_o = (address_overflow ? addr_i[0+:64] : addr_i[shamt * 64+:64]);
	assign fetch_entry_valid_o = ~(&instr_queue_empty);
	localparam [63:0] riscv_INSTR_ACCESS_FAULT = 1;
	localparam [63:0] riscv_INSTR_PAGE_FAULT = 12;
	always @(*) begin
		idx_ds_d = idx_ds_q;
		pop_instr = 1'sb0;
		fetch_entry_o[227-:32] = 1'sb0;
		fetch_entry_o[291-:64] = pc_q;
		fetch_entry_o[0] = 1'b0;
		fetch_entry_o[128-:64] = 1'sb0;
		fetch_entry_o[64-:64] = 1'sb0;
		fetch_entry_o[192-:riscv_VLEN] = address_out;
		fetch_entry_o[195-:3] = 3'd0;
		begin : sv2v_autoblock_1
			reg [31:0] i;
			for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1)
				if (idx_ds_q[i]) begin
					if (instr_data_out[(i * 101) + 65-:2] == 2'd1)
						fetch_entry_o[128-:64] = riscv_INSTR_ACCESS_FAULT;
					else
						fetch_entry_o[128-:64] = riscv_INSTR_PAGE_FAULT;
					fetch_entry_o[227-:32] = instr_data_out[(i * 101) + 100-:32];
					fetch_entry_o[0] = instr_data_out[(i * 101) + 65-:2] != 2'd0;
					fetch_entry_o[64-:64] = {instr_data_out[(i * 101) + 63-:riscv_VLEN]};
					fetch_entry_o[195-:3] = instr_data_out[(i * 101) + 68-:3];
					pop_instr[i] = fetch_entry_valid_o & fetch_entry_ready_i;
				end
		end
		if (fetch_entry_ready_i)
			idx_ds_d = {idx_ds_q[0:0], idx_ds_q[1]};
	end
	assign pop_address = (fetch_entry_o[195-:3] != 3'd0) & |pop_instr;
	always @(*) begin
		pc_d = pc_q;
		reset_address_d = (flush_i ? 1'b1 : reset_address_q);
		if (fetch_entry_ready_i)
			pc_d = pc_q + (fetch_entry_o[197:196] != 2'b11 ? 'd2 : 'd4);
		if (pop_address)
			pc_d = address_out;
		if (valid_i[0] && reset_address_q) begin
			pc_d = addr_i[0+:64];
			reset_address_d = 1'b0;
		end
	end
	generate
		for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1) begin : gen_instr_fifo
			assign push_instr_fifo[i] = push_instr[i] & ~address_overflow;
			fifo_v3_AECA2_3F763 #(
				.dtype_riscv_VLEN(riscv_VLEN),
				.DEPTH(ariane_pkg_FETCH_FIFO_DEPTH)
			) i_fifo_instr_data(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.testmode_i(1'b0),
				.full_o(instr_queue_full[i]),
				.empty_o(instr_queue_empty[i]),
				.usage_o(instr_queue_usage[i * 2+:2]),
				.data_i(instr_data_in[i * 101+:101]),
				.push_i(push_instr_fifo[i]),
				.data_o(instr_data_out[i * 101+:101]),
				.pop_i(pop_instr[i])
			);
		end
	endgenerate
	always @(*) begin
		push_address = 1'b0;
		begin : sv2v_autoblock_2
			reg signed [31:0] i;
			for (i = 0; i < ariane_pkg_INSTR_PER_FETCH; i = i + 1)
				push_address = push_address | (push_instr[i] & (instr_data_in[(i * 101) + 68-:3] != 3'd0));
		end
	end
	fifo_v3 #(
		.DEPTH(ariane_pkg_FETCH_FIFO_DEPTH),
		.DATA_WIDTH(riscv_VLEN)
	) i_fifo_address(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(flush_i),
		.testmode_i(1'b0),
		.full_o(full_address),
		.empty_o(empty_address),
		.usage_o(address_queue_usage),
		.data_i(predict_address_i),
		.push_i(push_address & ~full_address),
		.data_o(address_out),
		.pop_i(pop_address)
	);
	unread i_unread_address_fifo(.d_i(|{empty_address, address_queue_usage}));
	unread i_unread_branch_mask(.d_i(|branch_mask_extended));
	unread i_unread_lzc(.d_i(|{branch_empty}));
	unread i_unread_fifo_pos(.d_i(|fifo_pos_extended));
	unread i_unread_instr_fifo(.d_i(|instr_queue_usage));
	always @(posedge clk_i or negedge rst_ni)
		if (!rst_ni) begin
			idx_ds_q <= 'b1;
			idx_is_q <= 1'sb0;
			pc_q <= 1'sb0;
			reset_address_q <= 1'b1;
		end
		else begin
			pc_q <= pc_d;
			reset_address_q <= reset_address_d;
			if (flush_i) begin
				idx_ds_q <= 'b1;
				idx_is_q <= 1'sb0;
				reset_address_q <= 1'b1;
			end
			else begin
				idx_ds_q <= idx_ds_d;
				idx_is_q <= idx_is_d;
			end
		end
endmodule
module instr_scan (
	instr_i,
	rvi_return_o,
	rvi_call_o,
	rvi_branch_o,
	rvi_jalr_o,
	rvi_jump_o,
	rvi_imm_o,
	rvc_branch_o,
	rvc_jump_o,
	rvc_jr_o,
	rvc_return_o,
	rvc_jalr_o,
	rvc_call_o,
	rvc_imm_o
);
	input wire [31:0] instr_i;
	output wire rvi_return_o;
	output wire rvi_call_o;
	output wire rvi_branch_o;
	output wire rvi_jalr_o;
	output wire rvi_jump_o;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	output wire [63:0] rvi_imm_o;
	output wire rvc_branch_o;
	output wire rvc_jump_o;
	output wire rvc_jr_o;
	output wire rvc_return_o;
	output wire rvc_jalr_o;
	output wire rvc_call_o;
	output wire [63:0] rvc_imm_o;
	wire is_rvc;
	assign is_rvc = instr_i[1:0] != 2'b11;
	wire rv32_rvc_jal;
	localparam riscv_OpcodeC1 = 2'b01;
	localparam riscv_OpcodeC1Jal = 3'b001;
	assign rv32_rvc_jal = 1'd0 & (((instr_i[15:13] == riscv_OpcodeC1Jal) & is_rvc) & (instr_i[1:0] == riscv_OpcodeC1));
	assign rvi_return_o = (rvi_jalr_o & ((instr_i[19:15] == 5'd1) | (instr_i[19:15] == 5'd5))) & (instr_i[19:15] != instr_i[11:7]);
	assign rvi_call_o = (rvi_jalr_o | rvi_jump_o) & ((instr_i[11:7] == 5'd1) | (instr_i[11:7] == 5'd5));
	function automatic [63:0] ariane_pkg_sb_imm;
		input reg [31:0] instruction_i;
		ariane_pkg_sb_imm = {{51 {instruction_i[31]}}, instruction_i[31], instruction_i[7], instruction_i[30:25], instruction_i[11:8], 1'b0};
	endfunction
	function automatic [63:0] ariane_pkg_uj_imm;
		input reg [31:0] instruction_i;
		ariane_pkg_uj_imm = {{44 {instruction_i[31]}}, instruction_i[19:12], instruction_i[20], instruction_i[30:21], 1'b0};
	endfunction
	assign rvi_imm_o = (instr_i[3] ? ariane_pkg_uj_imm(instr_i) : ariane_pkg_sb_imm(instr_i));
	localparam riscv_OpcodeBranch = 7'b1100011;
	assign rvi_branch_o = instr_i[6:0] == riscv_OpcodeBranch;
	localparam riscv_OpcodeJalr = 7'b1100111;
	assign rvi_jalr_o = instr_i[6:0] == riscv_OpcodeJalr;
	localparam riscv_OpcodeJal = 7'b1101111;
	assign rvi_jump_o = instr_i[6:0] == riscv_OpcodeJal;
	localparam riscv_OpcodeC1J = 3'b101;
	assign rvc_jump_o = (((instr_i[15:13] == riscv_OpcodeC1J) & is_rvc) & (instr_i[1:0] == riscv_OpcodeC1)) | rv32_rvc_jal;
	wire is_jal_r;
	localparam riscv_OpcodeC2 = 2'b10;
	localparam riscv_OpcodeC2JalrMvAdd = 3'b100;
	assign is_jal_r = (((instr_i[15:13] == riscv_OpcodeC2JalrMvAdd) & (instr_i[6:2] == 5'b00000)) & (instr_i[1:0] == riscv_OpcodeC2)) & is_rvc;
	assign rvc_jr_o = is_jal_r & ~instr_i[12];
	assign rvc_jalr_o = is_jal_r & instr_i[12];
	assign rvc_call_o = rvc_jalr_o | rv32_rvc_jal;
	localparam riscv_OpcodeC1Beqz = 3'b110;
	localparam riscv_OpcodeC1Bnez = 3'b111;
	assign rvc_branch_o = (((instr_i[15:13] == riscv_OpcodeC1Beqz) | (instr_i[15:13] == riscv_OpcodeC1Bnez)) & (instr_i[1:0] == riscv_OpcodeC1)) & is_rvc;
	assign rvc_return_o = ((instr_i[11:7] == 5'd1) | (instr_i[11:7] == 5'd5)) & rvc_jr_o;
	assign rvc_imm_o = (instr_i[14] ? {{56 {instr_i[12]}}, instr_i[6:5], instr_i[2], instr_i[11:10], instr_i[4:3], 1'b0} : {{53 {instr_i[12]}}, instr_i[8], instr_i[10:9], instr_i[6], instr_i[7], instr_i[2], instr_i[11], instr_i[5:3], 1'b0});
endmodule
module ras (
	clk_i,
	rst_ni,
	flush_i,
	push_i,
	pop_i,
	data_i,
	data_o
);
	parameter [31:0] DEPTH = 2;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire push_i;
	input wire pop_i;
	localparam riscv_XLEN = 64;
	localparam riscv_VLEN = 64;
	input wire [63:0] data_i;
	output wire [64:0] data_o;
	reg [(DEPTH * 65) - 1:0] stack_d;
	reg [(DEPTH * 65) - 1:0] stack_q;
	assign data_o = stack_q[0+:65];
	always @(*) begin
		stack_d = stack_q;
		if (push_i) begin
			stack_d[63-:riscv_VLEN] = data_i;
			stack_d[64] = 1'b1;
			stack_d[65 * (((DEPTH - 1) >= 1 ? DEPTH - 1 : ((DEPTH - 1) + ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH) - 1))+:65 * ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)] = stack_q[65 * (((DEPTH - 2) >= 0 ? DEPTH - 2 : ((DEPTH - 2) + ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH) - 1))+:65 * ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)];
		end
		if (pop_i) begin
			stack_d[65 * (((DEPTH - 2) >= 0 ? DEPTH - 2 : ((DEPTH - 2) + ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH) - 1))+:65 * ((DEPTH - 2) >= 0 ? DEPTH - 1 : 3 - DEPTH)] = stack_q[65 * (((DEPTH - 1) >= 1 ? DEPTH - 1 : ((DEPTH - 1) + ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)) - 1) - (((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH) - 1))+:65 * ((DEPTH - 1) >= 1 ? DEPTH - 1 : 3 - DEPTH)];
			stack_d[((DEPTH - 1) * 65) + 64] = 1'b0;
			stack_d[((DEPTH - 1) * 65) + 63-:riscv_VLEN] = 'b0;
		end
		if (pop_i && push_i) begin
			stack_d = stack_q;
			stack_d[63-:riscv_VLEN] = data_i;
			stack_d[64] = 1'b1;
		end
		if (flush_i)
			stack_d = 1'sb0;
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			stack_q <= 1'sb0;
		else
			stack_q <= stack_d;
endmodule
module cva6_icache (
	clk_i,
	rst_ni,
	flush_i,
	en_i,
	miss_o,
	areq_i,
	areq_o,
	dreq_i,
	dreq_o,
	mem_rtrn_vld_i,
	mem_rtrn_i,
	mem_data_req_o,
	mem_data_ack_i,
	mem_data_o
);
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	parameter [1:0] RdTxId = 0;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire en_i;
	output reg miss_o;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	input wire [185:0] areq_i;
	localparam riscv_VLEN = 64;
	output reg [64:0] areq_o;
	input wire [67:0] dreq_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	output reg [226:0] dreq_o;
	input wire mem_rtrn_vld_i;
	localparam [31:0] ariane_pkg_ICACHE_LINE_WIDTH = 128;
	localparam [31:0] ariane_pkg_ICACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	localparam wt_cache_pkg_L15_SET_ASSOC = ariane_pkg_DCACHE_SET_ASSOC;
	localparam wt_cache_pkg_L15_WAY_WIDTH = 3;
	input wire [147:0] mem_rtrn_i;
	output reg mem_data_req_o;
	input wire mem_data_ack_i;
	localparam [31:0] ariane_pkg_ICACHE_SET_ASSOC = 4;
	output wire [60:0] mem_data_o;
	reg cache_en_d;
	reg cache_en_q;
	wire [63:0] vaddr_d;
	reg [63:0] vaddr_q;
	wire paddr_is_nc;
	wire [3:0] cl_hit;
	reg cache_rden;
	reg cache_wren;
	reg cmp_en_d;
	reg cmp_en_q;
	reg flush_d;
	reg flush_q;
	wire update_lfsr;
	wire [1:0] inv_way;
	wire [1:0] rnd_way;
	wire [1:0] repl_way;
	wire [3:0] repl_way_oh_d;
	reg [3:0] repl_way_oh_q;
	wire all_ways_valid;
	reg inv_en;
	wire inv_d;
	reg inv_q;
	reg flush_en;
	wire flush_done;
	localparam wt_cache_pkg_ICACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_ICACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_ICACHE_CL_IDX_WIDTH = 8;
	wire [7:0] flush_cnt_d;
	reg [7:0] flush_cnt_q;
	wire cl_we;
	wire [3:0] cl_req;
	wire [7:0] cl_index;
	wire [3:0] cl_offset_d;
	reg [3:0] cl_offset_q;
	localparam [31:0] ariane_pkg_ICACHE_TAG_WIDTH = 44;
	wire [43:0] cl_tag_d;
	reg [43:0] cl_tag_q;
	wire [43:0] cl_tag_rdata [3:0];
	wire [127:0] cl_rdata [3:0];
	wire [(ariane_pkg_ICACHE_SET_ASSOC * ariane_pkg_FETCH_WIDTH) - 1:0] cl_sel;
	wire [3:0] vld_req;
	wire vld_we;
	wire [3:0] vld_wdata;
	wire [3:0] vld_rdata;
	wire [7:0] vld_addr;
	reg [2:0] state_d;
	reg [2:0] state_q;
	assign cl_tag_d = (areq_i[185] ? areq_i[128 + (ariane_pkg_ICACHE_TAG_WIDTH + ariane_pkg_ICACHE_INDEX_WIDTH):141] : cl_tag_q);
	function automatic ariane_pkg_range_check;
		input reg [63:0] base;
		input reg [63:0] len;
		input reg [63:0] address;
		ariane_pkg_range_check = (address >= base) && (address < (base + len));
	endfunction
	function automatic ariane_pkg_is_inside_cacheable_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_1
				reg [31:0] k;
				for (k = 0; k < Cfg[2177-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[1122 + (k * 64)+:64], Cfg[98 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_cacheable_regions = |pass;
		end
	endfunction
	assign paddr_is_nc = ~cache_en_q | ~ariane_pkg_is_inside_cacheable_regions(ArianeCfg, {{'d8 {1'b0}}, cl_tag_d, {ariane_pkg_ICACHE_INDEX_WIDTH {1'b0}}});
	wire [129:1] sv2v_tmp_CBB03;
	assign sv2v_tmp_CBB03 = areq_i[128-:129];
	always @(*) dreq_o[128-:129] = sv2v_tmp_CBB03;
	assign vaddr_d = (dreq_o[226] & dreq_i[67] ? dreq_i[63-:riscv_VLEN] : vaddr_q);
	wire [64:1] sv2v_tmp_70A69;
	assign sv2v_tmp_70A69 = {vaddr_q >> 2, 2'b00};
	always @(*) areq_o[63-:riscv_VLEN] = sv2v_tmp_70A69;
	assign cl_index = vaddr_d[11:wt_cache_pkg_ICACHE_OFFSET_WIDTH];
	generate
		if (ArianeCfg[97]) begin : gen_axi_offset
			assign cl_offset_d = (dreq_o[226] & dreq_i[67] ? {dreq_i[63-:riscv_VLEN] >> 2, 2'b00} : (paddr_is_nc & mem_data_req_o ? cl_offset_q[2] << 2 : cl_offset_q));
			assign mem_data_o[58-:56] = (paddr_is_nc ? {cl_tag_d, vaddr_q[11:3], 3'b000} : {cl_tag_d, vaddr_q[11:wt_cache_pkg_ICACHE_OFFSET_WIDTH], {wt_cache_pkg_ICACHE_OFFSET_WIDTH {1'b0}}});
		end
		else begin : gen_piton_offset
			assign cl_offset_d = (dreq_o[226] & dreq_i[67] ? {dreq_i[63-:riscv_VLEN] >> 2, 2'b00} : cl_offset_q);
			assign mem_data_o[58-:56] = (paddr_is_nc ? {cl_tag_d, vaddr_q[11:2], 2'b00} : {cl_tag_d, vaddr_q[11:wt_cache_pkg_ICACHE_OFFSET_WIDTH], {wt_cache_pkg_ICACHE_OFFSET_WIDTH {1'b0}}});
		end
	endgenerate
	assign mem_data_o[1-:wt_cache_pkg_CACHE_ID_WIDTH] = RdTxId;
	assign mem_data_o[2] = paddr_is_nc;
	assign mem_data_o[60-:2] = repl_way;
	wire [64:1] sv2v_tmp_97904;
	assign sv2v_tmp_97904 = vaddr_q;
	always @(*) dreq_o[192-:64] = sv2v_tmp_97904;
	assign inv_d = inv_en;
	wire addr_ni;
	function automatic ariane_pkg_is_inside_nonidempotent_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_2
				reg [31:0] k;
				for (k = 0; k < Cfg[6337-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[5282 + (k * 64)+:64], Cfg[4258 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_nonidempotent_regions = |pass;
		end
	endfunction
	assign addr_ni = ariane_pkg_is_inside_nonidempotent_regions(ArianeCfg, areq_i[184-:56]);
	always @(*) begin : p_fsm
		state_d = state_q;
		cache_en_d = cache_en_q & en_i;
		flush_en = 1'b0;
		cmp_en_d = 1'b0;
		cache_rden = 1'b0;
		cache_wren = 1'b0;
		inv_en = 1'b0;
		flush_d = flush_q | flush_i;
		dreq_o[226] = 1'b0;
		areq_o[64] = 1'b0;
		dreq_o[225] = 1'b0;
		mem_data_req_o = 1'b0;
		miss_o = 1'b0;
		if (mem_rtrn_vld_i && (mem_rtrn_i[147] == 1'd0))
			inv_en = 1'b1;
		case (state_q)
			3'd0: begin
				flush_en = 1'b1;
				if (flush_done) begin
					state_d = 3'd1;
					flush_d = 1'b0;
					cache_en_d = en_i;
				end
			end
			3'd1: begin
				cmp_en_d = cache_en_q;
				if (flush_d || (en_i && !cache_en_q))
					state_d = 3'd0;
				else begin
					if (!mem_rtrn_vld_i) begin
						dreq_o[226] = 1'b1;
						if (dreq_i[67]) begin
							cache_rden = 1'b1;
							state_d = 3'd2;
						end
					end
					if (dreq_i[66])
						state_d = 3'd1;
				end
			end
			3'd2: begin
				areq_o[64] = 1'sb1;
				cmp_en_d = cache_en_q;
				cache_rden = cache_en_q;
				if (areq_i[185] && (!dreq_i[64] || !addr_ni)) begin
					if (flush_d)
						state_d = 3'd1;
					else if (((|cl_hit && cache_en_q) || areq_i[0]) && !inv_q) begin
						dreq_o[225] = ~dreq_i[65];
						state_d = 3'd1;
						if (!mem_rtrn_vld_i) begin
							dreq_o[226] = 1'b1;
							if (dreq_i[67])
								state_d = 3'd2;
						end
						if (dreq_i[66])
							state_d = 3'd1;
					end
					else if (dreq_i[65])
						state_d = 3'd1;
					else if (!inv_q) begin
						cmp_en_d = 1'b0;
						mem_data_req_o = 1'b1;
						if (mem_data_ack_i) begin
							miss_o = ~paddr_is_nc;
							state_d = 3'd3;
						end
					end
				end
				else if (dreq_i[65] || flush_d)
					state_d = 3'd4;
			end
			3'd3:
				if (mem_rtrn_vld_i && (mem_rtrn_i[147] == 1'd1)) begin
					state_d = 3'd1;
					if (!(dreq_i[65] || flush_d)) begin
						dreq_o[225] = 1'b1;
						cache_wren = ~paddr_is_nc;
					end
				end
				else if (dreq_i[65] || flush_d)
					state_d = 3'd5;
			3'd4: begin
				areq_o[64] = 1'sb1;
				if (areq_i[185])
					state_d = 3'd1;
			end
			3'd5:
				if (mem_rtrn_vld_i && (mem_rtrn_i[147] == 1'd1))
					state_d = 3'd1;
			default: state_d = 3'd0;
		endcase
	end
	assign flush_cnt_d = (flush_done ? {wt_cache_pkg_ICACHE_CL_IDX_WIDTH {1'sb0}} : (flush_en ? flush_cnt_q + 1 : flush_cnt_q));
	assign flush_done = flush_cnt_q == 255;
	assign vld_addr = (flush_en ? flush_cnt_q : (inv_en ? mem_rtrn_i[16:9] : cl_index));
	localparam wt_cache_pkg_L1I_WAY_WIDTH = 2;
	function automatic [3:0] wt_cache_pkg_icache_way_bin2oh;
		input reg [1:0] in;
		reg [3:0] out;
		begin
			out = 1'sb0;
			out[in] = 1'b1;
			wt_cache_pkg_icache_way_bin2oh = out;
		end
	endfunction
	assign vld_req = (flush_en || cache_rden ? {4 {1'sb1}} : (mem_rtrn_i[17] && inv_en ? {4 {1'sb1}} : (mem_rtrn_i[18] && inv_en ? wt_cache_pkg_icache_way_bin2oh(mem_rtrn_i[4-:wt_cache_pkg_L15_WAY_WIDTH]) : repl_way_oh_q)));
	assign vld_wdata = (cache_wren ? {4 {1'sb1}} : {4 {1'sb0}});
	assign vld_we = (cache_wren | inv_en) | flush_en;
	assign update_lfsr = cache_wren & all_ways_valid;
	assign repl_way = (all_ways_valid ? rnd_way : inv_way);
	assign repl_way_oh_d = (cmp_en_q ? wt_cache_pkg_icache_way_bin2oh(repl_way) : repl_way_oh_q);
	assign cl_req = (cache_rden ? {4 {1'sb1}} : (cache_wren ? repl_way_oh_q : {4 {1'sb0}}));
	assign cl_we = cache_wren;
	lzc #(.WIDTH(ariane_pkg_ICACHE_SET_ASSOC)) i_lzc(
		.in_i(~vld_rdata),
		.cnt_o(inv_way),
		.empty_o(all_ways_valid)
	);
	lfsr_8bit #(.WIDTH(ariane_pkg_ICACHE_SET_ASSOC)) i_lfsr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_i(update_lfsr),
		.refill_way_oh(),
		.refill_way_bin(rnd_way)
	);
	wire [1:0] hit_idx;
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_ICACHE_SET_ASSOC; i = i + 1) begin : gen_tag_cmpsel
			assign cl_hit[i] = (cl_tag_rdata[i] == cl_tag_d) & vld_rdata[i];
			assign cl_sel[i * ariane_pkg_FETCH_WIDTH+:ariane_pkg_FETCH_WIDTH] = cl_rdata[i][{cl_offset_q, 3'b000}+:ariane_pkg_FETCH_WIDTH];
		end
	endgenerate
	lzc #(.WIDTH(ariane_pkg_ICACHE_SET_ASSOC)) i_lzc_hit(
		.in_i(cl_hit),
		.cnt_o(hit_idx),
		.empty_o()
	);
	wire [32:1] sv2v_tmp_EAAF9;
	assign sv2v_tmp_EAAF9 = (cmp_en_q ? cl_sel[hit_idx * ariane_pkg_FETCH_WIDTH+:ariane_pkg_FETCH_WIDTH] : mem_rtrn_i[19 + {cl_offset_q, 3'b000}+:ariane_pkg_FETCH_WIDTH]);
	always @(*) dreq_o[224-:32] = sv2v_tmp_EAAF9;
	wire [ariane_pkg_ICACHE_TAG_WIDTH:0] cl_tag_valid_rdata [3:0];
	generate
		for (i = 0; i < ariane_pkg_ICACHE_SET_ASSOC; i = i + 1) begin : gen_sram
			localparam sv2v_uu_tag_sram_DATA_WIDTH = 45;
			localparam [5:0] sv2v_uu_tag_sram_ext_be_i_1 = 1'sb1;
			sram #(
				.DATA_WIDTH(45),
				.NUM_WORDS(wt_cache_pkg_ICACHE_NUM_WORDS)
			) tag_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(vld_req[i]),
				.we_i(vld_we),
				.addr_i(vld_addr),
				.wdata_i({vld_wdata[i], cl_tag_q}),
				.be_i(sv2v_uu_tag_sram_ext_be_i_1),
				.rdata_o(cl_tag_valid_rdata[i])
			);
			assign cl_tag_rdata[i] = cl_tag_valid_rdata[i][43:0];
			assign vld_rdata[i] = cl_tag_valid_rdata[i][ariane_pkg_ICACHE_TAG_WIDTH];
			localparam sv2v_uu_data_sram_DATA_WIDTH = ariane_pkg_ICACHE_LINE_WIDTH;
			localparam [15:0] sv2v_uu_data_sram_ext_be_i_1 = 1'sb1;
			sram #(
				.DATA_WIDTH(ariane_pkg_ICACHE_LINE_WIDTH),
				.NUM_WORDS(wt_cache_pkg_ICACHE_NUM_WORDS)
			) data_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(cl_req[i]),
				.we_i(cl_we),
				.addr_i(cl_index),
				.wdata_i(mem_rtrn_i[146-:128]),
				.be_i(sv2v_uu_data_sram_ext_be_i_1),
				.rdata_o(cl_rdata[i])
			);
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			cl_tag_q <= 1'sb0;
			flush_cnt_q <= 1'sb0;
			vaddr_q <= 1'sb0;
			cmp_en_q <= 1'sb0;
			cache_en_q <= 1'sb0;
			flush_q <= 1'sb0;
			state_q <= 3'd1;
			cl_offset_q <= 1'sb0;
			repl_way_oh_q <= 1'sb0;
			inv_q <= 1'sb0;
		end
		else begin
			cl_tag_q <= cl_tag_d;
			flush_cnt_q <= flush_cnt_d;
			vaddr_q <= vaddr_d;
			cmp_en_q <= cmp_en_d;
			cache_en_q <= cache_en_d;
			flush_q <= flush_d;
			state_q <= state_d;
			cl_offset_q <= cl_offset_d;
			repl_way_oh_q <= repl_way_oh_d;
			inv_q <= inv_d;
		end
	end
endmodule
module wt_dcache_wbuffer (
	clk_i,
	rst_ni,
	cache_en_i,
	empty_o,
	not_ni_o,
	req_port_i,
	req_port_o,
	miss_ack_i,
	miss_paddr_o,
	miss_req_o,
	miss_we_o,
	miss_wdata_o,
	miss_vld_bits_o,
	miss_nc_o,
	miss_size_o,
	miss_id_o,
	miss_rtrn_vld_i,
	miss_rtrn_id_i,
	rd_tag_o,
	rd_idx_o,
	rd_off_o,
	rd_req_o,
	rd_tag_only_o,
	rd_ack_i,
	rd_data_i,
	rd_vld_bits_i,
	rd_hit_oh_i,
	wr_cl_vld_i,
	wr_cl_idx_i,
	wr_req_o,
	wr_ack_i,
	wr_idx_o,
	wr_off_o,
	wr_data_o,
	wr_data_be_o,
	wbuffer_data_o,
	tx_paddr_o,
	tx_vld_o
);
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire cache_en_i;
	output wire empty_o;
	output wire not_ni_o;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	input wire [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_i;
	output reg [65:0] req_port_o;
	input wire miss_ack_i;
	output wire [55:0] miss_paddr_o;
	output wire miss_req_o;
	output wire miss_we_o;
	output wire [63:0] miss_wdata_o;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	output wire [7:0] miss_vld_bits_o;
	output wire miss_nc_o;
	output wire [2:0] miss_size_o;
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	output wire [1:0] miss_id_o;
	input wire miss_rtrn_vld_i;
	input wire [1:0] miss_rtrn_id_i;
	output wire [43:0] rd_tag_o;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	localparam wt_cache_pkg_DCACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_DCACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_DCACHE_CL_IDX_WIDTH = 8;
	output wire [7:0] rd_idx_o;
	output wire [3:0] rd_off_o;
	output wire rd_req_o;
	output wire rd_tag_only_o;
	input wire rd_ack_i;
	input wire [63:0] rd_data_i;
	input wire [7:0] rd_vld_bits_i;
	input wire [7:0] rd_hit_oh_i;
	input wire wr_cl_vld_i;
	input wire [7:0] wr_cl_idx_i;
	output reg [7:0] wr_req_o;
	input wire wr_ack_i;
	output wire [7:0] wr_idx_o;
	output wire [3:0] wr_off_o;
	output wire [63:0] wr_data_o;
	output wire [7:0] wr_data_be_o;
	localparam wt_cache_pkg_DCACHE_WBUF_DEPTH = 8;
	output wire [(8 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] wbuffer_data_o;
	localparam wt_cache_pkg_DCACHE_MAX_TX = 4;
	output wire [223:0] tx_paddr_o;
	output wire [3:0] tx_vld_o;
	reg [47:0] tx_stat_d;
	reg [47:0] tx_stat_q;
	reg [(8 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] wbuffer_d;
	reg [(8 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] wbuffer_q;
	wire [7:0] valid;
	wire [7:0] dirty;
	wire [7:0] tocheck;
	wire [7:0] wbuffer_hit_oh;
	wire [7:0] inval_hit;
	wire [63:0] bdirty;
	wire [2:0] next_ptr;
	wire [2:0] dirty_ptr;
	wire [2:0] hit_ptr;
	wire [2:0] wr_ptr;
	wire [2:0] check_ptr_d;
	reg [2:0] check_ptr_q;
	reg [2:0] check_ptr_q1;
	wire [2:0] rtrn_ptr;
	wire [1:0] tx_id;
	wire [1:0] rtrn_id;
	wire [2:0] bdirty_off;
	wire [7:0] tx_be;
	wire [55:0] wr_paddr;
	wire [55:0] rd_paddr;
	wire [43:0] rd_tag_d;
	reg [43:0] rd_tag_q;
	wire [7:0] rd_hit_oh_d;
	reg [7:0] rd_hit_oh_q;
	wire check_en_d;
	reg check_en_q;
	reg check_en_q1;
	wire full;
	reg dirty_rd_en;
	wire rdy;
	wire rtrn_empty;
	reg evict;
	reg [7:0] ni_pending_d;
	reg [7:0] ni_pending_q;
	reg wbuffer_wren;
	wire free_tx_slots;
	reg wr_cl_vld_q;
	wire wr_cl_vld_d;
	reg [7:0] wr_cl_idx_q;
	wire [7:0] wr_cl_idx_d;
	wire [55:0] debug_paddr [7:0];
	wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC) - 1:0] wbuffer_check_mux;
	wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC) - 1:0] wbuffer_dirty_mux;
	wire [43:0] miss_tag;
	wire is_nc_miss;
	wire is_ni;
	assign miss_tag = miss_paddr_o[ariane_pkg_DCACHE_INDEX_WIDTH+:ariane_pkg_DCACHE_TAG_WIDTH];
	function automatic ariane_pkg_range_check;
		input reg [63:0] base;
		input reg [63:0] len;
		input reg [63:0] address;
		ariane_pkg_range_check = (address >= base) && (address < (base + len));
	endfunction
	function automatic ariane_pkg_is_inside_cacheable_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_1
				reg [31:0] k;
				for (k = 0; k < Cfg[2177-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[1122 + (k * 64)+:64], Cfg[98 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_cacheable_regions = |pass;
		end
	endfunction
	assign is_nc_miss = !ariane_pkg_is_inside_cacheable_regions(ArianeCfg, {{20 {1'b0}}, miss_tag, {ariane_pkg_DCACHE_INDEX_WIDTH {1'b0}}});
	assign miss_nc_o = !cache_en_i || is_nc_miss;
	function automatic ariane_pkg_is_inside_nonidempotent_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_2
				reg [31:0] k;
				for (k = 0; k < Cfg[6337-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[5282 + (k * 64)+:64], Cfg[4258 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_nonidempotent_regions = |pass;
		end
	endfunction
	assign is_ni = ariane_pkg_is_inside_nonidempotent_regions(ArianeCfg, {{20 {1'b0}}, req_port_i[121-:44], {ariane_pkg_DCACHE_INDEX_WIDTH {1'b0}}});
	assign miss_we_o = 1'b1;
	assign miss_vld_bits_o = 1'sb0;
	assign wbuffer_data_o = wbuffer_q;
	genvar k;
	generate
		for (k = 0; k < wt_cache_pkg_DCACHE_MAX_TX; k = k + 1) begin : gen_tx_vld
			assign tx_vld_o[k] = tx_stat_q[(k * 12) + 11];
			assign tx_paddr_o[k * 56+:56] = wbuffer_q[(tx_stat_q[(k * 12) + 2-:3] * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] << 3;
		end
	endgenerate
	lzc #(.WIDTH(8)) i_vld_bdirty(
		.in_i(bdirty[dirty_ptr * 8+:8]),
		.cnt_o(bdirty_off),
		.empty_o()
	);
	assign miss_paddr_o = {wbuffer_dirty_mux[(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))], bdirty_off};
	assign miss_id_o = tx_id;
	assign miss_req_o = |dirty && free_tx_slots;
	function automatic [1:0] wt_cache_pkg_toSize64;
		input reg [7:0] be;
		reg [1:0] size;
		begin
			case (be)
				8'b11111111: size = 2'b11;
				8'b00001111, 8'b11110000: size = 2'b10;
				8'b11000000, 8'b00110000, 8'b00001100, 8'b00000011: size = 2'b01;
				default: size = 2'b00;
			endcase
			wt_cache_pkg_toSize64 = size;
		end
	endfunction
	assign miss_size_o = wt_cache_pkg_toSize64(bdirty[dirty_ptr * 8+:8]);
	function automatic [63:0] wt_cache_pkg_repData64;
		input reg [63:0] data;
		input reg [2:0] offset;
		input reg [1:0] size;
		reg [63:0] out;
		begin
			case (size)
				2'b00: begin : sv2v_autoblock_3
					reg signed [31:0] k;
					for (k = 0; k < 8; k = k + 1)
						out[k * 8+:8] = data[offset * 8+:8];
				end
				2'b01: begin : sv2v_autoblock_4
					reg signed [31:0] k;
					for (k = 0; k < 4; k = k + 1)
						out[k * 16+:16] = data[offset * 8+:16];
				end
				2'b10: begin : sv2v_autoblock_5
					reg signed [31:0] k;
					for (k = 0; k < 2; k = k + 1)
						out[k * 32+:32] = data[offset * 8+:32];
				end
				default: out = data;
			endcase
			wt_cache_pkg_repData64 = out;
		end
	endfunction
	assign miss_wdata_o = wt_cache_pkg_repData64(wbuffer_dirty_mux[96-:64], bdirty_off, miss_size_o[1:0]);
	function automatic [7:0] wt_cache_pkg_toByteEnable8;
		input reg [2:0] offset;
		input reg [1:0] size;
		reg [7:0] be;
		begin
			be = 1'sb0;
			case (size)
				2'b00: be[offset] = 1'sb1;
				2'b01: be[offset+:2] = 1'sb1;
				2'b10: be[offset+:4] = 1'sb1;
				default: be = 1'sb1;
			endcase
			wt_cache_pkg_toByteEnable8 = be;
		end
	endfunction
	assign tx_be = wt_cache_pkg_toByteEnable8(bdirty_off, miss_size_o[1:0]);
	fifo_v3 #(
		.FALL_THROUGH(1'b0),
		.DATA_WIDTH(2),
		.DEPTH(wt_cache_pkg_DCACHE_MAX_TX)
	) i_rtrn_id_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(),
		.empty_o(rtrn_empty),
		.usage_o(),
		.data_i(miss_rtrn_id_i),
		.push_i(miss_rtrn_vld_i),
		.data_o(rtrn_id),
		.pop_i(evict)
	);
	always @(*) begin : p_tx_stat
		tx_stat_d = tx_stat_q;
		evict = 1'b0;
		wr_req_o = 1'sb0;
		if (!rtrn_empty && wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8]) begin
			if (|wr_data_be_o && |wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 7-:ariane_pkg_DCACHE_SET_ASSOC]) begin
				wr_req_o = wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 7-:ariane_pkg_DCACHE_SET_ASSOC];
				if (wr_ack_i) begin
					evict = 1'b1;
					tx_stat_d[(rtrn_id * 12) + 11] = 1'b0;
				end
			end
			else begin
				evict = 1'b1;
				tx_stat_d[(rtrn_id * 12) + 11] = 1'b0;
			end
		end
		if (dirty_rd_en) begin
			tx_stat_d[(tx_id * 12) + 11] = 1'b1;
			tx_stat_d[(tx_id * 12) + 2-:3] = dirty_ptr;
			tx_stat_d[(tx_id * 12) + 10-:8] = tx_be;
		end
	end
	assign free_tx_slots = |(~tx_vld_o);
	localparam [0:0] sv2v_uu_i_tx_id_rr_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_tx_id_rr_NumIn = wt_cache_pkg_DCACHE_MAX_TX;
	localparam [1:0] sv2v_uu_i_tx_id_rr_ext_rr_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_tx_id_rr_DataWidth = 1;
	localparam [(sv2v_uu_i_tx_id_rr_NumIn * sv2v_uu_i_tx_id_rr_DataWidth) - 1:0] sv2v_uu_i_tx_id_rr_ext_data_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(wt_cache_pkg_DCACHE_MAX_TX),
		.LockIn(1'b1),
		.DataWidth(1)
	) i_tx_id_rr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_tx_id_rr_ext_flush_i_0),
		.rr_i(sv2v_uu_i_tx_id_rr_ext_rr_i_0),
		.req_i(~tx_vld_o),
		.gnt_o(),
		.data_i(sv2v_uu_i_tx_id_rr_ext_data_i_0),
		.gnt_i(dirty_rd_en),
		.req_o(),
		.data_o(),
		.idx_o(tx_id)
	);
	assign rd_tag_d = rd_paddr >> ariane_pkg_DCACHE_INDEX_WIDTH;
	assign rd_tag_only_o = 1'b1;
	assign rd_paddr = wbuffer_check_mux[(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] << 3;
	assign rd_req_o = |tocheck;
	assign rd_tag_o = rd_tag_q;
	assign rd_idx_o = rd_paddr[11:wt_cache_pkg_DCACHE_OFFSET_WIDTH];
	assign rd_off_o = rd_paddr[3:0];
	assign check_en_d = rd_req_o & rd_ack_i;
	assign rtrn_ptr = tx_stat_q[(rtrn_id * 12) + 2-:3];
	assign wr_data_be_o = tx_stat_q[(rtrn_id * 12) + 10-:8] & ~wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 32-:8];
	assign wr_paddr = wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] << 3;
	assign wr_idx_o = wr_paddr[11:wt_cache_pkg_DCACHE_OFFSET_WIDTH];
	assign wr_off_o = wr_paddr[3:0];
	assign wr_data_o = wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 96-:64];
	wire [63:0] wtag_comp;
	assign wr_cl_vld_d = wr_cl_vld_i;
	assign wr_cl_idx_d = wr_cl_idx_i;
	generate
		for (k = 0; k < wt_cache_pkg_DCACHE_WBUF_DEPTH; k = k + 1) begin : gen_flags
			assign debug_paddr[k] = wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] << 3;
			assign bdirty[k * 8+:8] = (|wbuffer_q[(k * ((32'd12 + 32'd44) + 97)) + 16-:8] ? {8 {1'sb0}} : wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 32-:8] & wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8]);
			assign dirty[k] = |bdirty[k * 8+:8];
			assign valid[k] = |wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8];
			assign wbuffer_hit_oh[k] = valid[k] & (wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] == {req_port_i[121-:44], req_port_i[133:125]});
			assign wtag_comp[k * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH] = wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 9)) >= (((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 2)) ? ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9) : ((((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9)) + ((((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 9)) >= (((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 2)) ? ((((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9)) - (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 2))) + 1 : ((((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 2)) - (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9))) + 1)) - 1)-:((((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 9)) >= (((32'd12 + 32'd44) + 96) - ((32'd12 + 32'd44) - 2)) ? ((((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9)) - (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 2))) + 1 : ((((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 2)) - (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) - 9))) + 1)];
			assign inval_hit[k] = ((wr_cl_vld_d & valid[k]) & (wtag_comp[k * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH] == wr_cl_idx_d)) | ((wr_cl_vld_q & valid[k]) & (wtag_comp[k * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH] == wr_cl_idx_q));
			assign tocheck[k] = ~wbuffer_q[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8] & valid[k];
		end
	endgenerate
	assign wr_ptr = (|wbuffer_hit_oh ? hit_ptr : next_ptr);
	assign rdy = |wbuffer_hit_oh | ~full;
	lzc #(.WIDTH(wt_cache_pkg_DCACHE_WBUF_DEPTH)) i_vld_lzc(
		.in_i(~valid),
		.cnt_o(next_ptr),
		.empty_o(full)
	);
	lzc #(.WIDTH(wt_cache_pkg_DCACHE_WBUF_DEPTH)) i_hit_lzc(
		.in_i(wbuffer_hit_oh),
		.cnt_o(hit_ptr),
		.empty_o()
	);
	localparam [0:0] sv2v_uu_i_dirty_rr_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_dirty_rr_NumIn = wt_cache_pkg_DCACHE_WBUF_DEPTH;
	localparam [2:0] sv2v_uu_i_dirty_rr_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_866BD_14B99 #(
		.DataType_ariane_pkg_DCACHE_INDEX_WIDTH(ariane_pkg_DCACHE_INDEX_WIDTH),
		.DataType_ariane_pkg_DCACHE_SET_ASSOC(ariane_pkg_DCACHE_SET_ASSOC),
		.DataType_ariane_pkg_DCACHE_TAG_WIDTH(ariane_pkg_DCACHE_TAG_WIDTH),
		.NumIn(wt_cache_pkg_DCACHE_WBUF_DEPTH),
		.LockIn(1'b1)
	) i_dirty_rr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_dirty_rr_ext_flush_i_0),
		.rr_i(sv2v_uu_i_dirty_rr_ext_rr_i_0),
		.req_i(dirty),
		.gnt_o(),
		.data_i(wbuffer_q),
		.gnt_i(dirty_rd_en),
		.req_o(),
		.data_o(wbuffer_dirty_mux),
		.idx_o(dirty_ptr)
	);
	localparam [0:0] sv2v_uu_i_clean_rr_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_clean_rr_NumIn = wt_cache_pkg_DCACHE_WBUF_DEPTH;
	localparam [2:0] sv2v_uu_i_clean_rr_ext_rr_i_0 = 1'sb0;
	rr_arb_tree_866BD_14B99 #(
		.DataType_ariane_pkg_DCACHE_INDEX_WIDTH(ariane_pkg_DCACHE_INDEX_WIDTH),
		.DataType_ariane_pkg_DCACHE_SET_ASSOC(ariane_pkg_DCACHE_SET_ASSOC),
		.DataType_ariane_pkg_DCACHE_TAG_WIDTH(ariane_pkg_DCACHE_TAG_WIDTH),
		.NumIn(wt_cache_pkg_DCACHE_WBUF_DEPTH)
	) i_clean_rr(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_clean_rr_ext_flush_i_0),
		.rr_i(sv2v_uu_i_clean_rr_ext_rr_i_0),
		.req_i(tocheck),
		.gnt_o(),
		.data_i(wbuffer_q),
		.gnt_i(check_en_d),
		.req_o(),
		.data_o(wbuffer_check_mux),
		.idx_o(check_ptr_d)
	);
	wire [1:1] sv2v_tmp_6DFA6;
	assign sv2v_tmp_6DFA6 = 1'sb0;
	always @(*) req_port_o[64] = sv2v_tmp_6DFA6;
	wire [64:1] sv2v_tmp_63D26;
	assign sv2v_tmp_63D26 = 1'sb0;
	always @(*) req_port_o[63-:64] = sv2v_tmp_63D26;
	assign rd_hit_oh_d = rd_hit_oh_i;
	wire ni_inside;
	wire ni_conflict;
	assign ni_inside = |ni_pending_q;
	assign ni_conflict = is_ni && ni_inside;
	assign not_ni_o = !ni_inside;
	assign empty_o = !(|valid);
	always @(*) begin : p_buffer
		wbuffer_d = wbuffer_q;
		ni_pending_d = ni_pending_q;
		dirty_rd_en = 1'b0;
		req_port_o[65] = 1'b0;
		wbuffer_wren = 1'b0;
		if (check_en_q1) begin
			if (wbuffer_q[(check_ptr_q1 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8]) begin
				wbuffer_d[(check_ptr_q1 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8] = 1'b1;
				wbuffer_d[(check_ptr_q1 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 7-:ariane_pkg_DCACHE_SET_ASSOC] = rd_hit_oh_q;
			end
		end
		begin : sv2v_autoblock_6
			reg signed [31:0] k;
			for (k = 0; k < wt_cache_pkg_DCACHE_WBUF_DEPTH; k = k + 1)
				if (inval_hit[k])
					wbuffer_d[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8] = 1'b0;
		end
		if (evict) begin
			begin : sv2v_autoblock_7
				reg signed [31:0] k;
				for (k = 0; k < 8; k = k + 1)
					if (tx_stat_q[(rtrn_id * 12) + (3 + k)]) begin
						wbuffer_d[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (9 + k)] = 1'b0;
						if (!wbuffer_q[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (25 + k)])
							wbuffer_d[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (17 + k)] = 1'b0;
					end
			end
			if (wbuffer_d[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8] == 0) begin
				wbuffer_d[(rtrn_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8] = 1'b0;
				ni_pending_d[rtrn_ptr] = 1'b0;
			end
		end
		if (miss_req_o && miss_ack_i) begin
			dirty_rd_en = 1'b1;
			begin : sv2v_autoblock_8
				reg signed [31:0] k;
				for (k = 0; k < 8; k = k + 1)
					if (tx_be[k]) begin
						wbuffer_d[(dirty_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (25 + k)] = 1'b0;
						wbuffer_d[(dirty_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (9 + k)] = 1'b1;
					end
			end
		end
		if (req_port_i[13] && rdy) begin
			if (!ni_conflict) begin
				wbuffer_wren = 1'b1;
				req_port_o[65] = 1'b1;
				ni_pending_d[wr_ptr] = is_ni;
				wbuffer_d[(wr_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 8] = 1'b0;
				wbuffer_d[(wr_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] = {req_port_i[121-:44], req_port_i[133:125]};
				begin : sv2v_autoblock_9
					reg signed [31:0] k;
					for (k = 0; k < 8; k = k + 1)
						if (req_port_i[4 + k]) begin
							wbuffer_d[(wr_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (17 + k)] = 1'b1;
							wbuffer_d[(wr_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (25 + k)] = 1'b1;
							wbuffer_d[(wr_ptr * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + (33 + (k * 8))+:8] = req_port_i[14 + (k * 8)+:8];
						end
				end
			end
		end
	end
	function automatic [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC) - 1:0] sv2v_cast_760D3;
		input reg [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC) - 1:0] inp;
		sv2v_cast_760D3 = inp;
	endfunction
	function automatic [11:0] sv2v_cast_78AC3;
		input reg [11:0] inp;
		sv2v_cast_78AC3 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			wbuffer_q <= {wt_cache_pkg_DCACHE_WBUF_DEPTH {sv2v_cast_760D3(1'sb0)}};
			tx_stat_q <= {wt_cache_pkg_DCACHE_MAX_TX {sv2v_cast_78AC3(1'sb0)}};
			ni_pending_q <= 1'sb0;
			check_ptr_q <= 1'sb0;
			check_ptr_q1 <= 1'sb0;
			check_en_q <= 1'sb0;
			check_en_q1 <= 1'sb0;
			rd_tag_q <= 1'sb0;
			rd_hit_oh_q <= 1'sb0;
			wr_cl_vld_q <= 1'sb0;
			wr_cl_idx_q <= 1'sb0;
		end
		else begin
			wbuffer_q <= wbuffer_d;
			tx_stat_q <= tx_stat_d;
			ni_pending_q <= ni_pending_d;
			check_ptr_q <= check_ptr_d;
			check_ptr_q1 <= check_ptr_q;
			check_en_q <= check_en_d;
			check_en_q1 <= check_en_q;
			rd_tag_q <= rd_tag_d;
			rd_hit_oh_q <= rd_hit_oh_d;
			wr_cl_vld_q <= wr_cl_vld_d;
			wr_cl_idx_q <= wr_cl_idx_d;
		end
	end
endmodule
module wt_dcache (
	clk_i,
	rst_ni,
	enable_i,
	flush_i,
	flush_ack_o,
	miss_o,
	wbuffer_empty_o,
	wbuffer_not_ni_o,
	amo_req_i,
	amo_resp_o,
	req_ports_i,
	req_ports_o,
	mem_rtrn_vld_i,
	mem_rtrn_i,
	mem_data_req_o,
	mem_data_ack_i,
	mem_data_o
);
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	parameter [1:0] RdAmoTxId = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire enable_i;
	input wire flush_i;
	output wire flush_ack_o;
	output wire miss_o;
	output wire wbuffer_empty_o;
	output wire wbuffer_not_ni_o;
	input wire [134:0] amo_req_i;
	output wire [64:0] amo_resp_o;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	input wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (3 * ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78)) - 1 : (3 * (1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 76)):(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)] req_ports_i;
	output wire [197:0] req_ports_o;
	input wire mem_rtrn_vld_i;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	localparam [31:0] ariane_pkg_ICACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	localparam wt_cache_pkg_L15_SET_ASSOC = ariane_pkg_DCACHE_SET_ASSOC;
	localparam wt_cache_pkg_L15_WAY_WIDTH = 3;
	input wire [149:0] mem_rtrn_i;
	output wire mem_data_req_o;
	input wire mem_data_ack_i;
	localparam wt_cache_pkg_L1D_WAY_WIDTH = 3;
	output wire [134:0] mem_data_o;
	localparam NumPorts = 3;
	wire cache_en;
	wire wr_cl_vld;
	wire wr_cl_nc;
	wire [7:0] wr_cl_we;
	wire [43:0] wr_cl_tag;
	localparam wt_cache_pkg_DCACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_DCACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_DCACHE_CL_IDX_WIDTH = 8;
	wire [7:0] wr_cl_idx;
	wire [3:0] wr_cl_off;
	wire [127:0] wr_cl_data;
	wire [15:0] wr_cl_data_be;
	wire [7:0] wr_vld_bits;
	wire [7:0] wr_req;
	wire wr_ack;
	wire [7:0] wr_idx;
	wire [3:0] wr_off;
	wire [63:0] wr_data;
	wire [7:0] wr_data_be;
	wire [2:0] miss_req;
	wire [2:0] miss_ack;
	wire [2:0] miss_nc;
	wire [2:0] miss_we;
	wire [191:0] miss_wdata;
	wire [167:0] miss_paddr;
	wire [23:0] miss_vld_bits;
	wire [8:0] miss_size;
	wire [5:0] miss_id;
	wire [2:0] miss_replay;
	wire [2:0] miss_rtrn_vld;
	wire [1:0] miss_rtrn_id;
	wire [2:0] rd_prio;
	wire [2:0] rd_tag_only;
	wire [2:0] rd_req;
	wire [2:0] rd_ack;
	wire [131:0] rd_tag;
	wire [23:0] rd_idx;
	wire [11:0] rd_off;
	wire [63:0] rd_data;
	wire [7:0] rd_vld_bits;
	wire [7:0] rd_hit_oh;
	localparam wt_cache_pkg_DCACHE_MAX_TX = 4;
	wire [223:0] tx_paddr;
	wire [3:0] tx_vld;
	localparam wt_cache_pkg_DCACHE_WBUF_DEPTH = 8;
	wire [(8 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] wbuffer_data;
	wt_dcache_missunit #(
		.Axi64BitCompliant(ArianeCfg[97]),
		.AmoTxId(RdAmoTxId),
		.NumPorts(NumPorts)
	) i_wt_dcache_missunit(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.enable_i(enable_i),
		.flush_i(flush_i),
		.flush_ack_o(flush_ack_o),
		.miss_o(miss_o),
		.wbuffer_empty_i(wbuffer_empty_o),
		.cache_en_o(cache_en),
		.amo_req_i(amo_req_i),
		.amo_resp_o(amo_resp_o),
		.miss_req_i(miss_req),
		.miss_ack_o(miss_ack),
		.miss_nc_i(miss_nc),
		.miss_we_i(miss_we),
		.miss_wdata_i(miss_wdata),
		.miss_paddr_i(miss_paddr),
		.miss_vld_bits_i(miss_vld_bits),
		.miss_size_i(miss_size),
		.miss_id_i(miss_id),
		.miss_replay_o(miss_replay),
		.miss_rtrn_vld_o(miss_rtrn_vld),
		.miss_rtrn_id_o(miss_rtrn_id),
		.tx_paddr_i(tx_paddr),
		.tx_vld_i(tx_vld),
		.wr_cl_vld_o(wr_cl_vld),
		.wr_cl_nc_o(wr_cl_nc),
		.wr_cl_we_o(wr_cl_we),
		.wr_cl_tag_o(wr_cl_tag),
		.wr_cl_idx_o(wr_cl_idx),
		.wr_cl_off_o(wr_cl_off),
		.wr_cl_data_o(wr_cl_data),
		.wr_cl_data_be_o(wr_cl_data_be),
		.wr_vld_bits_o(wr_vld_bits),
		.mem_rtrn_vld_i(mem_rtrn_vld_i),
		.mem_rtrn_i(mem_rtrn_i),
		.mem_data_req_o(mem_data_req_o),
		.mem_data_ack_i(mem_data_ack_i),
		.mem_data_o(mem_data_o)
	);
	genvar k;
	generate
		for (k = 0; k < 2; k = k + 1) begin : gen_rd_ports
			assign rd_prio[k] = 1'b1;
			wt_dcache_ctrl #(
				.RdTxId(RdAmoTxId),
				.ArianeCfg(ArianeCfg)
			) i_wt_dcache_ctrl(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.cache_en_i(cache_en),
				.req_port_i(req_ports_i[(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) + (k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)))+:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))]),
				.req_port_o(req_ports_o[k * 66+:66]),
				.miss_req_o(miss_req[k]),
				.miss_ack_i(miss_ack[k]),
				.miss_we_o(miss_we[k]),
				.miss_wdata_o(miss_wdata[k * 64+:64]),
				.miss_vld_bits_o(miss_vld_bits[k * ariane_pkg_DCACHE_SET_ASSOC+:ariane_pkg_DCACHE_SET_ASSOC]),
				.miss_paddr_o(miss_paddr[k * 56+:56]),
				.miss_nc_o(miss_nc[k]),
				.miss_size_o(miss_size[k * 3+:3]),
				.miss_id_o(miss_id[k * 2+:2]),
				.miss_replay_i(miss_replay[k]),
				.miss_rtrn_vld_i(miss_rtrn_vld[k]),
				.wr_cl_vld_i(wr_cl_vld),
				.rd_tag_o(rd_tag[k * ariane_pkg_DCACHE_TAG_WIDTH+:ariane_pkg_DCACHE_TAG_WIDTH]),
				.rd_idx_o(rd_idx[k * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH]),
				.rd_off_o(rd_off[k * wt_cache_pkg_DCACHE_OFFSET_WIDTH+:wt_cache_pkg_DCACHE_OFFSET_WIDTH]),
				.rd_req_o(rd_req[k]),
				.rd_tag_only_o(rd_tag_only[k]),
				.rd_ack_i(rd_ack[k]),
				.rd_data_i(rd_data),
				.rd_vld_bits_i(rd_vld_bits),
				.rd_hit_oh_i(rd_hit_oh)
			);
		end
	endgenerate
	assign rd_prio[2] = 1'b0;
	wt_dcache_wbuffer #(.ArianeCfg(ArianeCfg)) i_wt_dcache_wbuffer(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.empty_o(wbuffer_empty_o),
		.not_ni_o(wbuffer_not_ni_o),
		.cache_en_i(cache_en),
		.req_port_i(req_ports_i[(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) + (2 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)))+:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78 : 1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))]),
		.req_port_o(req_ports_o[132+:66]),
		.miss_req_o(miss_req[2]),
		.miss_ack_i(miss_ack[2]),
		.miss_we_o(miss_we[2]),
		.miss_wdata_o(miss_wdata[128+:64]),
		.miss_vld_bits_o(miss_vld_bits[16+:ariane_pkg_DCACHE_SET_ASSOC]),
		.miss_paddr_o(miss_paddr[112+:56]),
		.miss_nc_o(miss_nc[2]),
		.miss_size_o(miss_size[6+:3]),
		.miss_id_o(miss_id[4+:2]),
		.miss_rtrn_vld_i(miss_rtrn_vld[2]),
		.miss_rtrn_id_i(miss_rtrn_id),
		.rd_tag_o(rd_tag[88+:ariane_pkg_DCACHE_TAG_WIDTH]),
		.rd_idx_o(rd_idx[16+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH]),
		.rd_off_o(rd_off[8+:wt_cache_pkg_DCACHE_OFFSET_WIDTH]),
		.rd_req_o(rd_req[2]),
		.rd_tag_only_o(rd_tag_only[2]),
		.rd_ack_i(rd_ack[2]),
		.rd_data_i(rd_data),
		.rd_vld_bits_i(rd_vld_bits),
		.rd_hit_oh_i(rd_hit_oh),
		.wr_cl_vld_i(wr_cl_vld),
		.wr_cl_idx_i(wr_cl_idx),
		.wr_req_o(wr_req),
		.wr_ack_i(wr_ack),
		.wr_idx_o(wr_idx),
		.wr_off_o(wr_off),
		.wr_data_o(wr_data),
		.wr_data_be_o(wr_data_be),
		.wbuffer_data_o(wbuffer_data),
		.tx_paddr_o(tx_paddr),
		.tx_vld_o(tx_vld)
	);
	wt_dcache_mem #(
		.Axi64BitCompliant(ArianeCfg[97]),
		.NumPorts(NumPorts)
	) i_wt_dcache_mem(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rd_prio_i(rd_prio),
		.rd_tag_i(rd_tag),
		.rd_idx_i(rd_idx),
		.rd_off_i(rd_off),
		.rd_req_i(rd_req),
		.rd_tag_only_i(rd_tag_only),
		.rd_ack_o(rd_ack),
		.rd_vld_bits_o(rd_vld_bits),
		.rd_hit_oh_o(rd_hit_oh),
		.rd_data_o(rd_data),
		.wr_cl_vld_i(wr_cl_vld),
		.wr_cl_nc_i(wr_cl_nc),
		.wr_cl_we_i(wr_cl_we),
		.wr_cl_tag_i(wr_cl_tag),
		.wr_cl_idx_i(wr_cl_idx),
		.wr_cl_off_i(wr_cl_off),
		.wr_cl_data_i(wr_cl_data),
		.wr_cl_data_be_i(wr_cl_data_be),
		.wr_vld_bits_i(wr_vld_bits),
		.wr_req_i(wr_req),
		.wr_ack_o(wr_ack),
		.wr_idx_i(wr_idx),
		.wr_off_i(wr_off),
		.wr_data_i(wr_data),
		.wr_data_be_i(wr_data_be),
		.wbuffer_data_i(wbuffer_data)
	);
endmodule
module wt_dcache_missunit (
	clk_i,
	rst_ni,
	enable_i,
	flush_i,
	flush_ack_o,
	miss_o,
	wbuffer_empty_i,
	cache_en_o,
	amo_req_i,
	amo_resp_o,
	miss_req_i,
	miss_ack_o,
	miss_nc_i,
	miss_we_i,
	miss_wdata_i,
	miss_paddr_i,
	miss_vld_bits_i,
	miss_size_i,
	miss_id_i,
	miss_replay_o,
	miss_rtrn_vld_o,
	miss_rtrn_id_o,
	tx_paddr_i,
	tx_vld_i,
	wr_cl_vld_o,
	wr_cl_nc_o,
	wr_cl_we_o,
	wr_cl_tag_o,
	wr_cl_idx_o,
	wr_cl_off_o,
	wr_cl_data_o,
	wr_cl_data_be_o,
	wr_vld_bits_o,
	mem_rtrn_vld_i,
	mem_rtrn_i,
	mem_data_req_o,
	mem_data_ack_i,
	mem_data_o
);
	parameter [0:0] Axi64BitCompliant = 1'b0;
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	parameter [1:0] AmoTxId = 1;
	parameter [31:0] NumPorts = 3;
	input wire clk_i;
	input wire rst_ni;
	input wire enable_i;
	input wire flush_i;
	output reg flush_ack_o;
	output wire miss_o;
	input wire wbuffer_empty_i;
	output wire cache_en_o;
	input wire [134:0] amo_req_i;
	output reg [64:0] amo_resp_o;
	input wire [NumPorts - 1:0] miss_req_i;
	output reg [NumPorts - 1:0] miss_ack_o;
	input wire [NumPorts - 1:0] miss_nc_i;
	input wire [NumPorts - 1:0] miss_we_i;
	input wire [(NumPorts * 64) - 1:0] miss_wdata_i;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	input wire [(NumPorts * 56) - 1:0] miss_paddr_i;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	input wire [(NumPorts * ariane_pkg_DCACHE_SET_ASSOC) - 1:0] miss_vld_bits_i;
	input wire [(NumPorts * 3) - 1:0] miss_size_i;
	input wire [(NumPorts * 2) - 1:0] miss_id_i;
	output reg [NumPorts - 1:0] miss_replay_o;
	output reg [NumPorts - 1:0] miss_rtrn_vld_o;
	output wire [1:0] miss_rtrn_id_o;
	localparam wt_cache_pkg_DCACHE_MAX_TX = 4;
	input wire [223:0] tx_paddr_i;
	input wire [3:0] tx_vld_i;
	output wire wr_cl_vld_o;
	output wire wr_cl_nc_o;
	output wire [7:0] wr_cl_we_o;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	output wire [43:0] wr_cl_tag_o;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	localparam wt_cache_pkg_DCACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_DCACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_DCACHE_CL_IDX_WIDTH = 8;
	output wire [7:0] wr_cl_idx_o;
	output wire [3:0] wr_cl_off_o;
	output wire [127:0] wr_cl_data_o;
	output wire [15:0] wr_cl_data_be_o;
	output wire [7:0] wr_vld_bits_o;
	input wire mem_rtrn_vld_i;
	localparam [31:0] ariane_pkg_ICACHE_INDEX_WIDTH = 12;
	localparam wt_cache_pkg_L15_SET_ASSOC = ariane_pkg_DCACHE_SET_ASSOC;
	localparam wt_cache_pkg_L15_WAY_WIDTH = 3;
	input wire [149:0] mem_rtrn_i;
	output reg mem_data_req_o;
	input wire mem_data_ack_i;
	localparam wt_cache_pkg_L1D_WAY_WIDTH = 3;
	output reg [134:0] mem_data_o;
	reg [2:0] state_d;
	reg [2:0] state_q;
	wire [(73 + $clog2(NumPorts)) - 1:0] mshr_d;
	reg [(73 + $clog2(NumPorts)) - 1:0] mshr_q;
	wire [2:0] repl_way;
	wire [2:0] inv_way;
	wire [2:0] rnd_way;
	wire mshr_vld_d;
	reg mshr_vld_q;
	reg mshr_vld_q1;
	reg mshr_allocate;
	reg update_lfsr;
	wire all_ways_valid;
	reg enable_d;
	reg enable_q;
	reg flush_ack_d;
	reg flush_ack_q;
	reg flush_en;
	wire flush_done;
	reg mask_reads;
	reg lock_reqs;
	reg amo_sel;
	wire miss_is_write;
	wire amo_req_d;
	reg amo_req_q;
	wire [63:0] amo_data;
	wire [63:0] amo_rtrn_mux;
	wire [55:0] tmp_paddr;
	wire [$clog2(NumPorts) - 1:0] miss_port_idx;
	wire [7:0] cnt_d;
	reg [7:0] cnt_q;
	wire [NumPorts - 1:0] miss_req_masked_d;
	reg [NumPorts - 1:0] miss_req_masked_q;
	reg inv_vld;
	reg inv_vld_all;
	wire cl_write_en;
	reg load_ack;
	reg store_ack;
	reg amo_ack;
	wire [NumPorts - 1:0] mshr_rdrd_collision_d;
	reg [NumPorts - 1:0] mshr_rdrd_collision_q;
	wire [NumPorts - 1:0] mshr_rdrd_collision;
	reg tx_rdwr_collision;
	wire mshr_rdwr_collision;
	assign cache_en_o = enable_q;
	assign cnt_d = (flush_en ? cnt_q + 1 : {wt_cache_pkg_DCACHE_CL_IDX_WIDTH {1'sb0}});
	assign flush_done = cnt_q == 255;
	assign miss_req_masked_d = (lock_reqs ? miss_req_masked_q : (mask_reads ? miss_we_i & miss_req_i : miss_req_i));
	assign miss_is_write = miss_we_i[miss_port_idx];
	lzc #(.WIDTH(NumPorts)) i_lzc_reqs(
		.in_i(miss_req_masked_d),
		.cnt_o(miss_port_idx),
		.empty_o()
	);
	always @(*) begin : p_ack
		miss_ack_o = 1'sb0;
		if (!amo_sel)
			miss_ack_o[miss_port_idx] = mem_data_ack_i & mem_data_req_o;
	end
	lzc #(.WIDTH(ariane_pkg_DCACHE_SET_ASSOC)) i_lzc_inv(
		.in_i(~miss_vld_bits_i[miss_port_idx * ariane_pkg_DCACHE_SET_ASSOC+:ariane_pkg_DCACHE_SET_ASSOC]),
		.cnt_o(inv_way),
		.empty_o(all_ways_valid)
	);
	lfsr_8bit #(.WIDTH(ariane_pkg_DCACHE_SET_ASSOC)) i_lfsr_inv(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.en_i(update_lfsr),
		.refill_way_oh(),
		.refill_way_bin(rnd_way)
	);
	assign repl_way = (all_ways_valid ? rnd_way : inv_way);
	assign mshr_d[3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))-:((14 + ($clog2(NumPorts) + 2)) >= (14 + ($clog2(NumPorts) + 0)) ? ((3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))) - (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))))) + 1 : ((ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))) - (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) + 1)] = (mshr_allocate ? miss_size_i[miss_port_idx * 3+:3] : mshr_q[3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))-:((14 + ($clog2(NumPorts) + 2)) >= (14 + ($clog2(NumPorts) + 0)) ? ((3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))) - (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))))) + 1 : ((ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))) - (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) + 1)]);
	assign mshr_d[riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))-:((70 + ($clog2(NumPorts) + 2)) >= (17 + ($clog2(NumPorts) + 0)) ? ((riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))))) + 1 : ((3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))))) - (riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))))) + 1)] = (mshr_allocate ? miss_paddr_i[miss_port_idx * 56+:56] : mshr_q[riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))-:((70 + ($clog2(NumPorts) + 2)) >= (17 + ($clog2(NumPorts) + 0)) ? ((riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))))) + 1 : ((3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))))) - (riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))))) + 1)]);
	assign mshr_d[ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))-:((11 + ($clog2(NumPorts) + 2)) >= (6 + ($clog2(NumPorts) + 0)) ? ((ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))) - (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))) + 1 : ((wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))) - (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))) + 1)] = (mshr_allocate ? miss_vld_bits_i[miss_port_idx * ariane_pkg_DCACHE_SET_ASSOC+:ariane_pkg_DCACHE_SET_ASSOC] : mshr_q[ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))-:((11 + ($clog2(NumPorts) + 2)) >= (6 + ($clog2(NumPorts) + 0)) ? ((ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))) - (wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0)))) + 1 : ((wt_cache_pkg_CACHE_ID_WIDTH + (4 + ($clog2(NumPorts) + 0))) - (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))) + 1)]);
	assign mshr_d[wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))-:((3 + ($clog2(NumPorts) + 2)) >= (4 + ($clog2(NumPorts) + 0)) ? ((wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))) - (4 + ($clog2(NumPorts) + 0))) + 1 : ((4 + ($clog2(NumPorts) + 0)) - (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))) + 1)] = (mshr_allocate ? miss_id_i[miss_port_idx * 2+:2] : mshr_q[wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))-:((3 + ($clog2(NumPorts) + 2)) >= (4 + ($clog2(NumPorts) + 0)) ? ((wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))) - (4 + ($clog2(NumPorts) + 0))) + 1 : ((4 + ($clog2(NumPorts) + 0)) - (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))) + 1)]);
	assign mshr_d[1 + ($clog2(NumPorts) + 2)] = (mshr_allocate ? miss_nc_i[miss_port_idx] : mshr_q[1 + ($clog2(NumPorts) + 2)]);
	assign mshr_d[$clog2(NumPorts) + 2-:(($clog2(NumPorts) + 2) >= ($clog2(NumPorts) + 0) ? (($clog2(NumPorts) + 2) - ($clog2(NumPorts) + 0)) + 1 : (($clog2(NumPorts) + 0) - ($clog2(NumPorts) + 2)) + 1)] = (mshr_allocate ? repl_way : mshr_q[$clog2(NumPorts) + 2-:(($clog2(NumPorts) + 2) >= ($clog2(NumPorts) + 0) ? (($clog2(NumPorts) + 2) - ($clog2(NumPorts) + 0)) + 1 : (($clog2(NumPorts) + 0) - ($clog2(NumPorts) + 2)) + 1)]);
	assign mshr_d[$clog2(NumPorts) - 1-:$clog2(NumPorts)] = (mshr_allocate ? miss_port_idx : mshr_q[$clog2(NumPorts) - 1-:$clog2(NumPorts)]);
	assign mshr_vld_d = (mshr_allocate ? 1'b1 : (load_ack ? 1'b0 : mshr_vld_q));
	assign miss_o = (mshr_allocate ? ~miss_nc_i[miss_port_idx] : 1'b0);
	genvar k;
	generate
		for (k = 0; k < NumPorts; k = k + 1) begin : gen_rdrd_collision
			assign mshr_rdrd_collision[k] = (mshr_q[riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))):(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 51] == miss_paddr_i[(k * 56) + 55-:52]) && (mshr_vld_q | mshr_vld_q1);
			assign mshr_rdrd_collision_d[k] = (!miss_req_i[k] ? 1'b0 : mshr_rdrd_collision_q[k] | mshr_rdrd_collision[k]);
		end
	endgenerate
	assign mshr_rdwr_collision = (mshr_q[riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2))))):(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 51] == miss_paddr_i[((NumPorts - 1) * 56) + 55-:52]) && mshr_vld_q;
	always @(*) begin : p_tx_coll
		tx_rdwr_collision = 1'b0;
		begin : sv2v_autoblock_1
			reg signed [31:0] k;
			for (k = 0; k < wt_cache_pkg_DCACHE_MAX_TX; k = k + 1)
				tx_rdwr_collision = tx_rdwr_collision | ((miss_paddr_i[(miss_port_idx * 56) + 55-:52] == tx_paddr_i[(k * 56) + 55-:52]) && tx_vld_i[k]);
		end
	end
	assign amo_data = (amo_req_i[129-:2] == 2'b10 ? {amo_req_i[0+:32], amo_req_i[0+:32]} : amo_req_i[63-:64]);
	generate
		if (Axi64BitCompliant) begin : gen_axi_rtrn_mux
			assign amo_rtrn_mux = mem_rtrn_i[19+:64];
		end
		else begin : gen_piton_rtrn_mux
			assign amo_rtrn_mux = mem_rtrn_i[19 + (amo_req_i[67:67] * 64)+:64];
		end
	endgenerate
	wire [64:1] sv2v_tmp_EB343;
	assign sv2v_tmp_EB343 = (amo_req_i[129-:2] == 2'b10 ? {{32 {amo_rtrn_mux[(amo_req_i[66] * 32) + 31]}}, amo_rtrn_mux[amo_req_i[66] * 32+:32]} : amo_rtrn_mux);
	always @(*) amo_resp_o[63-:64] = sv2v_tmp_EB343;
	assign amo_req_d = amo_req_i[134];
	wire [2:1] sv2v_tmp_9C294;
	assign sv2v_tmp_9C294 = (amo_sel ? AmoTxId : miss_id_i[miss_port_idx * 2+:2]);
	always @(*) mem_data_o[5-:2] = sv2v_tmp_9C294;
	wire [1:1] sv2v_tmp_D3E03;
	assign sv2v_tmp_D3E03 = (amo_sel ? 1'b1 : miss_nc_i[miss_port_idx]);
	always @(*) mem_data_o[6] = sv2v_tmp_D3E03;
	wire [3:1] sv2v_tmp_1DA39;
	assign sv2v_tmp_1DA39 = (amo_sel ? {3 {1'sb0}} : repl_way);
	always @(*) mem_data_o[129-:3] = sv2v_tmp_1DA39;
	wire [64:1] sv2v_tmp_A5E70;
	assign sv2v_tmp_A5E70 = (amo_sel ? amo_data : miss_wdata_i[miss_port_idx * 64+:64]);
	always @(*) mem_data_o[70-:64] = sv2v_tmp_A5E70;
	wire [3:1] sv2v_tmp_75859;
	assign sv2v_tmp_75859 = (amo_sel ? amo_req_i[129-:2] : miss_size_i[miss_port_idx * 3+:3]);
	always @(*) mem_data_o[132-:3] = sv2v_tmp_75859;
	wire [4:1] sv2v_tmp_1AA7A;
	assign sv2v_tmp_1AA7A = (amo_sel ? amo_req_i[133-:4] : 4'b0000);
	always @(*) mem_data_o[3-:4] = sv2v_tmp_1AA7A;
	assign tmp_paddr = (amo_sel ? amo_req_i[119:64] : miss_paddr_i[miss_port_idx * 56+:56]);
	function automatic [55:0] wt_cache_pkg_paddrSizeAlign;
		input reg [55:0] paddr;
		input reg [2:0] size;
		reg [55:0] out;
		begin
			out = paddr;
			case (size)
				3'b001: out[0:0] = 1'sb0;
				3'b010: out[1:0] = 1'sb0;
				3'b011: out[2:0] = 1'sb0;
				3'b111: out[3:0] = 1'sb0;
				default:
					;
			endcase
			wt_cache_pkg_paddrSizeAlign = out;
		end
	endfunction
	wire [56:1] sv2v_tmp_1873E;
	assign sv2v_tmp_1873E = wt_cache_pkg_paddrSizeAlign(tmp_paddr, mem_data_o[132-:3]);
	always @(*) mem_data_o[126-:56] = sv2v_tmp_1873E;
	reg sc_fail;
	reg sc_pass;
	wire sc_backoff_over;
	exp_backoff #(
		.Seed(3),
		.MaxExp(16)
	) i_exp_backoff(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.set_i(sc_fail),
		.clr_i(sc_pass),
		.is_zero_o(sc_backoff_over)
	);
	wire store_sent;
	wire [2:0] stores_inflight_d;
	reg [2:0] stores_inflight_q;
	assign store_sent = (mem_data_req_o & mem_data_ack_i) & (mem_data_o[134-:2] == 2'd0);
	assign stores_inflight_d = (store_ack && store_sent ? stores_inflight_q : (store_ack ? stores_inflight_q - 1 : (store_sent ? stores_inflight_q + 1 : stores_inflight_q)));
	always @(*) begin : p_rtrn_logic
		load_ack = 1'b0;
		store_ack = 1'b0;
		amo_ack = 1'b0;
		inv_vld = 1'b0;
		inv_vld_all = 1'b0;
		sc_fail = 1'b0;
		sc_pass = 1'b0;
		miss_rtrn_vld_o = 1'sb0;
		if (mem_rtrn_vld_i)
			case (mem_rtrn_i[149-:3])
				3'd2:
					if (mshr_vld_q) begin
						load_ack = 1'b1;
						miss_rtrn_vld_o[mshr_q[$clog2(NumPorts) - 1-:$clog2(NumPorts)]] = 1'b1;
					end
				3'd1:
					if (stores_inflight_q) begin
						store_ack = 1'b1;
						miss_rtrn_vld_o[NumPorts - 1] = 1'b1;
					end
				3'd3:
					if (amo_req_q) begin
						amo_ack = 1'b1;
						if (amo_req_i[133-:4] == 4'b0010) begin
							if (amo_resp_o[63-:64])
								sc_fail = 1'b1;
							else
								sc_pass = 1'b1;
						end
					end
				3'd0: begin
					inv_vld = mem_rtrn_i[18] | mem_rtrn_i[17];
					inv_vld_all = mem_rtrn_i[17];
				end
				default:
					;
			endcase
	end
	assign miss_rtrn_id_o = mem_rtrn_i[1-:wt_cache_pkg_CACHE_ID_WIDTH];
	assign wr_cl_nc_o = mshr_q[1 + ($clog2(NumPorts) + 2)];
	assign wr_cl_vld_o = load_ack | |wr_cl_we_o;
	function automatic [7:0] wt_cache_pkg_dcache_way_bin2oh;
		input reg [2:0] in;
		reg [7:0] out;
		begin
			out = 1'sb0;
			out[in] = 1'b1;
			wt_cache_pkg_dcache_way_bin2oh = out;
		end
	endfunction
	assign wr_cl_we_o = (flush_en ? {8 {1'sb1}} : (inv_vld_all ? {8 {1'sb1}} : (inv_vld ? wt_cache_pkg_dcache_way_bin2oh(mem_rtrn_i[4-:wt_cache_pkg_L15_WAY_WIDTH]) : (cl_write_en ? wt_cache_pkg_dcache_way_bin2oh(mshr_q[$clog2(NumPorts) + 2-:(($clog2(NumPorts) + 2) >= ($clog2(NumPorts) + 0) ? (($clog2(NumPorts) + 2) - ($clog2(NumPorts) + 0)) + 1 : (($clog2(NumPorts) + 0) - ($clog2(NumPorts) + 2)) + 1)]) : {8 {1'sb0}}))));
	assign wr_vld_bits_o = (flush_en ? {8 {1'sb0}} : (inv_vld ? {8 {1'sb0}} : (cl_write_en ? wt_cache_pkg_dcache_way_bin2oh(mshr_q[$clog2(NumPorts) + 2-:(($clog2(NumPorts) + 2) >= ($clog2(NumPorts) + 0) ? (($clog2(NumPorts) + 2) - ($clog2(NumPorts) + 0)) + 1 : (($clog2(NumPorts) + 0) - ($clog2(NumPorts) + 2)) + 1)]) : {8 {1'sb0}})));
	assign wr_cl_idx_o = (flush_en ? cnt_q : (inv_vld ? mem_rtrn_i[16:9] : mshr_q[(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 44:(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 51]));
	assign wr_cl_tag_o = mshr_q[(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - (56 - (ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_INDEX_WIDTH)):(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 43];
	assign wr_cl_off_o = mshr_q[(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 52:(riscv_PLEN + (3 + (ariane_pkg_DCACHE_SET_ASSOC + (wt_cache_pkg_CACHE_ID_WIDTH + (1 + ($clog2(NumPorts) + 2)))))) - 55];
	assign wr_cl_data_o = mem_rtrn_i[146-:128];
	assign wr_cl_data_be_o = (cl_write_en ? {16 {1'sb1}} : {16 {1'sb0}});
	assign cl_write_en = load_ack & ~mshr_q[1 + ($clog2(NumPorts) + 2)];
	always @(*) begin : p_fsm
		state_d = state_q;
		flush_ack_o = 1'b0;
		mem_data_o[134-:2] = 2'd1;
		mem_data_req_o = 1'b0;
		amo_resp_o[64] = 1'b0;
		miss_replay_o = 1'sb0;
		enable_d = enable_q & enable_i;
		flush_ack_d = flush_ack_q;
		flush_en = 1'b0;
		amo_sel = 1'b0;
		update_lfsr = 1'b0;
		mshr_allocate = 1'b0;
		lock_reqs = 1'b0;
		mask_reads = mshr_vld_q;
		case (state_q)
			3'd0:
				if (flush_i || (enable_i && !enable_q)) begin
					if (wbuffer_empty_i && !mshr_vld_q) begin
						flush_ack_d = flush_i;
						state_d = 3'd3;
					end
					else
						state_d = 3'd1;
				end
				else if (amo_req_i[134]) begin
					if (wbuffer_empty_i && !mshr_vld_q)
						state_d = 3'd2;
					else
						state_d = 3'd1;
				end
				else if (|miss_req_masked_d) begin
					if (miss_is_write) begin
						if (!mshr_rdwr_collision) begin
							mem_data_req_o = 1'b1;
							mem_data_o[134-:2] = 2'd0;
							if (!mem_data_ack_i)
								state_d = 3'd4;
						end
					end
					else if (!mshr_vld_q || load_ack) begin
						if (mshr_rdrd_collision_d[miss_port_idx])
							miss_replay_o[miss_port_idx] = 1'b1;
						else if (!tx_rdwr_collision) begin
							mem_data_req_o = 1'b1;
							mem_data_o[134-:2] = 2'd1;
							update_lfsr = all_ways_valid & mem_data_ack_i;
							mshr_allocate = mem_data_ack_i;
							if (!mem_data_ack_i)
								state_d = 3'd5;
						end
					end
				end
			3'd4: begin
				lock_reqs = 1'b1;
				mem_data_req_o = 1'b1;
				mem_data_o[134-:2] = 2'd0;
				if (mem_data_ack_i)
					state_d = 3'd0;
			end
			3'd5: begin
				lock_reqs = 1'b1;
				mem_data_req_o = 1'b1;
				mem_data_o[134-:2] = 2'd1;
				if (mem_data_ack_i) begin
					update_lfsr = all_ways_valid;
					mshr_allocate = 1'b1;
					state_d = 3'd0;
				end
			end
			3'd1: begin
				mask_reads = 1'b1;
				if (|miss_req_masked_d && !mshr_rdwr_collision) begin
					mem_data_req_o = 1'b1;
					mem_data_o[134-:2] = 2'd0;
				end
				if (wbuffer_empty_i && !mshr_vld_q)
					state_d = 3'd0;
			end
			3'd3: begin
				flush_en = 1'b1;
				if (flush_done) begin
					state_d = 3'd0;
					flush_ack_o = flush_ack_q;
					flush_ack_d = 1'b0;
					enable_d = enable_i;
				end
			end
			3'd2: begin
				mem_data_o[134-:2] = 2'd2;
				amo_sel = 1'b1;
				if ((amo_req_i[133-:4] != 4'b0001) || sc_backoff_over) begin
					mem_data_req_o = 1'b1;
					if (mem_data_ack_i)
						state_d = 3'd6;
				end
			end
			3'd6: begin
				amo_sel = 1'b1;
				if (amo_ack) begin
					amo_resp_o[64] = 1'b1;
					state_d = 3'd0;
				end
			end
			default: state_d = 3'd0;
		endcase
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			state_q <= 3'd3;
			cnt_q <= 1'sb0;
			enable_q <= 1'sb0;
			flush_ack_q <= 1'sb0;
			mshr_vld_q <= 1'sb0;
			mshr_vld_q1 <= 1'sb0;
			mshr_q <= 1'sb0;
			mshr_rdrd_collision_q <= 1'sb0;
			miss_req_masked_q <= 1'sb0;
			amo_req_q <= 1'sb0;
			stores_inflight_q <= 1'sb0;
		end
		else begin
			state_q <= state_d;
			cnt_q <= cnt_d;
			enable_q <= enable_d;
			flush_ack_q <= flush_ack_d;
			mshr_vld_q <= mshr_vld_d;
			mshr_vld_q1 <= mshr_vld_q;
			mshr_q <= mshr_d;
			mshr_rdrd_collision_q <= mshr_rdrd_collision_d;
			miss_req_masked_q <= miss_req_masked_d;
			amo_req_q <= amo_req_d;
			stores_inflight_q <= stores_inflight_d;
		end
	end
endmodule
module wt_dcache_mem (
	clk_i,
	rst_ni,
	rd_tag_i,
	rd_idx_i,
	rd_off_i,
	rd_req_i,
	rd_tag_only_i,
	rd_prio_i,
	rd_ack_o,
	rd_vld_bits_o,
	rd_hit_oh_o,
	rd_data_o,
	wr_cl_vld_i,
	wr_cl_nc_i,
	wr_cl_we_i,
	wr_cl_tag_i,
	wr_cl_idx_i,
	wr_cl_off_i,
	wr_cl_data_i,
	wr_cl_data_be_i,
	wr_vld_bits_i,
	wr_req_i,
	wr_ack_o,
	wr_idx_i,
	wr_off_i,
	wr_data_i,
	wr_data_be_i,
	wbuffer_data_i
);
	parameter [0:0] Axi64BitCompliant = 1'b0;
	parameter [31:0] NumPorts = 3;
	input wire clk_i;
	input wire rst_ni;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	input wire [(NumPorts * ariane_pkg_DCACHE_TAG_WIDTH) - 1:0] rd_tag_i;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	localparam wt_cache_pkg_DCACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_DCACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_DCACHE_CL_IDX_WIDTH = 8;
	input wire [(NumPorts * wt_cache_pkg_DCACHE_CL_IDX_WIDTH) - 1:0] rd_idx_i;
	input wire [(NumPorts * wt_cache_pkg_DCACHE_OFFSET_WIDTH) - 1:0] rd_off_i;
	input wire [NumPorts - 1:0] rd_req_i;
	input wire [NumPorts - 1:0] rd_tag_only_i;
	input wire [NumPorts - 1:0] rd_prio_i;
	output wire [NumPorts - 1:0] rd_ack_o;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	output wire [7:0] rd_vld_bits_o;
	output wire [7:0] rd_hit_oh_o;
	output wire [63:0] rd_data_o;
	input wire wr_cl_vld_i;
	input wire wr_cl_nc_i;
	input wire [7:0] wr_cl_we_i;
	input wire [43:0] wr_cl_tag_i;
	input wire [7:0] wr_cl_idx_i;
	input wire [3:0] wr_cl_off_i;
	input wire [127:0] wr_cl_data_i;
	input wire [15:0] wr_cl_data_be_i;
	input wire [7:0] wr_vld_bits_i;
	input wire [7:0] wr_req_i;
	output reg wr_ack_o;
	input wire [7:0] wr_idx_i;
	input wire [3:0] wr_off_i;
	input wire [63:0] wr_data_i;
	input wire [7:0] wr_data_be_i;
	localparam wt_cache_pkg_DCACHE_WBUF_DEPTH = 8;
	input wire [(8 * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] wbuffer_data_i;
	localparam wt_cache_pkg_DCACHE_NUM_BANKS = 2;
	reg [1:0] bank_req;
	reg [1:0] bank_we;
	wire [127:0] bank_be;
	reg [15:0] bank_idx;
	wire [7:0] bank_idx_d;
	reg [7:0] bank_idx_q;
	wire [3:0] bank_off_d;
	reg [3:0] bank_off_q;
	wire [1023:0] bank_wdata;
	wire [1023:0] bank_rdata;
	wire [511:0] rdata_cl;
	wire [43:0] rd_tag;
	wire [7:0] vld_req;
	reg vld_we;
	wire [7:0] vld_wdata;
	wire [(ariane_pkg_DCACHE_SET_ASSOC * ariane_pkg_DCACHE_TAG_WIDTH) - 1:0] tag_rdata;
	wire [7:0] vld_addr;
	wire [$clog2(NumPorts) - 1:0] vld_sel_d;
	reg [$clog2(NumPorts) - 1:0] vld_sel_q;
	wire [7:0] wbuffer_hit_oh;
	wire [7:0] wbuffer_be;
	wire [63:0] wbuffer_rdata;
	wire [63:0] rdata;
	wire [63:0] wbuffer_cmp_addr;
	wire cmp_en_d;
	reg cmp_en_q;
	wire rd_acked;
	reg [NumPorts - 1:0] bank_collision;
	wire [NumPorts - 1:0] rd_req_masked;
	wire [NumPorts - 1:0] rd_req_prio;
	genvar k;
	generate
		for (k = 0; k < wt_cache_pkg_DCACHE_NUM_BANKS; k = k + 1) begin : gen_bank
			genvar j;
			for (j = 0; j < ariane_pkg_DCACHE_SET_ASSOC; j = j + 1) begin : gen_bank_way
				assign bank_be[((k * ariane_pkg_DCACHE_SET_ASSOC) + j) * 8+:8] = (wr_cl_we_i[j] & wr_cl_vld_i ? wr_cl_data_be_i[k * 8+:8] : (wr_req_i[j] & wr_ack_o ? wr_data_be_i : {8 {1'sb0}}));
				assign bank_wdata[((k * ariane_pkg_DCACHE_SET_ASSOC) + j) * 64+:64] = (wr_cl_we_i[j] & wr_cl_vld_i ? wr_cl_data_i[k * 64+:64] : wr_data_i);
			end
		end
	endgenerate
	assign vld_wdata = wr_vld_bits_i;
	assign vld_addr = (wr_cl_vld_i ? wr_cl_idx_i : rd_idx_i[vld_sel_d * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH]);
	assign rd_tag = rd_tag_i[vld_sel_q * ariane_pkg_DCACHE_TAG_WIDTH+:ariane_pkg_DCACHE_TAG_WIDTH];
	assign bank_off_d = (wr_cl_vld_i ? wr_cl_off_i : rd_off_i[vld_sel_d * wt_cache_pkg_DCACHE_OFFSET_WIDTH+:wt_cache_pkg_DCACHE_OFFSET_WIDTH]);
	assign bank_idx_d = (wr_cl_vld_i ? wr_cl_idx_i : rd_idx_i[vld_sel_d * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH]);
	assign vld_req = (wr_cl_vld_i ? wr_cl_we_i : (rd_acked ? {8 {1'sb1}} : {8 {1'sb0}}));
	assign rd_req_prio = rd_req_i & rd_prio_i;
	assign rd_req_masked = (|rd_req_prio ? rd_req_prio : rd_req_i);
	wire rd_req;
	localparam [0:0] sv2v_uu_i_rr_arb_tree_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_NumIn = NumPorts;
	localparam [$clog2(sv2v_uu_i_rr_arb_tree_NumIn) - 1:0] sv2v_uu_i_rr_arb_tree_ext_rr_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_DataWidth = 1;
	localparam [(sv2v_uu_i_rr_arb_tree_NumIn * sv2v_uu_i_rr_arb_tree_DataWidth) - 1:0] sv2v_uu_i_rr_arb_tree_ext_data_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(NumPorts),
		.DataWidth(1)
	) i_rr_arb_tree(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_rr_arb_tree_ext_flush_i_0),
		.rr_i(sv2v_uu_i_rr_arb_tree_ext_rr_i_0),
		.req_i(rd_req_masked),
		.gnt_o(rd_ack_o),
		.data_i(sv2v_uu_i_rr_arb_tree_ext_data_i_0),
		.gnt_i(~wr_cl_vld_i),
		.req_o(rd_req),
		.data_o(),
		.idx_o(vld_sel_d)
	);
	assign rd_acked = rd_req & ~wr_cl_vld_i;
	localparam wt_cache_pkg_DCACHE_NUM_BANKS_WIDTH = 1;
	function automatic [1:0] wt_cache_pkg_dcache_cl_bin2oh;
		input reg [0:0] in;
		reg [1:0] out;
		begin
			out = 1'sb0;
			out[in] = 1'b1;
			wt_cache_pkg_dcache_cl_bin2oh = out;
		end
	endfunction
	function automatic [7:0] sv2v_cast_680C3;
		input reg [7:0] inp;
		sv2v_cast_680C3 = inp;
	endfunction
	always @(*) begin : p_bank_req
		vld_we = wr_cl_vld_i;
		bank_req = 1'sb0;
		wr_ack_o = 1'sb0;
		bank_we = 1'sb0;
		bank_idx = {wt_cache_pkg_DCACHE_NUM_BANKS {sv2v_cast_680C3(wr_idx_i)}};
		begin : sv2v_autoblock_1
			reg signed [31:0] k;
			for (k = 0; k < NumPorts; k = k + 1)
				bank_collision[k] = rd_off_i[(k * wt_cache_pkg_DCACHE_OFFSET_WIDTH) + 3-:1] == wr_off_i[3:3];
		end
		if (wr_cl_vld_i & |wr_cl_we_i) begin
			bank_req = 1'sb1;
			bank_we = 1'sb1;
			bank_idx = {wt_cache_pkg_DCACHE_NUM_BANKS {sv2v_cast_680C3(wr_cl_idx_i)}};
		end
		else begin
			if (rd_acked) begin
				if (!rd_tag_only_i[vld_sel_d]) begin
					bank_req = wt_cache_pkg_dcache_cl_bin2oh(rd_off_i[(vld_sel_d * wt_cache_pkg_DCACHE_OFFSET_WIDTH) + 3-:1]);
					bank_idx[rd_off_i[(vld_sel_d * wt_cache_pkg_DCACHE_OFFSET_WIDTH) + 3-:1] * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH] = rd_idx_i[vld_sel_d * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH];
				end
			end
			if (|wr_req_i) begin
				if (rd_tag_only_i[vld_sel_d] || !(rd_ack_o[vld_sel_d] && bank_collision[vld_sel_d])) begin
					wr_ack_o = 1'b1;
					bank_req = bank_req | wt_cache_pkg_dcache_cl_bin2oh(wr_off_i[3:3]);
					bank_we = wt_cache_pkg_dcache_cl_bin2oh(wr_off_i[3:3]);
				end
			end
		end
	end
	wire [3:0] wr_cl_off;
	wire [2:0] wbuffer_hit_idx;
	wire [2:0] rd_hit_idx;
	assign cmp_en_d = |vld_req & ~vld_we;
	assign wbuffer_cmp_addr = (wr_cl_vld_i ? {wr_cl_tag_i, wr_cl_idx_i, wr_cl_off_i} : {rd_tag, bank_idx_q, bank_off_q});
	genvar i;
	generate
		for (i = 0; i < ariane_pkg_DCACHE_SET_ASSOC; i = i + 1) begin : gen_tag_cmpsel
			assign rd_hit_oh_o[i] = ((rd_tag == tag_rdata[i * ariane_pkg_DCACHE_TAG_WIDTH+:ariane_pkg_DCACHE_TAG_WIDTH]) & rd_vld_bits_o[i]) & cmp_en_q;
			assign rdata_cl[i * 64+:64] = bank_rdata[((bank_off_q[3:3] * ariane_pkg_DCACHE_SET_ASSOC) + i) * 64+:64];
		end
		for (k = 0; k < wt_cache_pkg_DCACHE_WBUF_DEPTH; k = k + 1) begin : gen_wbuffer_hit
			assign wbuffer_hit_oh[k] = |wbuffer_data_i[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8] & (wbuffer_data_i[(k * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96)-:(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96) >= 97 ? ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH : 98 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 96))] == (wbuffer_cmp_addr >> 3));
		end
	endgenerate
	lzc #(.WIDTH(wt_cache_pkg_DCACHE_WBUF_DEPTH)) i_lzc_wbuffer_hit(
		.in_i(wbuffer_hit_oh),
		.cnt_o(wbuffer_hit_idx),
		.empty_o()
	);
	lzc #(.WIDTH(ariane_pkg_DCACHE_SET_ASSOC)) i_lzc_rd_hit(
		.in_i(rd_hit_oh_o),
		.cnt_o(rd_hit_idx),
		.empty_o()
	);
	assign wbuffer_rdata = wbuffer_data_i[(wbuffer_hit_idx * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 96-:64];
	assign wbuffer_be = (|wbuffer_hit_oh ? wbuffer_data_i[(wbuffer_hit_idx * (((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 89) + ariane_pkg_DCACHE_SET_ASSOC)) + 24-:8] : {8 {1'sb0}});
	generate
		if (Axi64BitCompliant) begin : gen_axi_off
			assign wr_cl_off = (wr_cl_nc_i ? {wt_cache_pkg_DCACHE_OFFSET_WIDTH {1'sb0}} : wr_cl_off_i[3:3]);
		end
		else begin : gen_piton_off
			assign wr_cl_off = wr_cl_off_i[3:3];
		end
	endgenerate
	assign rdata = (wr_cl_vld_i ? wr_cl_data_i[wr_cl_off * 64+:64] : rdata_cl[rd_hit_idx * 64+:64]);
	generate
		for (k = 0; k < 8; k = k + 1) begin : gen_rd_data
			assign rd_data_o[8 * k+:8] = (wbuffer_be[k] ? wbuffer_rdata[8 * k+:8] : rdata[8 * k+:8]);
		end
	endgenerate
	wire [ariane_pkg_DCACHE_TAG_WIDTH:0] vld_tag_rdata [7:0];
	generate
		for (k = 0; k < wt_cache_pkg_DCACHE_NUM_BANKS; k = k + 1) begin : gen_data_banks
			sram #(
				.DATA_WIDTH(512),
				.NUM_WORDS(wt_cache_pkg_DCACHE_NUM_WORDS)
			) i_data_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(bank_req[k]),
				.we_i(bank_we[k]),
				.addr_i(bank_idx[k * wt_cache_pkg_DCACHE_CL_IDX_WIDTH+:wt_cache_pkg_DCACHE_CL_IDX_WIDTH]),
				.wdata_i(bank_wdata[64 * (k * ariane_pkg_DCACHE_SET_ASSOC)+:512]),
				.be_i(bank_be[8 * (k * ariane_pkg_DCACHE_SET_ASSOC)+:64]),
				.rdata_o(bank_rdata[64 * (k * ariane_pkg_DCACHE_SET_ASSOC)+:512])
			);
		end
		for (i = 0; i < ariane_pkg_DCACHE_SET_ASSOC; i = i + 1) begin : gen_tag_srams
			assign tag_rdata[i * ariane_pkg_DCACHE_TAG_WIDTH+:ariane_pkg_DCACHE_TAG_WIDTH] = vld_tag_rdata[i][43:0];
			assign rd_vld_bits_o[i] = vld_tag_rdata[i][ariane_pkg_DCACHE_TAG_WIDTH];
			localparam sv2v_uu_i_tag_sram_DATA_WIDTH = 45;
			localparam [5:0] sv2v_uu_i_tag_sram_ext_be_i_1 = 1'sb1;
			sram #(
				.DATA_WIDTH(45),
				.NUM_WORDS(wt_cache_pkg_DCACHE_NUM_WORDS)
			) i_tag_sram(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.req_i(vld_req[i]),
				.we_i(vld_we),
				.addr_i(vld_addr),
				.wdata_i({vld_wdata[i], wr_cl_tag_i}),
				.be_i(sv2v_uu_i_tag_sram_ext_be_i_1),
				.rdata_o(vld_tag_rdata[i])
			);
		end
	endgenerate
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			bank_idx_q <= 1'sb0;
			bank_off_q <= 1'sb0;
			vld_sel_q <= 1'sb0;
			cmp_en_q <= 1'sb0;
		end
		else begin
			bank_idx_q <= bank_idx_d;
			bank_off_q <= bank_off_d;
			vld_sel_q <= vld_sel_d;
			cmp_en_q <= cmp_en_d;
		end
	end
endmodule
module wt_dcache_ctrl (
	clk_i,
	rst_ni,
	cache_en_i,
	req_port_i,
	req_port_o,
	miss_req_o,
	miss_ack_i,
	miss_we_o,
	miss_wdata_o,
	miss_vld_bits_o,
	miss_paddr_o,
	miss_nc_o,
	miss_size_o,
	miss_id_o,
	miss_replay_i,
	miss_rtrn_vld_i,
	wr_cl_vld_i,
	rd_tag_o,
	rd_idx_o,
	rd_off_o,
	rd_req_o,
	rd_tag_only_o,
	rd_ack_i,
	rd_data_i,
	rd_vld_bits_i,
	rd_hit_oh_i
);
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	parameter [1:0] RdTxId = 1;
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire cache_en_i;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	input wire [(ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77:0] req_port_i;
	output reg [65:0] req_port_o;
	output reg miss_req_o;
	input wire miss_ack_i;
	output wire miss_we_o;
	output wire [63:0] miss_wdata_o;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	output wire [7:0] miss_vld_bits_o;
	output wire [55:0] miss_paddr_o;
	output wire miss_nc_o;
	output wire [2:0] miss_size_o;
	output wire [1:0] miss_id_o;
	input wire miss_replay_i;
	input wire miss_rtrn_vld_i;
	input wire wr_cl_vld_i;
	output wire [43:0] rd_tag_o;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	localparam wt_cache_pkg_DCACHE_OFFSET_WIDTH = 4;
	localparam wt_cache_pkg_DCACHE_NUM_WORDS = 256;
	localparam wt_cache_pkg_DCACHE_CL_IDX_WIDTH = 8;
	output wire [7:0] rd_idx_o;
	output wire [3:0] rd_off_o;
	output reg rd_req_o;
	output wire rd_tag_only_o;
	input wire rd_ack_i;
	input wire [63:0] rd_data_i;
	input wire [7:0] rd_vld_bits_i;
	input wire [7:0] rd_hit_oh_i;
	reg [2:0] state_d;
	reg [2:0] state_q;
	wire [43:0] address_tag_d;
	reg [43:0] address_tag_q;
	wire [7:0] address_idx_d;
	reg [7:0] address_idx_q;
	wire [3:0] address_off_d;
	reg [3:0] address_off_q;
	wire [7:0] vld_data_d;
	reg [7:0] vld_data_q;
	reg save_tag;
	wire rd_req_d;
	reg rd_req_q;
	wire rd_ack_d;
	reg rd_ack_q;
	wire [1:0] data_size_d;
	reg [1:0] data_size_q;
	assign vld_data_d = (rd_req_q ? rd_vld_bits_i : vld_data_q);
	assign address_tag_d = (save_tag ? req_port_i[121-:44] : address_tag_q);
	assign address_idx_d = (req_port_o[65] ? req_port_i[133:126] : address_idx_q);
	assign address_off_d = (req_port_o[65] ? req_port_i[125:122] : address_off_q);
	assign data_size_d = (req_port_o[65] ? req_port_i[3-:2] : data_size_q);
	assign rd_tag_o = address_tag_d;
	assign rd_idx_o = address_idx_d;
	assign rd_off_o = address_off_d;
	wire [64:1] sv2v_tmp_2BF52;
	assign sv2v_tmp_2BF52 = rd_data_i;
	always @(*) req_port_o[63-:64] = sv2v_tmp_2BF52;
	assign miss_vld_bits_o = vld_data_q;
	assign miss_paddr_o = {address_tag_q, address_idx_q, address_off_q};
	assign miss_size_o = (miss_nc_o ? data_size_q : 3'b111);
	function automatic ariane_pkg_range_check;
		input reg [63:0] base;
		input reg [63:0] len;
		input reg [63:0] address;
		ariane_pkg_range_check = (address >= base) && (address < (base + len));
	endfunction
	function automatic ariane_pkg_is_inside_cacheable_regions;
		input reg [6433:0] Cfg;
		input reg [63:0] address;
		reg [15:0] pass;
		begin
			pass = 1'sb0;
			begin : sv2v_autoblock_1
				reg [31:0] k;
				for (k = 0; k < Cfg[2177-:32]; k = k + 1)
					pass[k] = ariane_pkg_range_check(Cfg[1122 + (k * 64)+:64], Cfg[98 + (k * 64)+:64], address);
			end
			ariane_pkg_is_inside_cacheable_regions = |pass;
		end
	endfunction
	assign miss_nc_o = ~cache_en_i | ~ariane_pkg_is_inside_cacheable_regions(ArianeCfg, {{'d20 {1'b0}}, address_tag_q, {ariane_pkg_DCACHE_INDEX_WIDTH {1'b0}}});
	assign miss_we_o = 1'sb0;
	assign miss_wdata_o = 1'sb0;
	assign miss_id_o = RdTxId;
	assign rd_req_d = rd_req_o;
	assign rd_ack_d = rd_ack_i;
	assign rd_tag_only_o = 1'sb0;
	always @(*) begin : p_fsm
		state_d = state_q;
		save_tag = 1'b0;
		rd_req_o = 1'b0;
		miss_req_o = 1'b0;
		req_port_o[64] = 1'b0;
		req_port_o[65] = 1'b0;
		case (state_q)
			3'd0:
				if (req_port_i[13]) begin
					rd_req_o = 1'b1;
					if (rd_ack_i) begin
						state_d = 3'd1;
						req_port_o[65] = 1'b1;
					end
				end
			3'd1, 3'd7: begin
				rd_req_o = 1'b1;
				if (req_port_i[1]) begin
					state_d = 3'd0;
					req_port_o[64] = 1'b1;
				end
				else if (req_port_i[0] | (state_q == 3'd7)) begin
					save_tag = state_q != 3'd7;
					if (wr_cl_vld_i || !rd_ack_q)
						state_d = 3'd6;
					else if (|rd_hit_oh_i && cache_en_i) begin
						state_d = 3'd0;
						req_port_o[64] = 1'b1;
						if (rd_ack_i && req_port_i[13]) begin
							state_d = 3'd1;
							req_port_o[65] = 1'b1;
						end
					end
					else
						state_d = 3'd2;
				end
			end
			3'd2: begin
				miss_req_o = 1'b1;
				if (req_port_i[1]) begin
					req_port_o[64] = 1'b1;
					if (miss_ack_i)
						state_d = 3'd4;
					else
						state_d = 3'd5;
				end
				else if (miss_replay_i)
					state_d = 3'd6;
				else if (miss_ack_i)
					state_d = 3'd3;
			end
			3'd3:
				if (req_port_i[1]) begin
					req_port_o[64] = 1'b1;
					if (miss_rtrn_vld_i)
						state_d = 3'd0;
					else
						state_d = 3'd4;
				end
				else if (miss_rtrn_vld_i) begin
					state_d = 3'd0;
					req_port_o[64] = 1'b1;
				end
			3'd6: begin
				rd_req_o = 1'b1;
				if (req_port_i[1]) begin
					req_port_o[64] = 1'b1;
					state_d = 3'd0;
				end
				else if (rd_ack_i)
					state_d = 3'd7;
			end
			3'd5: begin
				miss_req_o = 1'b1;
				if (miss_replay_i)
					state_d = 3'd0;
				else if (miss_ack_i)
					state_d = 3'd4;
			end
			3'd4:
				if (miss_rtrn_vld_i)
					state_d = 3'd0;
			default: state_d = 3'd0;
		endcase
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			state_q <= 3'd0;
			address_tag_q <= 1'sb0;
			address_idx_q <= 1'sb0;
			address_off_q <= 1'sb0;
			vld_data_q <= 1'sb0;
			data_size_q <= 1'sb0;
			rd_req_q <= 1'sb0;
			rd_ack_q <= 1'sb0;
		end
		else begin
			state_q <= state_d;
			address_tag_q <= address_tag_d;
			address_idx_q <= address_idx_d;
			address_off_q <= address_off_d;
			vld_data_q <= vld_data_d;
			data_size_q <= data_size_d;
			rd_req_q <= rd_req_d;
			rd_ack_q <= rd_ack_d;
		end
	end
endmodule
module wt_cache_subsystem (
	clk_i,
	rst_ni,
	icache_en_i,
	icache_flush_i,
	icache_miss_o,
	icache_areq_i,
	icache_areq_o,
	icache_dreq_i,
	icache_dreq_o,
	dcache_enable_i,
	dcache_flush_i,
	dcache_flush_ack_o,
	dcache_miss_o,
	dcache_amo_req_i,
	dcache_amo_resp_o,
	dcache_req_ports_i,
	dcache_req_ports_o,
	wbuffer_empty_o,
	wbuffer_not_ni_o,
	axi_req_o,
	axi_resp_i
);
	localparam ariane_pkg_NrMaxRules = 16;
	localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 6434'h8000000800000020000000008000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000040000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000004000000000000000040000000000400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000002000000000000000000000008;
	parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
	input wire clk_i;
	input wire rst_ni;
	input wire icache_en_i;
	input wire icache_flush_i;
	output wire icache_miss_o;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	input wire [185:0] icache_areq_i;
	localparam riscv_VLEN = 64;
	output wire [64:0] icache_areq_o;
	input wire [67:0] icache_dreq_i;
	localparam [31:0] ariane_pkg_FETCH_WIDTH = 32;
	output wire [226:0] icache_dreq_o;
	input wire dcache_enable_i;
	input wire dcache_flush_i;
	output wire dcache_flush_ack_o;
	output wire dcache_miss_o;
	input wire [134:0] dcache_amo_req_i;
	output wire [64:0] dcache_amo_resp_o;
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = 44;
	input wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? (3 * ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 78)) - 1 : (3 * (1 - ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77))) + ((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 76)):(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77) >= 0 ? 0 : (ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + 77)] dcache_req_ports_i;
	output wire [197:0] dcache_req_ports_o;
	output wire wbuffer_empty_o;
	output wire wbuffer_not_ni_o;
	localparam ariane_axi_AddrWidth = 64;
	localparam ariane_axi_IdWidth = 4;
	localparam ariane_axi_UserWidth = 1;
	localparam ariane_axi_DataWidth = 64;
	localparam ariane_axi_StrbWidth = 8;
	output wire [280:0] axi_req_o;
	input wire [83:0] axi_resp_i;
	wire icache_adapter_data_req;
	wire adapter_icache_data_ack;
	wire adapter_icache_rtrn_vld;
	localparam [31:0] ariane_pkg_ICACHE_SET_ASSOC = 4;
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	wire [60:0] icache_adapter;
	localparam [31:0] ariane_pkg_ICACHE_LINE_WIDTH = 128;
	localparam [31:0] ariane_pkg_ICACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	localparam wt_cache_pkg_L15_SET_ASSOC = ariane_pkg_DCACHE_SET_ASSOC;
	localparam wt_cache_pkg_L15_WAY_WIDTH = 3;
	wire [147:0] adapter_icache;
	wire dcache_adapter_data_req;
	wire adapter_dcache_data_ack;
	wire adapter_dcache_rtrn_vld;
	localparam wt_cache_pkg_L1D_WAY_WIDTH = 3;
	wire [134:0] dcache_adapter;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	wire [149:0] adapter_dcache;
	cva6_icache #(
		.RdTxId(0),
		.ArianeCfg(ArianeCfg)
	) i_cva6_icache(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(icache_flush_i),
		.en_i(icache_en_i),
		.miss_o(icache_miss_o),
		.areq_i(icache_areq_i),
		.areq_o(icache_areq_o),
		.dreq_i(icache_dreq_i),
		.dreq_o(icache_dreq_o),
		.mem_rtrn_vld_i(adapter_icache_rtrn_vld),
		.mem_rtrn_i(adapter_icache),
		.mem_data_req_o(icache_adapter_data_req),
		.mem_data_ack_i(adapter_icache_data_ack),
		.mem_data_o(icache_adapter)
	);
	wt_dcache #(
		.RdAmoTxId(1),
		.ArianeCfg(ArianeCfg)
	) i_wt_dcache(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.enable_i(dcache_enable_i),
		.flush_i(dcache_flush_i),
		.flush_ack_o(dcache_flush_ack_o),
		.miss_o(dcache_miss_o),
		.wbuffer_empty_o(wbuffer_empty_o),
		.wbuffer_not_ni_o(wbuffer_not_ni_o),
		.amo_req_i(dcache_amo_req_i),
		.amo_resp_o(dcache_amo_resp_o),
		.req_ports_i(dcache_req_ports_i),
		.req_ports_o(dcache_req_ports_o),
		.mem_rtrn_vld_i(adapter_dcache_rtrn_vld),
		.mem_rtrn_i(adapter_dcache),
		.mem_data_req_o(dcache_adapter_data_req),
		.mem_data_ack_i(adapter_dcache_data_ack),
		.mem_data_o(dcache_adapter)
	);
	wt_axi_adapter i_adapter(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.icache_data_req_i(icache_adapter_data_req),
		.icache_data_ack_o(adapter_icache_data_ack),
		.icache_data_i(icache_adapter),
		.icache_rtrn_vld_o(adapter_icache_rtrn_vld),
		.icache_rtrn_o(adapter_icache),
		.dcache_data_req_i(dcache_adapter_data_req),
		.dcache_data_ack_o(adapter_dcache_data_ack),
		.dcache_data_i(dcache_adapter),
		.dcache_rtrn_vld_o(adapter_dcache_rtrn_vld),
		.dcache_rtrn_o(adapter_dcache),
		.axi_req_o(axi_req_o),
		.axi_resp_i(axi_resp_i)
	);
endmodule
module wt_axi_adapter (
	clk_i,
	rst_ni,
	icache_data_req_i,
	icache_data_ack_o,
	icache_data_i,
	icache_rtrn_vld_o,
	icache_rtrn_o,
	dcache_data_req_i,
	dcache_data_ack_o,
	dcache_data_i,
	dcache_rtrn_vld_o,
	dcache_rtrn_o,
	axi_req_o,
	axi_resp_i
);
	parameter [31:0] ReqFifoDepth = 2;
	localparam wt_cache_pkg_L15_TID_WIDTH = 2;
	localparam wt_cache_pkg_DCACHE_MAX_TX = 4;
	parameter [31:0] MetaFifoDepth = wt_cache_pkg_DCACHE_MAX_TX;
	input wire clk_i;
	input wire rst_ni;
	input wire icache_data_req_i;
	output wire icache_data_ack_o;
	localparam [31:0] ariane_pkg_ICACHE_SET_ASSOC = 4;
	localparam riscv_XLEN = 64;
	localparam riscv_PLEN = 56;
	localparam wt_cache_pkg_CACHE_ID_WIDTH = wt_cache_pkg_L15_TID_WIDTH;
	input wire [60:0] icache_data_i;
	output reg icache_rtrn_vld_o;
	localparam [31:0] ariane_pkg_ICACHE_LINE_WIDTH = 128;
	localparam [31:0] ariane_pkg_ICACHE_INDEX_WIDTH = 12;
	localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
	localparam wt_cache_pkg_L15_SET_ASSOC = ariane_pkg_DCACHE_SET_ASSOC;
	localparam wt_cache_pkg_L15_WAY_WIDTH = 3;
	output reg [147:0] icache_rtrn_o;
	input wire dcache_data_req_i;
	output wire dcache_data_ack_o;
	localparam wt_cache_pkg_L1D_WAY_WIDTH = 3;
	input wire [134:0] dcache_data_i;
	output reg dcache_rtrn_vld_o;
	localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
	output reg [149:0] dcache_rtrn_o;
	localparam ariane_axi_AddrWidth = 64;
	localparam ariane_axi_IdWidth = 4;
	localparam ariane_axi_UserWidth = 1;
	localparam ariane_axi_DataWidth = 64;
	localparam ariane_axi_StrbWidth = 8;
	output wire [280:0] axi_req_o;
	input wire [83:0] axi_resp_i;
	localparam AxiNumWords = (2 * 1'd0) + (2 * 1'd1);
	wire [60:0] icache_data;
	wire icache_data_full;
	wire icache_data_empty;
	wire [134:0] dcache_data;
	wire dcache_data_full;
	wire dcache_data_empty;
	wire [1:0] arb_req;
	wire [1:0] arb_ack;
	wire arb_idx;
	wire arb_gnt;
	reg axi_rd_req;
	wire axi_rd_gnt;
	reg axi_wr_req;
	wire axi_wr_gnt;
	wire axi_wr_valid;
	wire axi_rd_valid;
	reg axi_rd_rdy;
	wire axi_wr_rdy;
	reg axi_rd_lock;
	reg axi_wr_lock;
	wire axi_rd_exokay;
	wire axi_wr_exokay;
	wire wr_exokay;
	reg [63:0] axi_rd_addr;
	reg [63:0] axi_wr_addr;
	reg [$clog2(AxiNumWords) - 1:0] axi_rd_blen;
	reg [$clog2(AxiNumWords) - 1:0] axi_wr_blen;
	reg [1:0] axi_rd_size;
	reg [1:0] axi_wr_size;
	reg [3:0] axi_rd_id_in;
	reg [3:0] axi_wr_id_in;
	wire [3:0] axi_rd_id_out;
	wire [3:0] axi_wr_id_out;
	wire [3:0] wr_id_out;
	reg [(AxiNumWords * 64) - 1:0] axi_wr_data;
	wire [63:0] axi_rd_data;
	reg [(AxiNumWords * 8) - 1:0] axi_wr_be;
	reg [5:0] axi_wr_atop;
	reg invalidate;
	reg [2:0] amo_off_d;
	reg [2:0] amo_off_q;
	reg amo_gen_r_d;
	reg amo_gen_r_q;
	wire [1:0] icache_rtrn_tid_d;
	reg [1:0] icache_rtrn_tid_q;
	wire [1:0] dcache_rtrn_tid_d;
	reg [1:0] dcache_rtrn_tid_q;
	wire [1:0] dcache_rtrn_rd_tid;
	wire [1:0] dcache_rtrn_wr_tid;
	reg dcache_rd_pop;
	reg dcache_wr_pop;
	wire icache_rd_full;
	wire icache_rd_empty;
	wire dcache_rd_full;
	wire dcache_rd_empty;
	wire dcache_wr_full;
	wire dcache_wr_empty;
	assign icache_data_ack_o = icache_data_req_i & ~icache_data_full;
	assign dcache_data_ack_o = dcache_data_req_i & ~dcache_data_full;
	assign arb_req = {~((dcache_data_empty | dcache_wr_full) | dcache_rd_full), ~(icache_data_empty | icache_rd_full)};
	assign arb_gnt = axi_rd_gnt | axi_wr_gnt;
	localparam [0:0] sv2v_uu_i_rr_arb_tree_ext_flush_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_NumIn = 2;
	localparam [0:0] sv2v_uu_i_rr_arb_tree_ext_rr_i_0 = 1'sb0;
	localparam [31:0] sv2v_uu_i_rr_arb_tree_DataWidth = 1;
	localparam [(sv2v_uu_i_rr_arb_tree_NumIn * sv2v_uu_i_rr_arb_tree_DataWidth) - 1:0] sv2v_uu_i_rr_arb_tree_ext_data_i_0 = 1'sb0;
	rr_arb_tree #(
		.NumIn(2),
		.DataWidth(1),
		.AxiVldRdy(1'b1),
		.LockIn(1'b1)
	) i_rr_arb_tree(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(sv2v_uu_i_rr_arb_tree_ext_flush_i_0),
		.rr_i(sv2v_uu_i_rr_arb_tree_ext_rr_i_0),
		.req_i(arb_req),
		.gnt_o(arb_ack),
		.data_i(sv2v_uu_i_rr_arb_tree_ext_data_i_0),
		.gnt_i(arb_gnt),
		.req_o(),
		.data_o(),
		.idx_o(arb_idx)
	);
	localparam axi_pkg_ATOP_ADD = 3'b000;
	localparam axi_pkg_ATOP_ATOMICLOAD = 2'b10;
	localparam axi_pkg_ATOP_ATOMICSWAP = 6'b110000;
	localparam axi_pkg_ATOP_CLR = 3'b001;
	localparam axi_pkg_ATOP_EOR = 3'b010;
	localparam axi_pkg_ATOP_LITTLE_END = 1'b0;
	localparam axi_pkg_ATOP_SET = 3'b011;
	localparam axi_pkg_ATOP_SMAX = 3'b100;
	localparam axi_pkg_ATOP_SMIN = 3'b101;
	localparam axi_pkg_ATOP_UMAX = 3'b110;
	localparam axi_pkg_ATOP_UMIN = 3'b111;
	function automatic [7:0] wt_cache_pkg_toByteEnable8;
		input reg [2:0] offset;
		input reg [1:0] size;
		reg [7:0] be;
		begin
			be = 1'sb0;
			case (size)
				2'b00: be[offset] = 1'sb1;
				2'b01: be[offset+:2] = 1'sb1;
				2'b10: be[offset+:4] = 1'sb1;
				default: be = 1'sb1;
			endcase
			wt_cache_pkg_toByteEnable8 = be;
		end
	endfunction
	always @(*) begin : p_axi_req
		axi_wr_id_in = arb_idx;
		axi_wr_data = dcache_data[70-:64];
		axi_wr_addr = {{8 {1'b0}}, dcache_data[126-:56]};
		axi_wr_size = dcache_data[131:130];
		axi_wr_req = 1'b0;
		axi_wr_blen = 1'sb0;
		axi_wr_be = 1'sb0;
		axi_wr_lock = 1'sb0;
		axi_wr_atop = 1'sb0;
		amo_off_d = 1'sb0;
		amo_gen_r_d = amo_gen_r_q;
		axi_rd_id_in = arb_idx;
		axi_rd_req = 1'b0;
		axi_rd_lock = 1'sb0;
		axi_rd_blen = 1'sb0;
		if (arb_idx) begin
			axi_rd_addr = {{8 {1'b0}}, dcache_data[126-:56]};
			axi_rd_size = dcache_data[131:130];
			if (dcache_data[132])
				axi_rd_blen = 1;
		end
		else begin
			axi_rd_addr = {{8 {1'b0}}, icache_data[58-:56]};
			axi_rd_size = 2'b11;
			if (!icache_data[2])
				axi_rd_blen = 1;
		end
		invalidate = 1'b0;
		if (|arb_req) begin
			if (arb_idx == 0)
				axi_rd_req = 1'b1;
			else
				case (dcache_data[134-:2])
					2'd1: axi_rd_req = 1'b1;
					2'd0: begin
						axi_wr_req = 1'b1;
						axi_wr_be = wt_cache_pkg_toByteEnable8(dcache_data[73:71], dcache_data[131:130]);
					end
					2'd2: begin
						invalidate = arb_gnt;
						axi_wr_req = 1'b1;
						axi_wr_be = wt_cache_pkg_toByteEnable8(dcache_data[73:71], dcache_data[131:130]);
						amo_gen_r_d = 1'b1;
						axi_wr_id_in[1] = 1'b1;
						case (dcache_data[3-:4])
							4'b0001: begin
								axi_rd_lock = 1'b1;
								axi_rd_req = 1'b1;
								axi_rd_id_in[1] = 1'b1;
								axi_wr_req = 1'b0;
								axi_wr_be = 1'sb0;
							end
							4'b0010: begin
								axi_wr_lock = 1'b1;
								amo_gen_r_d = 1'b0;
								case (dcache_data[131:130])
									2'b00: amo_off_d = dcache_data[73:71];
									2'b01: amo_off_d = {dcache_data[73:72], 1'b0};
									2'b10: amo_off_d = {dcache_data[73], 2'b00};
									2'b11: amo_off_d = 1'sb0;
								endcase
							end
							4'b0011: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_ATOMICSWAP};
							4'b0100: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_ADD};
							4'b0101: begin
								axi_wr_data = ~dcache_data[70-:64];
								axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_CLR};
							end
							4'b0110: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SET};
							4'b0111: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_EOR};
							4'b1000: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SMAX};
							4'b1001: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_UMAX};
							4'b1010: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_SMIN};
							4'b1011: axi_wr_atop = {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END, axi_pkg_ATOP_UMIN};
						endcase
					end
				endcase
		end
	end
	localparam signed [31:0] i_icache_data_fifo_sv2v_pfunc_651B1 = 2;
	fifo_v3_6C4C9_25B33 #(
		.dtype_i_icache_data_fifo_sv2v_pfunc_651B1(i_icache_data_fifo_sv2v_pfunc_651B1),
		.dtype_riscv_PLEN(riscv_PLEN),
		.dtype_wt_cache_pkg_CACHE_ID_WIDTH(wt_cache_pkg_CACHE_ID_WIDTH),
		.DEPTH(ReqFifoDepth)
	) i_icache_data_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(icache_data_full),
		.empty_o(icache_data_empty),
		.usage_o(),
		.data_i(icache_data_i),
		.push_i(icache_data_ack_o),
		.data_o(icache_data),
		.pop_i(arb_ack[0])
	);
	fifo_v3_77734_A8EA3 #(
		.dtype_riscv_PLEN(riscv_PLEN),
		.dtype_wt_cache_pkg_CACHE_ID_WIDTH(wt_cache_pkg_CACHE_ID_WIDTH),
		.dtype_wt_cache_pkg_L1D_WAY_WIDTH(wt_cache_pkg_L1D_WAY_WIDTH),
		.DEPTH(ReqFifoDepth)
	) i_dcache_data_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(dcache_data_full),
		.empty_o(dcache_data_empty),
		.usage_o(),
		.data_i(dcache_data_i),
		.push_i(dcache_data_ack_o),
		.data_o(dcache_data),
		.pop_i(arb_ack[1])
	);
	reg icache_rtrn_rd_en;
	reg dcache_rtrn_rd_en;
	reg icache_rtrn_vld_d;
	reg icache_rtrn_vld_q;
	reg dcache_rtrn_vld_d;
	reg dcache_rtrn_vld_q;
	fifo_v3 #(
		.DATA_WIDTH(wt_cache_pkg_CACHE_ID_WIDTH),
		.DEPTH(MetaFifoDepth)
	) i_rd_icache_id(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(icache_rd_full),
		.empty_o(icache_rd_empty),
		.usage_o(),
		.data_i(icache_data[1-:wt_cache_pkg_CACHE_ID_WIDTH]),
		.push_i(arb_ack[0] & axi_rd_gnt),
		.data_o(icache_rtrn_tid_d),
		.pop_i(icache_rtrn_vld_d)
	);
	fifo_v3 #(
		.DATA_WIDTH(wt_cache_pkg_CACHE_ID_WIDTH),
		.DEPTH(MetaFifoDepth)
	) i_rd_dcache_id(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(dcache_rd_full),
		.empty_o(dcache_rd_empty),
		.usage_o(),
		.data_i(dcache_data[5-:2]),
		.push_i(arb_ack[1] & axi_rd_gnt),
		.data_o(dcache_rtrn_rd_tid),
		.pop_i(dcache_rd_pop)
	);
	fifo_v3 #(
		.DATA_WIDTH(wt_cache_pkg_CACHE_ID_WIDTH),
		.DEPTH(MetaFifoDepth)
	) i_wr_dcache_id(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(dcache_wr_full),
		.empty_o(dcache_wr_empty),
		.usage_o(),
		.data_i(dcache_data[5-:2]),
		.push_i(arb_ack[1] & axi_wr_gnt),
		.data_o(dcache_rtrn_wr_tid),
		.pop_i(dcache_wr_pop)
	);
	assign dcache_rtrn_tid_d = (dcache_wr_pop ? dcache_rtrn_wr_tid : dcache_rtrn_rd_tid);
	wire b_full;
	wire b_empty;
	wire b_push;
	reg b_pop;
	assign axi_wr_rdy = ~b_full;
	assign b_push = axi_wr_valid & axi_wr_rdy;
	fifo_v3 #(
		.DATA_WIDTH(5),
		.DEPTH(MetaFifoDepth),
		.FALL_THROUGH(1'b1)
	) i_b_fifo(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.testmode_i(1'b0),
		.full_o(b_full),
		.empty_o(b_empty),
		.usage_o(),
		.data_i({axi_wr_exokay, axi_wr_id_out}),
		.push_i(b_push),
		.data_o({wr_exokay, wr_id_out}),
		.pop_i(b_pop)
	);
	reg icache_first_d;
	reg icache_first_q;
	reg dcache_first_d;
	reg dcache_first_q;
	reg [127:0] icache_rd_shift_d;
	reg [127:0] icache_rd_shift_q;
	reg [127:0] dcache_rd_shift_d;
	reg [127:0] dcache_rd_shift_q;
	reg [2:0] dcache_rtrn_type_d;
	reg [2:0] dcache_rtrn_type_q;
	reg [16:0] dcache_rtrn_inv_d;
	reg [16:0] dcache_rtrn_inv_q;
	reg dcache_sc_rtrn;
	wire axi_rd_last;
	always @(*) begin : p_axi_rtrn_shift
		icache_rtrn_o = 1'sb0;
		icache_rtrn_o[147] = 1'd1;
		icache_rtrn_o[1-:wt_cache_pkg_CACHE_ID_WIDTH] = icache_rtrn_tid_q;
		icache_rtrn_o[146-:128] = icache_rd_shift_q;
		icache_rtrn_vld_o = icache_rtrn_vld_q;
		dcache_rtrn_o = 1'sb0;
		dcache_rtrn_o[149-:3] = dcache_rtrn_type_q;
		dcache_rtrn_o[18-:17] = dcache_rtrn_inv_q;
		dcache_rtrn_o[1-:wt_cache_pkg_CACHE_ID_WIDTH] = dcache_rtrn_tid_q;
		dcache_rtrn_o[146-:128] = dcache_rd_shift_q;
		dcache_rtrn_vld_o = dcache_rtrn_vld_q;
		icache_rd_shift_d = icache_rd_shift_q;
		dcache_rd_shift_d = dcache_rd_shift_q;
		icache_first_d = icache_first_q;
		dcache_first_d = dcache_first_q;
		if (icache_rtrn_rd_en) begin
			icache_first_d = axi_rd_last;
			icache_rd_shift_d = {axi_rd_data, icache_rd_shift_q[64+:64]};
			if (icache_first_q)
				icache_rd_shift_d[0+:64] = axi_rd_data;
		end
		if (dcache_rtrn_rd_en) begin
			dcache_first_d = axi_rd_last;
			dcache_rd_shift_d = {axi_rd_data, dcache_rd_shift_q[64+:64]};
			if (dcache_first_q)
				dcache_rd_shift_d[0+:64] = axi_rd_data;
		end
		else if (dcache_sc_rtrn) begin
			dcache_rd_shift_d[0+:64] = 1'sb0;
			dcache_rd_shift_d[0 + (amo_off_q * 8)] = (wr_exokay ? 1'b0 : 1'b1);
		end
	end
	localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = 12;
	always @(*) begin : p_axi_rtrn_decode
		axi_rd_rdy = ~invalidate;
		icache_rtrn_rd_en = 1'b0;
		icache_rtrn_vld_d = 1'b0;
		if ((axi_rd_valid && (axi_rd_id_out == 0)) && axi_rd_rdy) begin
			icache_rtrn_rd_en = 1'b1;
			icache_rtrn_vld_d = axi_rd_last;
		end
		dcache_rtrn_rd_en = 1'b0;
		dcache_rtrn_vld_d = 1'b0;
		dcache_rd_pop = 1'b0;
		dcache_wr_pop = 1'b0;
		dcache_rtrn_inv_d = 1'sb0;
		dcache_rtrn_type_d = 3'd2;
		b_pop = 1'b0;
		dcache_sc_rtrn = 1'b0;
		if (invalidate) begin
			dcache_rtrn_type_d = 3'd0;
			dcache_rtrn_vld_d = 1'b1;
			dcache_rtrn_inv_d[15] = 1'b1;
			dcache_rtrn_inv_d[14-:12] = dcache_data[82:71];
		end
		else if ((axi_rd_valid && axi_rd_id_out[0]) && axi_rd_rdy) begin
			dcache_rtrn_rd_en = 1'b1;
			dcache_rtrn_vld_d = axi_rd_last;
			if (axi_rd_id_out[1]) begin
				dcache_rtrn_type_d = 3'd3;
				if (!dcache_wr_empty)
					dcache_wr_pop = axi_rd_last;
				else
					dcache_rd_pop = axi_rd_last;
			end
			else
				dcache_rd_pop = axi_rd_last;
		end
		else if (!b_empty) begin
			b_pop = 1'b1;
			if (wr_id_out[1]) begin
				dcache_rtrn_type_d = 3'd3;
				if (!amo_gen_r_q) begin
					dcache_rtrn_vld_d = 1'b1;
					dcache_wr_pop = 1'b1;
					dcache_sc_rtrn = 1'b1;
				end
			end
			else begin
				dcache_rtrn_type_d = 3'd1;
				dcache_rtrn_vld_d = 1'b1;
				dcache_wr_pop = 1'b1;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : p_rd_buf
		if (!rst_ni) begin
			icache_first_q <= 1'b1;
			dcache_first_q <= 1'b1;
			icache_rd_shift_q <= 1'sb0;
			dcache_rd_shift_q <= 1'sb0;
			icache_rtrn_vld_q <= 1'sb0;
			dcache_rtrn_vld_q <= 1'sb0;
			icache_rtrn_tid_q <= 1'sb0;
			dcache_rtrn_tid_q <= 1'sb0;
			dcache_rtrn_type_q <= 3'd2;
			dcache_rtrn_inv_q <= 1'sb0;
			amo_off_q <= 1'sb0;
			amo_gen_r_q <= 1'b0;
		end
		else begin
			icache_first_q <= icache_first_d;
			dcache_first_q <= dcache_first_d;
			icache_rd_shift_q <= icache_rd_shift_d;
			dcache_rd_shift_q <= dcache_rd_shift_d;
			icache_rtrn_vld_q <= icache_rtrn_vld_d;
			dcache_rtrn_vld_q <= dcache_rtrn_vld_d;
			icache_rtrn_tid_q <= icache_rtrn_tid_d;
			dcache_rtrn_tid_q <= dcache_rtrn_tid_d;
			dcache_rtrn_type_q <= dcache_rtrn_type_d;
			dcache_rtrn_inv_q <= dcache_rtrn_inv_d;
			amo_off_q <= amo_off_d;
			amo_gen_r_q <= amo_gen_r_d;
		end
	end
	axi_shim #(
		.AxiNumWords(AxiNumWords),
		.AxiIdWidth(4)
	) i_axi_shim(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.rd_req_i(axi_rd_req),
		.rd_gnt_o(axi_rd_gnt),
		.rd_addr_i(axi_rd_addr),
		.rd_blen_i(axi_rd_blen),
		.rd_size_i(axi_rd_size),
		.rd_id_i(axi_rd_id_in),
		.rd_rdy_i(axi_rd_rdy),
		.rd_lock_i(axi_rd_lock),
		.rd_last_o(axi_rd_last),
		.rd_valid_o(axi_rd_valid),
		.rd_data_o(axi_rd_data),
		.rd_id_o(axi_rd_id_out),
		.rd_exokay_o(axi_rd_exokay),
		.wr_req_i(axi_wr_req),
		.wr_gnt_o(axi_wr_gnt),
		.wr_addr_i(axi_wr_addr),
		.wr_data_i(axi_wr_data),
		.wr_be_i(axi_wr_be),
		.wr_blen_i(axi_wr_blen),
		.wr_size_i(axi_wr_size),
		.wr_id_i(axi_wr_id_in),
		.wr_lock_i(axi_wr_lock),
		.wr_atop_i(axi_wr_atop),
		.wr_rdy_i(axi_wr_rdy),
		.wr_valid_o(axi_wr_valid),
		.wr_id_o(axi_wr_id_out),
		.wr_exokay_o(axi_wr_exokay),
		.axi_req_o(axi_req_o),
		.axi_resp_i(axi_resp_i)
	);
endmodule
module axi_res_tbl (
	clk_i,
	rst_ni,
	clr_addr_i,
	clr_req_i,
	clr_gnt_o,
	set_addr_i,
	set_id_i,
	set_req_i,
	set_gnt_o,
	check_addr_i,
	check_id_i,
	check_res_o,
	check_req_i,
	check_gnt_o
);
	parameter [31:0] AXI_ADDR_WIDTH = 0;
	parameter [31:0] AXI_ID_WIDTH = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire [AXI_ADDR_WIDTH - 1:0] clr_addr_i;
	input wire clr_req_i;
	output reg clr_gnt_o;
	input wire [AXI_ADDR_WIDTH - 1:0] set_addr_i;
	input wire [AXI_ID_WIDTH - 1:0] set_id_i;
	input wire set_req_i;
	output reg set_gnt_o;
	input wire [AXI_ADDR_WIDTH - 1:0] check_addr_i;
	input wire [AXI_ID_WIDTH - 1:0] check_id_i;
	output reg check_res_o;
	input wire check_req_i;
	output reg check_gnt_o;
	localparam integer N_IDS = 2 ** AXI_ID_WIDTH;
	reg [(N_IDS * AXI_ADDR_WIDTH) - 1:0] tbl_d;
	reg [(N_IDS * AXI_ADDR_WIDTH) - 1:0] tbl_q;
	reg clr;
	reg set;
	genvar i;
	generate
		for (i = 0; i < N_IDS; i = i + 1) begin : gen_tbl
			always @(*) begin
				tbl_d[i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH] = tbl_q[i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH];
				if (set && (i == set_id_i))
					tbl_d[i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH] = set_addr_i;
				else if (clr && (tbl_q[i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH] == clr_addr_i))
					tbl_d[i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH] = 1'sb0;
			end
		end
	endgenerate
	always @(*) begin
		clr = 1'b0;
		set = 1'b0;
		clr_gnt_o = 1'b0;
		set_gnt_o = 1'b0;
		check_res_o = 1'b0;
		check_gnt_o = 1'b0;
		if (clr_req_i) begin
			clr = 1'b1;
			clr_gnt_o = 1'b1;
		end
		else if (set_req_i) begin
			set = 1'b1;
			set_gnt_o = 1'b1;
		end
		else if (check_req_i) begin
			check_res_o = tbl_q[check_id_i * AXI_ADDR_WIDTH+:AXI_ADDR_WIDTH] == check_addr_i;
			check_gnt_o = 1'b1;
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			tbl_q <= 1'sb0;
		else
			tbl_q <= tbl_d;
endmodule
module axi_riscv_amos_alu (
	amo_op_i,
	amo_operand_a_i,
	amo_operand_b_i,
	amo_result_o
);
	parameter [31:0] DATA_WIDTH = 0;
	input wire [5:0] amo_op_i;
	input wire [DATA_WIDTH - 1:0] amo_operand_a_i;
	input wire [DATA_WIDTH - 1:0] amo_operand_b_i;
	output reg [DATA_WIDTH - 1:0] amo_result_o;
	wire [DATA_WIDTH:0] adder_sum;
	reg [DATA_WIDTH:0] adder_operand_a;
	reg [DATA_WIDTH:0] adder_operand_b;
	assign adder_sum = adder_operand_a + adder_operand_b;
	localparam axi_pkg_ATOP_ADD = 3'b000;
	localparam axi_pkg_ATOP_ATOMICLOAD = 2'b10;
	localparam axi_pkg_ATOP_ATOMICSTORE = 2'b01;
	localparam axi_pkg_ATOP_ATOMICSWAP = 6'b110000;
	localparam axi_pkg_ATOP_CLR = 3'b001;
	localparam axi_pkg_ATOP_EOR = 3'b010;
	localparam axi_pkg_ATOP_SET = 3'b011;
	localparam axi_pkg_ATOP_SMAX = 3'b100;
	localparam axi_pkg_ATOP_SMIN = 3'b101;
	localparam axi_pkg_ATOP_UMAX = 3'b110;
	localparam axi_pkg_ATOP_UMIN = 3'b111;
	always @(*) begin
		adder_operand_a = $signed(amo_operand_a_i);
		adder_operand_b = $signed(amo_operand_b_i);
		amo_result_o = amo_operand_a_i;
		if (amo_op_i == axi_pkg_ATOP_ATOMICSWAP)
			amo_result_o = amo_operand_b_i;
		else if ((amo_op_i[5:4] == axi_pkg_ATOP_ATOMICLOAD) | (amo_op_i[5:4] == axi_pkg_ATOP_ATOMICSTORE))
			case (amo_op_i[2:0])
				axi_pkg_ATOP_ADD: amo_result_o = adder_sum[DATA_WIDTH - 1:0];
				axi_pkg_ATOP_CLR: amo_result_o = amo_operand_a_i & ~amo_operand_b_i;
				axi_pkg_ATOP_SET: amo_result_o = amo_operand_a_i | amo_operand_b_i;
				axi_pkg_ATOP_EOR: amo_result_o = amo_operand_a_i ^ amo_operand_b_i;
				axi_pkg_ATOP_SMAX: begin
					adder_operand_b = -$signed(amo_operand_b_i);
					amo_result_o = (adder_sum[DATA_WIDTH] ? amo_operand_b_i : amo_operand_a_i);
				end
				axi_pkg_ATOP_SMIN: begin
					adder_operand_b = -$signed(amo_operand_b_i);
					amo_result_o = (adder_sum[DATA_WIDTH] ? amo_operand_a_i : amo_operand_b_i);
				end
				axi_pkg_ATOP_UMAX: begin
					adder_operand_a = $unsigned(amo_operand_a_i);
					adder_operand_b = -$unsigned(amo_operand_b_i);
					amo_result_o = (adder_sum[DATA_WIDTH] ? amo_operand_b_i : amo_operand_a_i);
				end
				axi_pkg_ATOP_UMIN: begin
					adder_operand_a = $unsigned(amo_operand_a_i);
					adder_operand_b = -$unsigned(amo_operand_b_i);
					amo_result_o = (adder_sum[DATA_WIDTH] ? amo_operand_a_i : amo_operand_b_i);
				end
				default: amo_result_o = 1'sb0;
			endcase
	end
endmodule
module axi_riscv_amos (
	clk_i,
	rst_ni,
	slv_aw_addr_i,
	slv_aw_prot_i,
	slv_aw_region_i,
	slv_aw_atop_i,
	slv_aw_len_i,
	slv_aw_size_i,
	slv_aw_burst_i,
	slv_aw_lock_i,
	slv_aw_cache_i,
	slv_aw_qos_i,
	slv_aw_id_i,
	slv_aw_user_i,
	slv_aw_ready_o,
	slv_aw_valid_i,
	slv_ar_addr_i,
	slv_ar_prot_i,
	slv_ar_region_i,
	slv_ar_len_i,
	slv_ar_size_i,
	slv_ar_burst_i,
	slv_ar_lock_i,
	slv_ar_cache_i,
	slv_ar_qos_i,
	slv_ar_id_i,
	slv_ar_user_i,
	slv_ar_ready_o,
	slv_ar_valid_i,
	slv_w_data_i,
	slv_w_strb_i,
	slv_w_user_i,
	slv_w_last_i,
	slv_w_ready_o,
	slv_w_valid_i,
	slv_r_data_o,
	slv_r_resp_o,
	slv_r_last_o,
	slv_r_id_o,
	slv_r_user_o,
	slv_r_ready_i,
	slv_r_valid_o,
	slv_b_resp_o,
	slv_b_id_o,
	slv_b_user_o,
	slv_b_ready_i,
	slv_b_valid_o,
	mst_aw_addr_o,
	mst_aw_prot_o,
	mst_aw_region_o,
	mst_aw_atop_o,
	mst_aw_len_o,
	mst_aw_size_o,
	mst_aw_burst_o,
	mst_aw_lock_o,
	mst_aw_cache_o,
	mst_aw_qos_o,
	mst_aw_id_o,
	mst_aw_user_o,
	mst_aw_ready_i,
	mst_aw_valid_o,
	mst_ar_addr_o,
	mst_ar_prot_o,
	mst_ar_region_o,
	mst_ar_len_o,
	mst_ar_size_o,
	mst_ar_burst_o,
	mst_ar_lock_o,
	mst_ar_cache_o,
	mst_ar_qos_o,
	mst_ar_id_o,
	mst_ar_user_o,
	mst_ar_ready_i,
	mst_ar_valid_o,
	mst_w_data_o,
	mst_w_strb_o,
	mst_w_user_o,
	mst_w_last_o,
	mst_w_ready_i,
	mst_w_valid_o,
	mst_r_data_i,
	mst_r_resp_i,
	mst_r_last_i,
	mst_r_id_i,
	mst_r_user_i,
	mst_r_ready_o,
	mst_r_valid_i,
	mst_b_resp_i,
	mst_b_id_i,
	mst_b_user_i,
	mst_b_ready_o,
	mst_b_valid_i
);
	parameter [31:0] AXI_ADDR_WIDTH = 0;
	parameter [31:0] AXI_DATA_WIDTH = 0;
	parameter [31:0] AXI_ID_WIDTH = 0;
	parameter [31:0] AXI_USER_WIDTH = 0;
	parameter [31:0] AXI_MAX_WRITE_TXNS = 0;
	parameter [31:0] RISCV_WORD_WIDTH = 0;
	localparam [31:0] AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
	input wire clk_i;
	input wire rst_ni;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_aw_addr_i;
	input wire [2:0] slv_aw_prot_i;
	input wire [3:0] slv_aw_region_i;
	input wire [5:0] slv_aw_atop_i;
	input wire [7:0] slv_aw_len_i;
	input wire [2:0] slv_aw_size_i;
	input wire [1:0] slv_aw_burst_i;
	input wire slv_aw_lock_i;
	input wire [3:0] slv_aw_cache_i;
	input wire [3:0] slv_aw_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_aw_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_aw_user_i;
	output reg slv_aw_ready_o;
	input wire slv_aw_valid_i;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_ar_addr_i;
	input wire [2:0] slv_ar_prot_i;
	input wire [3:0] slv_ar_region_i;
	input wire [7:0] slv_ar_len_i;
	input wire [2:0] slv_ar_size_i;
	input wire [1:0] slv_ar_burst_i;
	input wire slv_ar_lock_i;
	input wire [3:0] slv_ar_cache_i;
	input wire [3:0] slv_ar_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_ar_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_ar_user_i;
	output reg slv_ar_ready_o;
	input wire slv_ar_valid_i;
	input wire [AXI_DATA_WIDTH - 1:0] slv_w_data_i;
	input wire [AXI_STRB_WIDTH - 1:0] slv_w_strb_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_w_user_i;
	input wire slv_w_last_i;
	output reg slv_w_ready_o;
	input wire slv_w_valid_i;
	output reg [AXI_DATA_WIDTH - 1:0] slv_r_data_o;
	output reg [1:0] slv_r_resp_o;
	output reg slv_r_last_o;
	output reg [AXI_ID_WIDTH - 1:0] slv_r_id_o;
	output reg [AXI_USER_WIDTH - 1:0] slv_r_user_o;
	input wire slv_r_ready_i;
	output reg slv_r_valid_o;
	output reg [1:0] slv_b_resp_o;
	output reg [AXI_ID_WIDTH - 1:0] slv_b_id_o;
	output reg [AXI_USER_WIDTH - 1:0] slv_b_user_o;
	input wire slv_b_ready_i;
	output reg slv_b_valid_o;
	output reg [AXI_ADDR_WIDTH - 1:0] mst_aw_addr_o;
	output reg [2:0] mst_aw_prot_o;
	output reg [3:0] mst_aw_region_o;
	output reg [5:0] mst_aw_atop_o;
	output reg [7:0] mst_aw_len_o;
	output reg [2:0] mst_aw_size_o;
	output reg [1:0] mst_aw_burst_o;
	output reg mst_aw_lock_o;
	output reg [3:0] mst_aw_cache_o;
	output reg [3:0] mst_aw_qos_o;
	output reg [AXI_ID_WIDTH - 1:0] mst_aw_id_o;
	output reg [AXI_USER_WIDTH - 1:0] mst_aw_user_o;
	input wire mst_aw_ready_i;
	output reg mst_aw_valid_o;
	output reg [AXI_ADDR_WIDTH - 1:0] mst_ar_addr_o;
	output reg [2:0] mst_ar_prot_o;
	output reg [3:0] mst_ar_region_o;
	output reg [7:0] mst_ar_len_o;
	output reg [2:0] mst_ar_size_o;
	output reg [1:0] mst_ar_burst_o;
	output reg mst_ar_lock_o;
	output reg [3:0] mst_ar_cache_o;
	output reg [3:0] mst_ar_qos_o;
	output reg [AXI_ID_WIDTH - 1:0] mst_ar_id_o;
	output reg [AXI_USER_WIDTH - 1:0] mst_ar_user_o;
	input wire mst_ar_ready_i;
	output reg mst_ar_valid_o;
	output reg [AXI_DATA_WIDTH - 1:0] mst_w_data_o;
	output reg [AXI_STRB_WIDTH - 1:0] mst_w_strb_o;
	output reg [AXI_USER_WIDTH - 1:0] mst_w_user_o;
	output reg mst_w_last_o;
	input wire mst_w_ready_i;
	output reg mst_w_valid_o;
	input wire [AXI_DATA_WIDTH - 1:0] mst_r_data_i;
	input wire [1:0] mst_r_resp_i;
	input wire mst_r_last_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_r_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_r_user_i;
	output reg mst_r_ready_o;
	input wire mst_r_valid_i;
	input wire [1:0] mst_b_resp_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_b_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_b_user_i;
	output reg mst_b_ready_o;
	input wire mst_b_valid_i;
	localparam [31:0] OUTSTND_BURSTS_WIDTH = $clog2(AXI_MAX_WRITE_TXNS + 1);
	localparam [31:0] AXI_ALU_RATIO = AXI_DATA_WIDTH / RISCV_WORD_WIDTH;
	reg [1:0] aw_state_d;
	reg [1:0] aw_state_q;
	reg [2:0] w_state_d;
	reg [2:0] w_state_q;
	reg [1:0] b_state_d;
	reg [1:0] b_state_q;
	reg [1:0] ar_state_d;
	reg [1:0] ar_state_q;
	reg [1:0] r_state_d;
	reg [1:0] r_state_q;
	reg [1:0] atop_valid_d;
	reg [1:0] atop_valid_q;
	reg [AXI_ADDR_WIDTH - 1:0] addr_d;
	reg [AXI_ADDR_WIDTH - 1:0] addr_q;
	reg [AXI_ID_WIDTH - 1:0] id_d;
	reg [AXI_ID_WIDTH - 1:0] id_q;
	reg [AXI_STRB_WIDTH - 1:0] strb_d;
	reg [AXI_STRB_WIDTH - 1:0] strb_q;
	reg [2:0] size_d;
	reg [2:0] size_q;
	reg [5:0] atop_d;
	reg [5:0] atop_q;
	reg [3:0] cache_d;
	reg [3:0] cache_q;
	reg [2:0] prot_d;
	reg [2:0] prot_q;
	reg [3:0] qos_d;
	reg [3:0] qos_q;
	reg [3:0] region_d;
	reg [3:0] region_q;
	reg [1:0] r_resp_d;
	reg [1:0] r_resp_q;
	reg [AXI_USER_WIDTH - 1:0] aw_user_d;
	reg [AXI_USER_WIDTH - 1:0] aw_user_q;
	reg [AXI_USER_WIDTH - 1:0] w_user_d;
	reg [AXI_USER_WIDTH - 1:0] w_user_q;
	reg [AXI_USER_WIDTH - 1:0] r_user_d;
	reg [AXI_USER_WIDTH - 1:0] r_user_q;
	reg [AXI_DATA_WIDTH - 1:0] w_data_d;
	reg [AXI_DATA_WIDTH - 1:0] w_data_q;
	reg [AXI_DATA_WIDTH - 1:0] r_data_d;
	reg [AXI_DATA_WIDTH - 1:0] r_data_q;
	reg [AXI_DATA_WIDTH - 1:0] result_d;
	reg [AXI_DATA_WIDTH - 1:0] result_q;
	reg w_d_valid_d;
	reg w_d_valid_q;
	reg r_d_valid_d;
	reg r_d_valid_q;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_d;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_q;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_req_d;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_req_q;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_inj_d;
	reg [OUTSTND_BURSTS_WIDTH - 1:0] w_cnt_inj_q;
	wire adapter_ready;
	wire transaction_collision;
	reg aw_valid;
	reg aw_ready;
	wire aw_free;
	reg w_valid;
	reg w_ready;
	wire w_free;
	reg b_valid;
	reg b_ready;
	wire b_free;
	reg ar_valid;
	reg ar_ready;
	wire ar_free;
	reg r_valid;
	reg r_ready;
	wire r_free;
	reg [RISCV_WORD_WIDTH - 1:0] alu_operand_a;
	reg [RISCV_WORD_WIDTH - 1:0] alu_operand_b;
	wire [RISCV_WORD_WIDTH - 1:0] alu_result;
	wire [AXI_DATA_WIDTH - 1:0] alu_result_ext;
	wire [(AXI_ALU_RATIO * RISCV_WORD_WIDTH) - 1:0] op_a;
	wire [(AXI_ALU_RATIO * RISCV_WORD_WIDTH) - 1:0] op_b;
	reg [(AXI_ALU_RATIO * RISCV_WORD_WIDTH) - 1:0] op_a_sign_ext;
	reg [(AXI_ALU_RATIO * RISCV_WORD_WIDTH) - 1:0] op_b_sign_ext;
	reg [(AXI_ALU_RATIO * RISCV_WORD_WIDTH) - 1:0] res;
	reg [(AXI_STRB_WIDTH * 8) - 1:0] strb_ext;
	wire sign_a;
	wire sign_b;
	assign adapter_ready = ((((aw_state_q == 2'd0) && (w_state_q == 3'd0)) && (b_state_q == 2'd0)) && (ar_state_q == 2'd0)) && (r_state_q == 2'd0);
	assign aw_free = ~aw_valid | aw_ready;
	assign w_free = ~w_valid | w_ready;
	assign b_free = ~b_valid | b_ready;
	assign ar_free = ~ar_valid | ar_ready;
	assign r_free = ~r_valid | r_ready;
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			aw_valid <= 0;
			aw_ready <= 0;
			w_valid <= 0;
			w_ready <= 0;
			b_valid <= 0;
			b_ready <= 0;
			ar_valid <= 0;
			ar_ready <= 0;
			r_valid <= 0;
			r_ready <= 0;
		end
		else begin
			aw_valid <= mst_aw_valid_o;
			aw_ready <= mst_aw_ready_i;
			w_valid <= mst_w_valid_o;
			w_ready <= mst_w_ready_i;
			b_valid <= slv_b_valid_o;
			b_ready <= slv_b_ready_i;
			ar_valid <= mst_ar_valid_o;
			ar_ready <= mst_ar_ready_i;
			r_valid <= slv_r_valid_o;
			r_ready <= slv_r_ready_i;
		end
	assign transaction_collision = (slv_aw_addr_i < (addr_q + (8'h01 << size_q))) & (addr_q < (slv_aw_addr_i + (8'h01 << slv_aw_size_i)));
	localparam axi_pkg_ATOP_ATOMICLOAD = 2'b10;
	localparam axi_pkg_ATOP_ATOMICSTORE = 2'b01;
	localparam axi_pkg_ATOP_ATOMICSWAP = 6'b110000;
	localparam axi_pkg_ATOP_LITTLE_END = 1'b0;
	always @(*) begin : calc_atop_valid
		atop_valid_d = atop_valid_q;
		if (adapter_ready) begin
			atop_valid_d = 2'd0;
			if (slv_aw_valid_i && slv_aw_atop_i) begin
				atop_valid_d = 2'd1;
				if ((slv_aw_atop_i == axi_pkg_ATOP_ATOMICSWAP) || (slv_aw_atop_i[5:3] == {axi_pkg_ATOP_ATOMICLOAD, axi_pkg_ATOP_LITTLE_END}))
					atop_valid_d = 2'd2;
				if (slv_aw_atop_i[5:3] == {axi_pkg_ATOP_ATOMICSTORE, axi_pkg_ATOP_LITTLE_END})
					atop_valid_d = 2'd3;
				if (slv_aw_len_i | slv_aw_lock_i)
					atop_valid_d = 2'd1;
				if (slv_aw_size_i > $clog2(RISCV_WORD_WIDTH / 8))
					atop_valid_d = 2'd1;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni) begin : proc_atop_valid
		if (~rst_ni)
			atop_valid_q <= 2'd0;
		else
			atop_valid_q <= atop_valid_d;
	end
	always @(*) begin : axi_aw_channel
		mst_aw_id_o = slv_aw_id_i;
		mst_aw_addr_o = slv_aw_addr_i;
		mst_aw_len_o = slv_aw_len_i;
		mst_aw_size_o = slv_aw_size_i;
		mst_aw_burst_o = slv_aw_burst_i;
		mst_aw_lock_o = slv_aw_lock_i;
		mst_aw_cache_o = slv_aw_cache_i;
		mst_aw_prot_o = slv_aw_prot_i;
		mst_aw_qos_o = slv_aw_qos_i;
		mst_aw_region_o = slv_aw_region_i;
		mst_aw_atop_o = 6'b000000;
		mst_aw_user_o = slv_aw_user_i;
		addr_d = addr_q;
		id_d = id_q;
		size_d = size_q;
		atop_d = atop_q;
		cache_d = cache_q;
		prot_d = prot_q;
		qos_d = qos_q;
		region_d = region_q;
		aw_user_d = aw_user_q;
		w_cnt_inj_d = w_cnt_inj_q;
		aw_state_d = aw_state_q;
		if (slv_aw_valid_i && slv_aw_atop_i) begin
			mst_aw_valid_o = 1'b0;
			slv_aw_ready_o = 1'b0;
		end
		else if (w_cnt_q == AXI_MAX_WRITE_TXNS) begin
			mst_aw_valid_o = 1'b0;
			slv_aw_ready_o = 1'b0;
		end
		else if ((slv_aw_valid_i && transaction_collision) && !adapter_ready) begin
			mst_aw_valid_o = 1'b0;
			slv_aw_ready_o = 1'b0;
		end
		else begin
			mst_aw_valid_o = slv_aw_valid_i;
			slv_aw_ready_o = mst_aw_ready_i;
		end
		if (((w_cnt_inj_q && mst_w_valid_o) && mst_w_ready_i) && mst_w_last_o)
			w_cnt_inj_d = w_cnt_inj_q - 1;
		case (aw_state_q)
			2'd0:
				if ((slv_aw_valid_i && slv_aw_atop_i) && adapter_ready) begin
					slv_aw_ready_o = 1'b1;
					atop_d = slv_aw_atop_i;
					addr_d = slv_aw_addr_i;
					id_d = slv_aw_id_i;
					size_d = slv_aw_size_i;
					cache_d = slv_aw_cache_i;
					prot_d = slv_aw_prot_i;
					qos_d = slv_aw_qos_i;
					region_d = slv_aw_region_i;
					aw_user_d = slv_aw_user_i;
					if (atop_valid_d != 2'd1)
						aw_state_d = 2'd1;
				end
			2'd1, 2'd2:
				if (((r_d_valid_q && w_d_valid_q) && aw_free) || (aw_state_q == 2'd2)) begin
					slv_aw_ready_o = 1'b0;
					mst_aw_valid_o = 1'b1;
					mst_aw_addr_o = addr_q;
					mst_aw_len_o = 8'h00;
					mst_aw_id_o = id_q;
					mst_aw_size_o = size_q;
					mst_aw_burst_o = 2'b00;
					mst_aw_lock_o = 1'b0;
					mst_aw_cache_o = cache_q;
					mst_aw_prot_o = prot_q;
					mst_aw_qos_o = qos_q;
					mst_aw_region_o = region_q;
					mst_aw_user_o = aw_user_q;
					if (mst_aw_ready_i)
						aw_state_d = 2'd0;
					else
						aw_state_d = 2'd2;
					if (aw_state_q == 2'd1) begin
						if (((w_cnt_q && mst_w_valid_o) && mst_w_ready_i) && mst_w_last_o)
							w_cnt_inj_d = w_cnt_q - 1;
						else
							w_cnt_inj_d = w_cnt_q;
					end
				end
			default: aw_state_d = 2'd0;
		endcase
	end
	always @(*) begin : axi_w_channel
		mst_w_data_o = slv_w_data_i;
		mst_w_strb_o = slv_w_strb_i;
		mst_w_last_o = slv_w_last_i;
		mst_w_user_o = slv_w_user_i;
		strb_d = strb_q;
		w_user_d = w_user_q;
		w_data_d = w_data_q;
		result_d = result_q;
		w_d_valid_d = w_d_valid_q;
		w_cnt_req_d = w_cnt_req_q;
		w_state_d = w_state_q;
		if (w_cnt_q == 0) begin
			slv_w_ready_o = 1'b0;
			mst_w_valid_o = 1'b0;
		end
		else begin
			mst_w_valid_o = slv_w_valid_i;
			slv_w_ready_o = mst_w_ready_i;
		end
		case (w_state_q)
			3'd0:
				if (adapter_ready) begin
					w_d_valid_d = 1'b0;
					result_d = 1'sb0;
					if (atop_valid_d != 2'd0) begin
						if (w_cnt_q == 0) begin
							mst_w_valid_o = 1'b0;
							slv_w_ready_o = 1'b1;
							if (slv_w_valid_i) begin
								if (atop_valid_d != 2'd1) begin
									w_data_d = slv_w_data_i;
									strb_d = slv_w_strb_i;
									w_user_d = slv_w_user_i;
									w_d_valid_d = 1'b1;
									w_state_d = 3'd2;
								end
							end
							else begin
								w_cnt_req_d = 1'sb0;
								w_state_d = 3'd1;
							end
						end
						else begin
							if ((mst_w_valid_o && mst_w_ready_i) && mst_w_last_o)
								w_cnt_req_d = w_cnt_q - 1;
							else
								w_cnt_req_d = w_cnt_q;
							w_state_d = 3'd1;
						end
					end
				end
			3'd1:
				if (w_cnt_req_q == 0) begin
					mst_w_valid_o = 1'b0;
					slv_w_ready_o = 1'b1;
					if (slv_w_valid_i) begin
						if (atop_valid_q == 2'd1)
							w_state_d = 3'd0;
						else begin
							w_data_d = slv_w_data_i;
							strb_d = slv_w_strb_i;
							w_user_d = slv_w_user_i;
							w_d_valid_d = 1'b1;
							w_state_d = 3'd2;
						end
					end
				end
				else if ((mst_w_valid_o && mst_w_ready_i) && mst_w_last_o)
					w_cnt_req_d = w_cnt_req_q - 1;
			3'd2:
				if ((r_d_valid_q && w_d_valid_q) && aw_free) begin
					result_d = alu_result_ext;
					if (w_free && (w_cnt_q == 0)) begin
						slv_w_ready_o = 1'b0;
						mst_w_valid_o = 1'b1;
						mst_w_data_o = alu_result_ext;
						mst_w_last_o = 1'b1;
						mst_w_strb_o = strb_q;
						mst_w_user_o = w_user_q;
						if (mst_w_ready_i)
							w_state_d = 3'd0;
						else
							w_state_d = 3'd4;
					end
					else
						w_state_d = 3'd3;
				end
			3'd3, 3'd4:
				if ((w_free && (w_cnt_inj_q == 0)) || (w_state_q == 3'd4)) begin
					slv_w_ready_o = 1'b0;
					mst_w_valid_o = 1'b1;
					mst_w_data_o = result_q;
					mst_w_last_o = 1'b1;
					mst_w_strb_o = strb_q;
					mst_w_user_o = w_user_q;
					if (mst_w_ready_i)
						w_state_d = 3'd0;
					else
						w_state_d = 3'd4;
				end
			default: w_state_d = 3'd0;
		endcase
	end
	localparam axi_pkg_RESP_SLVERR = 2'b10;
	always @(*) begin : axi_b_channel
		mst_b_ready_o = slv_b_ready_i;
		slv_b_id_o = mst_b_id_i;
		slv_b_resp_o = mst_b_resp_i;
		slv_b_user_o = mst_b_user_i;
		slv_b_valid_o = mst_b_valid_i;
		b_state_d = b_state_q;
		case (b_state_q)
			2'd0:
				if (adapter_ready) begin
					if ((atop_valid_d == 2'd2) || (atop_valid_d == 2'd3))
						b_state_d = 2'd1;
					else if (atop_valid_d == 2'd1) begin
						if (b_free) begin
							mst_b_ready_o = 1'b0;
							slv_b_valid_o = 1'b1;
							slv_b_id_o = slv_aw_id_i;
							slv_b_resp_o = axi_pkg_RESP_SLVERR;
							slv_b_user_o = 1'sb0;
							if (!slv_b_ready_i)
								b_state_d = 2'd3;
						end
						else
							b_state_d = 2'd2;
					end
				end
			2'd2, 2'd3:
				if (b_free || (b_state_q == 2'd3)) begin
					mst_b_ready_o = 1'b0;
					slv_b_valid_o = 1'b1;
					slv_b_id_o = id_q;
					slv_b_resp_o = axi_pkg_RESP_SLVERR;
					slv_b_user_o = 1'sb0;
					if (slv_b_ready_i)
						b_state_d = 2'd0;
					else
						b_state_d = 2'd3;
				end
			2'd1:
				if (mst_b_valid_i && (mst_b_id_i == id_q))
					b_state_d = 2'd0;
			default: b_state_d = 2'd0;
		endcase
	end
	always @(*) begin
		w_cnt_d = w_cnt_q;
		if (mst_aw_valid_o && mst_aw_ready_i)
			w_cnt_d = w_cnt_d + 1;
		if ((mst_w_valid_o && mst_w_ready_i) && mst_w_last_o)
			w_cnt_d = w_cnt_d - 1;
	end
	always @(posedge clk_i or negedge rst_ni) begin : axi_write_channel_ff
		if (~rst_ni) begin
			aw_state_q <= 2'd0;
			w_state_q <= 3'd0;
			b_state_q <= 2'd0;
			w_cnt_q <= 1'sb0;
			w_cnt_req_q <= 1'sb0;
			w_cnt_inj_q <= 1'sb0;
			addr_q <= 1'sb0;
			id_q <= 1'sb0;
			size_q <= 1'sb0;
			strb_q <= 1'sb0;
			cache_q <= 1'sb0;
			prot_q <= 1'sb0;
			qos_q <= 1'sb0;
			region_q <= 1'sb0;
			aw_user_q <= 1'sb0;
			w_user_q <= 1'sb0;
			w_data_q <= 1'sb0;
			result_q <= 1'sb0;
			w_d_valid_q <= 1'sb0;
			atop_q <= 6'b000000;
		end
		else begin
			aw_state_q <= aw_state_d;
			w_state_q <= w_state_d;
			b_state_q <= b_state_d;
			w_cnt_q <= w_cnt_d;
			w_cnt_req_q <= w_cnt_req_d;
			w_cnt_inj_q <= w_cnt_inj_d;
			addr_q <= addr_d;
			id_q <= id_d;
			size_q <= size_d;
			strb_q <= strb_d;
			cache_q <= cache_d;
			prot_q <= prot_d;
			qos_q <= qos_d;
			region_q <= region_d;
			aw_user_q <= aw_user_d;
			w_user_q <= w_user_d;
			w_data_q <= w_data_d;
			result_q <= result_d;
			w_d_valid_q <= w_d_valid_d;
			atop_q <= atop_d;
		end
	end
	always @(*) begin : axi_ar_channel
		mst_ar_id_o = slv_ar_id_i;
		mst_ar_addr_o = slv_ar_addr_i;
		mst_ar_len_o = slv_ar_len_i;
		mst_ar_size_o = slv_ar_size_i;
		mst_ar_burst_o = slv_ar_burst_i;
		mst_ar_lock_o = slv_ar_lock_i;
		mst_ar_cache_o = slv_ar_cache_i;
		mst_ar_prot_o = slv_ar_prot_i;
		mst_ar_qos_o = slv_ar_qos_i;
		mst_ar_region_o = slv_ar_region_i;
		mst_ar_user_o = slv_ar_user_i;
		mst_ar_valid_o = 1'b0;
		slv_ar_ready_o = 1'b0;
		ar_state_d = ar_state_q;
		case (ar_state_q)
			2'd0: begin
				mst_ar_valid_o = slv_ar_valid_i;
				slv_ar_ready_o = mst_ar_ready_i;
				if (adapter_ready) begin
					if ((atop_valid_d == 2'd2) | (atop_valid_d == 2'd3)) begin
						if (ar_free) begin
							slv_ar_ready_o = 1'b0;
							mst_ar_valid_o = 1'b1;
							mst_ar_addr_o = slv_aw_addr_i;
							mst_ar_id_o = slv_aw_id_i;
							mst_ar_len_o = 8'h00;
							mst_ar_size_o = slv_aw_size_i;
							mst_ar_burst_o = 2'b00;
							mst_ar_lock_o = 1'h0;
							mst_ar_cache_o = slv_aw_cache_i;
							mst_ar_prot_o = slv_aw_prot_i;
							mst_ar_qos_o = slv_aw_qos_i;
							mst_ar_region_o = slv_aw_region_i;
							mst_ar_user_o = slv_aw_user_i;
							if (!mst_ar_ready_i)
								ar_state_d = 2'd2;
						end
						else
							ar_state_d = 2'd1;
					end
				end
			end
			2'd1, 2'd2:
				if (ar_free || (ar_state_q == 2'd2)) begin
					mst_ar_valid_o = 1'b1;
					mst_ar_addr_o = addr_q;
					mst_ar_id_o = id_q;
					mst_ar_len_o = 8'h00;
					mst_ar_size_o = size_q;
					mst_ar_burst_o = 2'b00;
					mst_ar_lock_o = 1'h0;
					mst_ar_cache_o = cache_q;
					mst_ar_prot_o = prot_q;
					mst_ar_qos_o = qos_q;
					mst_ar_region_o = region_q;
					mst_ar_user_o = aw_user_q;
					if (mst_ar_ready_i)
						ar_state_d = 2'd0;
					else
						ar_state_d = 2'd2;
				end
				else begin
					mst_ar_valid_o = slv_ar_valid_i;
					slv_ar_ready_o = mst_ar_ready_i;
				end
			default: ar_state_d = 2'd0;
		endcase
	end
	always @(*) begin : axi_r_channel
		mst_r_ready_o = slv_r_ready_i;
		slv_r_id_o = mst_r_id_i;
		slv_r_data_o = mst_r_data_i;
		slv_r_resp_o = mst_r_resp_i;
		slv_r_last_o = mst_r_last_i;
		slv_r_user_o = mst_r_user_i;
		slv_r_valid_o = mst_r_valid_i;
		r_data_d = r_data_q;
		r_resp_d = r_resp_q;
		r_user_d = r_user_q;
		r_d_valid_d = r_d_valid_q;
		r_state_d = r_state_q;
		case (r_state_q)
			2'd0:
				if (adapter_ready) begin
					r_d_valid_d = 1'b0;
					if ((atop_valid_d == 2'd2) || (atop_valid_d == 2'd3))
						r_state_d = 2'd1;
					else if (atop_valid_d == 2'd1) begin
						if (r_free) begin
							mst_r_ready_o = 1'b0;
							slv_r_valid_o = 1'b1;
							slv_r_data_o = 1'sb0;
							slv_r_id_o = slv_aw_id_i;
							slv_r_last_o = 1'b1;
							slv_r_resp_o = axi_pkg_RESP_SLVERR;
							slv_r_user_o = 1'sb0;
							if (!slv_r_ready_i)
								r_state_d = 2'd3;
						end
						else
							r_state_d = 2'd2;
					end
				end
			2'd1:
				if (mst_r_valid_i && (mst_r_id_i == id_q)) begin
					mst_r_ready_o = 1'b1;
					slv_r_valid_o = 1'b0;
					r_data_d = mst_r_data_i;
					r_resp_d = mst_r_resp_i;
					r_user_d = mst_r_user_i;
					r_d_valid_d = 1'b1;
					if (atop_valid_q == 2'd3)
						r_state_d = 2'd0;
					else
						r_state_d = 2'd2;
				end
			2'd2, 2'd3:
				if ((r_free && (b_state_q != 2'd1)) || (r_state_q == 2'd3)) begin
					mst_r_ready_o = 1'b0;
					slv_r_valid_o = 1'b1;
					slv_r_data_o = r_data_q;
					slv_r_id_o = id_q;
					slv_r_last_o = 1'b1;
					slv_r_resp_o = r_resp_q;
					slv_r_user_o = r_user_q;
					if (atop_valid_q == 2'd1) begin
						slv_r_data_o = 1'sb0;
						slv_r_resp_o = axi_pkg_RESP_SLVERR;
						slv_r_user_o = 1'sb0;
					end
					if (slv_r_ready_i)
						r_state_d = 2'd0;
					else
						r_state_d = 2'd3;
				end
			default: r_state_d = 2'd0;
		endcase
	end
	always @(posedge clk_i or negedge rst_ni) begin : axi_read_channel_ff
		if (~rst_ni) begin
			ar_state_q <= 2'd0;
			r_state_q <= 2'd0;
			r_data_q <= 1'sb0;
			r_resp_q <= 1'sb0;
			r_user_q <= 1'sb0;
			r_d_valid_q <= 1'b0;
		end
		else begin
			ar_state_q <= ar_state_d;
			r_state_q <= r_state_d;
			r_data_q <= r_data_d;
			r_resp_q <= r_resp_d;
			r_user_q <= r_user_d;
			r_d_valid_q <= r_d_valid_d;
		end
	end
	assign op_a = r_data_q & strb_ext;
	assign op_b = w_data_q & strb_ext;
	assign sign_a = |(op_a & ~(strb_ext >> 1));
	assign sign_b = |(op_b & ~(strb_ext >> 1));
	assign alu_result_ext = res;
	localparam axi_pkg_ATOP_SMAX = 3'b100;
	localparam axi_pkg_ATOP_SMIN = 3'b101;
	generate
		if ((AXI_ALU_RATIO == 1) && (RISCV_WORD_WIDTH == 32)) begin : genblk1
			wire [RISCV_WORD_WIDTH:1] sv2v_tmp_96078;
			assign sv2v_tmp_96078 = op_a;
			always @(*) alu_operand_a = sv2v_tmp_96078;
			wire [RISCV_WORD_WIDTH:1] sv2v_tmp_A90DA;
			assign sv2v_tmp_A90DA = op_b;
			always @(*) alu_operand_b = sv2v_tmp_A90DA;
			wire [AXI_ALU_RATIO * RISCV_WORD_WIDTH:1] sv2v_tmp_7D7E9;
			assign sv2v_tmp_7D7E9 = alu_result;
			always @(*) res = sv2v_tmp_7D7E9;
		end
		else if ((AXI_ALU_RATIO == 1) && (RISCV_WORD_WIDTH == 64)) begin : genblk1
			wire [AXI_ALU_RATIO * RISCV_WORD_WIDTH:1] sv2v_tmp_7D7E9;
			assign sv2v_tmp_7D7E9 = alu_result;
			always @(*) res = sv2v_tmp_7D7E9;
			always @(*) begin
				op_a_sign_ext = op_a | ({AXI_ALU_RATIO * RISCV_WORD_WIDTH {sign_a}} & ~strb_ext);
				op_b_sign_ext = op_b | ({AXI_ALU_RATIO * RISCV_WORD_WIDTH {sign_b}} & ~strb_ext);
				if ((atop_q[2:0] == axi_pkg_ATOP_SMAX) || (atop_q[2:0] == axi_pkg_ATOP_SMIN)) begin
					alu_operand_a = op_a_sign_ext;
					alu_operand_b = op_b_sign_ext;
				end
				else begin
					alu_operand_a = op_a;
					alu_operand_b = op_b;
				end
			end
		end
		else begin : genblk1
			always @(*) begin
				op_a_sign_ext = op_a | ({AXI_ALU_RATIO * RISCV_WORD_WIDTH {sign_a}} & ~strb_ext);
				op_b_sign_ext = op_b | ({AXI_ALU_RATIO * RISCV_WORD_WIDTH {sign_b}} & ~strb_ext);
				if ((atop_q[2:0] == axi_pkg_ATOP_SMAX) || (atop_q[2:0] == axi_pkg_ATOP_SMIN)) begin
					alu_operand_a = op_a_sign_ext[addr_q[$clog2(AXI_DATA_WIDTH / 8) - 1:$clog2(RISCV_WORD_WIDTH / 8)] * RISCV_WORD_WIDTH+:RISCV_WORD_WIDTH];
					alu_operand_b = op_b_sign_ext[addr_q[$clog2(AXI_DATA_WIDTH / 8) - 1:$clog2(RISCV_WORD_WIDTH / 8)] * RISCV_WORD_WIDTH+:RISCV_WORD_WIDTH];
				end
				else begin
					alu_operand_a = op_a[addr_q[$clog2(AXI_DATA_WIDTH / 8) - 1:$clog2(RISCV_WORD_WIDTH / 8)] * RISCV_WORD_WIDTH+:RISCV_WORD_WIDTH];
					alu_operand_b = op_b[addr_q[$clog2(AXI_DATA_WIDTH / 8) - 1:$clog2(RISCV_WORD_WIDTH / 8)] * RISCV_WORD_WIDTH+:RISCV_WORD_WIDTH];
				end
				res = 1'sb0;
				res[addr_q[$clog2(AXI_DATA_WIDTH / 8) - 1:$clog2(RISCV_WORD_WIDTH / 8)] * RISCV_WORD_WIDTH+:RISCV_WORD_WIDTH] = alu_result;
			end
		end
	endgenerate
	genvar i;
	generate
		for (i = 0; i < AXI_STRB_WIDTH; i = i + 1) begin : genblk2
			always @(*)
				if (strb_q[i])
					strb_ext[i * 8+:8] = 8'hff;
				else
					strb_ext[i * 8+:8] = 8'h00;
		end
	endgenerate
	axi_riscv_amos_alu #(.DATA_WIDTH(RISCV_WORD_WIDTH)) i_amo_alu(
		.amo_op_i(atop_q),
		.amo_operand_a_i(alu_operand_a),
		.amo_operand_b_i(alu_operand_b),
		.amo_result_o(alu_result)
	);
endmodule
module axi_riscv_atomics (
	clk_i,
	rst_ni,
	slv_aw_addr_i,
	slv_aw_prot_i,
	slv_aw_region_i,
	slv_aw_atop_i,
	slv_aw_len_i,
	slv_aw_size_i,
	slv_aw_burst_i,
	slv_aw_lock_i,
	slv_aw_cache_i,
	slv_aw_qos_i,
	slv_aw_id_i,
	slv_aw_user_i,
	slv_aw_ready_o,
	slv_aw_valid_i,
	slv_ar_addr_i,
	slv_ar_prot_i,
	slv_ar_region_i,
	slv_ar_len_i,
	slv_ar_size_i,
	slv_ar_burst_i,
	slv_ar_lock_i,
	slv_ar_cache_i,
	slv_ar_qos_i,
	slv_ar_id_i,
	slv_ar_user_i,
	slv_ar_ready_o,
	slv_ar_valid_i,
	slv_w_data_i,
	slv_w_strb_i,
	slv_w_user_i,
	slv_w_last_i,
	slv_w_ready_o,
	slv_w_valid_i,
	slv_r_data_o,
	slv_r_resp_o,
	slv_r_last_o,
	slv_r_id_o,
	slv_r_user_o,
	slv_r_ready_i,
	slv_r_valid_o,
	slv_b_resp_o,
	slv_b_id_o,
	slv_b_user_o,
	slv_b_ready_i,
	slv_b_valid_o,
	mst_aw_addr_o,
	mst_aw_prot_o,
	mst_aw_region_o,
	mst_aw_atop_o,
	mst_aw_len_o,
	mst_aw_size_o,
	mst_aw_burst_o,
	mst_aw_lock_o,
	mst_aw_cache_o,
	mst_aw_qos_o,
	mst_aw_id_o,
	mst_aw_user_o,
	mst_aw_ready_i,
	mst_aw_valid_o,
	mst_ar_addr_o,
	mst_ar_prot_o,
	mst_ar_region_o,
	mst_ar_len_o,
	mst_ar_size_o,
	mst_ar_burst_o,
	mst_ar_lock_o,
	mst_ar_cache_o,
	mst_ar_qos_o,
	mst_ar_id_o,
	mst_ar_user_o,
	mst_ar_ready_i,
	mst_ar_valid_o,
	mst_w_data_o,
	mst_w_strb_o,
	mst_w_user_o,
	mst_w_last_o,
	mst_w_ready_i,
	mst_w_valid_o,
	mst_r_data_i,
	mst_r_resp_i,
	mst_r_last_i,
	mst_r_id_i,
	mst_r_user_i,
	mst_r_ready_o,
	mst_r_valid_i,
	mst_b_resp_i,
	mst_b_id_i,
	mst_b_user_i,
	mst_b_ready_o,
	mst_b_valid_i
);
	parameter [31:0] AXI_ADDR_WIDTH = 0;
	parameter [31:0] AXI_DATA_WIDTH = 0;
	parameter [31:0] AXI_ID_WIDTH = 0;
	parameter [31:0] AXI_USER_WIDTH = 0;
	parameter [31:0] AXI_MAX_WRITE_TXNS = 0;
	parameter [31:0] RISCV_WORD_WIDTH = 0;
	localparam [31:0] AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
	input wire clk_i;
	input wire rst_ni;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_aw_addr_i;
	input wire [2:0] slv_aw_prot_i;
	input wire [3:0] slv_aw_region_i;
	input wire [5:0] slv_aw_atop_i;
	input wire [7:0] slv_aw_len_i;
	input wire [2:0] slv_aw_size_i;
	input wire [1:0] slv_aw_burst_i;
	input wire slv_aw_lock_i;
	input wire [3:0] slv_aw_cache_i;
	input wire [3:0] slv_aw_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_aw_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_aw_user_i;
	output wire slv_aw_ready_o;
	input wire slv_aw_valid_i;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_ar_addr_i;
	input wire [2:0] slv_ar_prot_i;
	input wire [3:0] slv_ar_region_i;
	input wire [7:0] slv_ar_len_i;
	input wire [2:0] slv_ar_size_i;
	input wire [1:0] slv_ar_burst_i;
	input wire slv_ar_lock_i;
	input wire [3:0] slv_ar_cache_i;
	input wire [3:0] slv_ar_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_ar_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_ar_user_i;
	output wire slv_ar_ready_o;
	input wire slv_ar_valid_i;
	input wire [AXI_DATA_WIDTH - 1:0] slv_w_data_i;
	input wire [AXI_STRB_WIDTH - 1:0] slv_w_strb_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_w_user_i;
	input wire slv_w_last_i;
	output wire slv_w_ready_o;
	input wire slv_w_valid_i;
	output wire [AXI_DATA_WIDTH - 1:0] slv_r_data_o;
	output wire [1:0] slv_r_resp_o;
	output wire slv_r_last_o;
	output wire [AXI_ID_WIDTH - 1:0] slv_r_id_o;
	output wire [AXI_USER_WIDTH - 1:0] slv_r_user_o;
	input wire slv_r_ready_i;
	output wire slv_r_valid_o;
	output wire [1:0] slv_b_resp_o;
	output wire [AXI_ID_WIDTH - 1:0] slv_b_id_o;
	output wire [AXI_USER_WIDTH - 1:0] slv_b_user_o;
	input wire slv_b_ready_i;
	output wire slv_b_valid_o;
	output wire [AXI_ADDR_WIDTH - 1:0] mst_aw_addr_o;
	output wire [2:0] mst_aw_prot_o;
	output wire [3:0] mst_aw_region_o;
	output wire [5:0] mst_aw_atop_o;
	output wire [7:0] mst_aw_len_o;
	output wire [2:0] mst_aw_size_o;
	output wire [1:0] mst_aw_burst_o;
	output wire mst_aw_lock_o;
	output wire [3:0] mst_aw_cache_o;
	output wire [3:0] mst_aw_qos_o;
	output wire [AXI_ID_WIDTH - 1:0] mst_aw_id_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_aw_user_o;
	input wire mst_aw_ready_i;
	output wire mst_aw_valid_o;
	output wire [AXI_ADDR_WIDTH - 1:0] mst_ar_addr_o;
	output wire [2:0] mst_ar_prot_o;
	output wire [3:0] mst_ar_region_o;
	output wire [7:0] mst_ar_len_o;
	output wire [2:0] mst_ar_size_o;
	output wire [1:0] mst_ar_burst_o;
	output wire mst_ar_lock_o;
	output wire [3:0] mst_ar_cache_o;
	output wire [3:0] mst_ar_qos_o;
	output wire [AXI_ID_WIDTH - 1:0] mst_ar_id_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_ar_user_o;
	input wire mst_ar_ready_i;
	output wire mst_ar_valid_o;
	output wire [AXI_DATA_WIDTH - 1:0] mst_w_data_o;
	output wire [AXI_STRB_WIDTH - 1:0] mst_w_strb_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_w_user_o;
	output wire mst_w_last_o;
	input wire mst_w_ready_i;
	output wire mst_w_valid_o;
	input wire [AXI_DATA_WIDTH - 1:0] mst_r_data_i;
	input wire [1:0] mst_r_resp_i;
	input wire mst_r_last_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_r_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_r_user_i;
	output wire mst_r_ready_o;
	input wire mst_r_valid_i;
	input wire [1:0] mst_b_resp_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_b_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_b_user_i;
	output wire mst_b_ready_o;
	input wire mst_b_valid_i;
	localparam [63:0] ADDR_BEGIN = 1'sb0;
	localparam [63:0] ADDR_END = {AXI_ADDR_WIDTH {1'b1}};
	wire [AXI_ADDR_WIDTH - 1:0] int_axi_aw_addr;
	wire [2:0] int_axi_aw_prot;
	wire [3:0] int_axi_aw_region;
	wire [5:0] int_axi_aw_atop;
	wire [7:0] int_axi_aw_len;
	wire [2:0] int_axi_aw_size;
	wire [1:0] int_axi_aw_burst;
	wire int_axi_aw_lock;
	wire [3:0] int_axi_aw_cache;
	wire [3:0] int_axi_aw_qos;
	wire [AXI_ID_WIDTH - 1:0] int_axi_aw_id;
	wire [AXI_USER_WIDTH - 1:0] int_axi_aw_user;
	wire int_axi_aw_ready;
	wire int_axi_aw_valid;
	wire [AXI_ADDR_WIDTH - 1:0] int_axi_ar_addr;
	wire [2:0] int_axi_ar_prot;
	wire [3:0] int_axi_ar_region;
	wire [7:0] int_axi_ar_len;
	wire [2:0] int_axi_ar_size;
	wire [1:0] int_axi_ar_burst;
	wire int_axi_ar_lock;
	wire [3:0] int_axi_ar_cache;
	wire [3:0] int_axi_ar_qos;
	wire [AXI_ID_WIDTH - 1:0] int_axi_ar_id;
	wire [AXI_USER_WIDTH - 1:0] int_axi_ar_user;
	wire int_axi_ar_ready;
	wire int_axi_ar_valid;
	wire [AXI_DATA_WIDTH - 1:0] int_axi_w_data;
	wire [AXI_STRB_WIDTH - 1:0] int_axi_w_strb;
	wire [AXI_USER_WIDTH - 1:0] int_axi_w_user;
	wire int_axi_w_last;
	wire int_axi_w_ready;
	wire int_axi_w_valid;
	wire [AXI_DATA_WIDTH - 1:0] int_axi_r_data;
	wire [1:0] int_axi_r_resp;
	wire int_axi_r_last;
	wire [AXI_ID_WIDTH - 1:0] int_axi_r_id;
	wire [AXI_USER_WIDTH - 1:0] int_axi_r_user;
	wire int_axi_r_ready;
	wire int_axi_r_valid;
	wire [1:0] int_axi_b_resp;
	wire [AXI_ID_WIDTH - 1:0] int_axi_b_id;
	wire [AXI_USER_WIDTH - 1:0] int_axi_b_user;
	wire int_axi_b_ready;
	wire int_axi_b_valid;
	axi_riscv_amos #(
		.AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
		.AXI_DATA_WIDTH(AXI_DATA_WIDTH),
		.AXI_ID_WIDTH(AXI_ID_WIDTH),
		.AXI_USER_WIDTH(AXI_USER_WIDTH),
		.AXI_MAX_WRITE_TXNS(AXI_MAX_WRITE_TXNS),
		.RISCV_WORD_WIDTH(RISCV_WORD_WIDTH)
	) i_amos(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.slv_aw_addr_i(slv_aw_addr_i),
		.slv_aw_prot_i(slv_aw_prot_i),
		.slv_aw_region_i(slv_aw_region_i),
		.slv_aw_atop_i(slv_aw_atop_i),
		.slv_aw_len_i(slv_aw_len_i),
		.slv_aw_size_i(slv_aw_size_i),
		.slv_aw_burst_i(slv_aw_burst_i),
		.slv_aw_lock_i(slv_aw_lock_i),
		.slv_aw_cache_i(slv_aw_cache_i),
		.slv_aw_qos_i(slv_aw_qos_i),
		.slv_aw_id_i(slv_aw_id_i),
		.slv_aw_user_i(slv_aw_user_i),
		.slv_aw_ready_o(slv_aw_ready_o),
		.slv_aw_valid_i(slv_aw_valid_i),
		.slv_ar_addr_i(slv_ar_addr_i),
		.slv_ar_prot_i(slv_ar_prot_i),
		.slv_ar_region_i(slv_ar_region_i),
		.slv_ar_len_i(slv_ar_len_i),
		.slv_ar_size_i(slv_ar_size_i),
		.slv_ar_burst_i(slv_ar_burst_i),
		.slv_ar_lock_i(slv_ar_lock_i),
		.slv_ar_cache_i(slv_ar_cache_i),
		.slv_ar_qos_i(slv_ar_qos_i),
		.slv_ar_id_i(slv_ar_id_i),
		.slv_ar_user_i(slv_ar_user_i),
		.slv_ar_ready_o(slv_ar_ready_o),
		.slv_ar_valid_i(slv_ar_valid_i),
		.slv_w_data_i(slv_w_data_i),
		.slv_w_strb_i(slv_w_strb_i),
		.slv_w_user_i(slv_w_user_i),
		.slv_w_last_i(slv_w_last_i),
		.slv_w_ready_o(slv_w_ready_o),
		.slv_w_valid_i(slv_w_valid_i),
		.slv_r_data_o(slv_r_data_o),
		.slv_r_resp_o(slv_r_resp_o),
		.slv_r_last_o(slv_r_last_o),
		.slv_r_id_o(slv_r_id_o),
		.slv_r_user_o(slv_r_user_o),
		.slv_r_ready_i(slv_r_ready_i),
		.slv_r_valid_o(slv_r_valid_o),
		.slv_b_resp_o(slv_b_resp_o),
		.slv_b_id_o(slv_b_id_o),
		.slv_b_user_o(slv_b_user_o),
		.slv_b_ready_i(slv_b_ready_i),
		.slv_b_valid_o(slv_b_valid_o),
		.mst_aw_addr_o(int_axi_aw_addr),
		.mst_aw_prot_o(int_axi_aw_prot),
		.mst_aw_region_o(int_axi_aw_region),
		.mst_aw_atop_o(int_axi_aw_atop),
		.mst_aw_len_o(int_axi_aw_len),
		.mst_aw_size_o(int_axi_aw_size),
		.mst_aw_burst_o(int_axi_aw_burst),
		.mst_aw_lock_o(int_axi_aw_lock),
		.mst_aw_cache_o(int_axi_aw_cache),
		.mst_aw_qos_o(int_axi_aw_qos),
		.mst_aw_id_o(int_axi_aw_id),
		.mst_aw_user_o(int_axi_aw_user),
		.mst_aw_ready_i(int_axi_aw_ready),
		.mst_aw_valid_o(int_axi_aw_valid),
		.mst_ar_addr_o(int_axi_ar_addr),
		.mst_ar_prot_o(int_axi_ar_prot),
		.mst_ar_region_o(int_axi_ar_region),
		.mst_ar_len_o(int_axi_ar_len),
		.mst_ar_size_o(int_axi_ar_size),
		.mst_ar_burst_o(int_axi_ar_burst),
		.mst_ar_lock_o(int_axi_ar_lock),
		.mst_ar_cache_o(int_axi_ar_cache),
		.mst_ar_qos_o(int_axi_ar_qos),
		.mst_ar_id_o(int_axi_ar_id),
		.mst_ar_user_o(int_axi_ar_user),
		.mst_ar_ready_i(int_axi_ar_ready),
		.mst_ar_valid_o(int_axi_ar_valid),
		.mst_w_data_o(int_axi_w_data),
		.mst_w_strb_o(int_axi_w_strb),
		.mst_w_user_o(int_axi_w_user),
		.mst_w_last_o(int_axi_w_last),
		.mst_w_ready_i(int_axi_w_ready),
		.mst_w_valid_o(int_axi_w_valid),
		.mst_r_data_i(int_axi_r_data),
		.mst_r_resp_i(int_axi_r_resp),
		.mst_r_last_i(int_axi_r_last),
		.mst_r_id_i(int_axi_r_id),
		.mst_r_user_i(int_axi_r_user),
		.mst_r_ready_o(int_axi_r_ready),
		.mst_r_valid_i(int_axi_r_valid),
		.mst_b_resp_i(int_axi_b_resp),
		.mst_b_id_i(int_axi_b_id),
		.mst_b_user_i(int_axi_b_user),
		.mst_b_ready_o(int_axi_b_ready),
		.mst_b_valid_i(int_axi_b_valid)
	);
	axi_riscv_lrsc #(
		.ADDR_BEGIN(ADDR_BEGIN),
		.ADDR_END(ADDR_END),
		.AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
		.AXI_DATA_WIDTH(AXI_DATA_WIDTH),
		.AXI_ID_WIDTH(AXI_ID_WIDTH),
		.AXI_USER_WIDTH(AXI_USER_WIDTH)
	) i_lrsc(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.slv_aw_addr_i(int_axi_aw_addr),
		.slv_aw_prot_i(int_axi_aw_prot),
		.slv_aw_region_i(int_axi_aw_region),
		.slv_aw_atop_i(int_axi_aw_atop),
		.slv_aw_len_i(int_axi_aw_len),
		.slv_aw_size_i(int_axi_aw_size),
		.slv_aw_burst_i(int_axi_aw_burst),
		.slv_aw_lock_i(int_axi_aw_lock),
		.slv_aw_cache_i(int_axi_aw_cache),
		.slv_aw_qos_i(int_axi_aw_qos),
		.slv_aw_id_i(int_axi_aw_id),
		.slv_aw_user_i(int_axi_aw_user),
		.slv_aw_ready_o(int_axi_aw_ready),
		.slv_aw_valid_i(int_axi_aw_valid),
		.slv_ar_addr_i(int_axi_ar_addr),
		.slv_ar_prot_i(int_axi_ar_prot),
		.slv_ar_region_i(int_axi_ar_region),
		.slv_ar_len_i(int_axi_ar_len),
		.slv_ar_size_i(int_axi_ar_size),
		.slv_ar_burst_i(int_axi_ar_burst),
		.slv_ar_lock_i(int_axi_ar_lock),
		.slv_ar_cache_i(int_axi_ar_cache),
		.slv_ar_qos_i(int_axi_ar_qos),
		.slv_ar_id_i(int_axi_ar_id),
		.slv_ar_user_i(int_axi_ar_user),
		.slv_ar_ready_o(int_axi_ar_ready),
		.slv_ar_valid_i(int_axi_ar_valid),
		.slv_w_data_i(int_axi_w_data),
		.slv_w_strb_i(int_axi_w_strb),
		.slv_w_user_i(int_axi_w_user),
		.slv_w_last_i(int_axi_w_last),
		.slv_w_ready_o(int_axi_w_ready),
		.slv_w_valid_i(int_axi_w_valid),
		.slv_r_data_o(int_axi_r_data),
		.slv_r_resp_o(int_axi_r_resp),
		.slv_r_last_o(int_axi_r_last),
		.slv_r_id_o(int_axi_r_id),
		.slv_r_user_o(int_axi_r_user),
		.slv_r_ready_i(int_axi_r_ready),
		.slv_r_valid_o(int_axi_r_valid),
		.slv_b_resp_o(int_axi_b_resp),
		.slv_b_id_o(int_axi_b_id),
		.slv_b_user_o(int_axi_b_user),
		.slv_b_ready_i(int_axi_b_ready),
		.slv_b_valid_o(int_axi_b_valid),
		.mst_aw_addr_o(mst_aw_addr_o),
		.mst_aw_prot_o(mst_aw_prot_o),
		.mst_aw_region_o(mst_aw_region_o),
		.mst_aw_atop_o(mst_aw_atop_o),
		.mst_aw_len_o(mst_aw_len_o),
		.mst_aw_size_o(mst_aw_size_o),
		.mst_aw_burst_o(mst_aw_burst_o),
		.mst_aw_lock_o(mst_aw_lock_o),
		.mst_aw_cache_o(mst_aw_cache_o),
		.mst_aw_qos_o(mst_aw_qos_o),
		.mst_aw_id_o(mst_aw_id_o),
		.mst_aw_user_o(mst_aw_user_o),
		.mst_aw_ready_i(mst_aw_ready_i),
		.mst_aw_valid_o(mst_aw_valid_o),
		.mst_ar_addr_o(mst_ar_addr_o),
		.mst_ar_prot_o(mst_ar_prot_o),
		.mst_ar_region_o(mst_ar_region_o),
		.mst_ar_len_o(mst_ar_len_o),
		.mst_ar_size_o(mst_ar_size_o),
		.mst_ar_burst_o(mst_ar_burst_o),
		.mst_ar_lock_o(mst_ar_lock_o),
		.mst_ar_cache_o(mst_ar_cache_o),
		.mst_ar_qos_o(mst_ar_qos_o),
		.mst_ar_id_o(mst_ar_id_o),
		.mst_ar_user_o(mst_ar_user_o),
		.mst_ar_ready_i(mst_ar_ready_i),
		.mst_ar_valid_o(mst_ar_valid_o),
		.mst_w_data_o(mst_w_data_o),
		.mst_w_strb_o(mst_w_strb_o),
		.mst_w_user_o(mst_w_user_o),
		.mst_w_last_o(mst_w_last_o),
		.mst_w_ready_i(mst_w_ready_i),
		.mst_w_valid_o(mst_w_valid_o),
		.mst_r_data_i(mst_r_data_i),
		.mst_r_resp_i(mst_r_resp_i),
		.mst_r_last_i(mst_r_last_i),
		.mst_r_id_i(mst_r_id_i),
		.mst_r_user_i(mst_r_user_i),
		.mst_r_ready_o(mst_r_ready_o),
		.mst_r_valid_i(mst_r_valid_i),
		.mst_b_resp_i(mst_b_resp_i),
		.mst_b_id_i(mst_b_id_i),
		.mst_b_user_i(mst_b_user_i),
		.mst_b_ready_o(mst_b_ready_o),
		.mst_b_valid_i(mst_b_valid_i)
	);
endmodule
module axi_riscv_lrsc (
	clk_i,
	rst_ni,
	slv_aw_addr_i,
	slv_aw_prot_i,
	slv_aw_region_i,
	slv_aw_atop_i,
	slv_aw_len_i,
	slv_aw_size_i,
	slv_aw_burst_i,
	slv_aw_lock_i,
	slv_aw_cache_i,
	slv_aw_qos_i,
	slv_aw_id_i,
	slv_aw_user_i,
	slv_aw_ready_o,
	slv_aw_valid_i,
	slv_ar_addr_i,
	slv_ar_prot_i,
	slv_ar_region_i,
	slv_ar_len_i,
	slv_ar_size_i,
	slv_ar_burst_i,
	slv_ar_lock_i,
	slv_ar_cache_i,
	slv_ar_qos_i,
	slv_ar_id_i,
	slv_ar_user_i,
	slv_ar_ready_o,
	slv_ar_valid_i,
	slv_w_data_i,
	slv_w_strb_i,
	slv_w_user_i,
	slv_w_last_i,
	slv_w_ready_o,
	slv_w_valid_i,
	slv_r_data_o,
	slv_r_resp_o,
	slv_r_last_o,
	slv_r_id_o,
	slv_r_user_o,
	slv_r_ready_i,
	slv_r_valid_o,
	slv_b_resp_o,
	slv_b_id_o,
	slv_b_user_o,
	slv_b_ready_i,
	slv_b_valid_o,
	mst_aw_addr_o,
	mst_aw_prot_o,
	mst_aw_region_o,
	mst_aw_atop_o,
	mst_aw_len_o,
	mst_aw_size_o,
	mst_aw_burst_o,
	mst_aw_lock_o,
	mst_aw_cache_o,
	mst_aw_qos_o,
	mst_aw_id_o,
	mst_aw_user_o,
	mst_aw_ready_i,
	mst_aw_valid_o,
	mst_ar_addr_o,
	mst_ar_prot_o,
	mst_ar_region_o,
	mst_ar_len_o,
	mst_ar_size_o,
	mst_ar_burst_o,
	mst_ar_lock_o,
	mst_ar_cache_o,
	mst_ar_qos_o,
	mst_ar_id_o,
	mst_ar_user_o,
	mst_ar_ready_i,
	mst_ar_valid_o,
	mst_w_data_o,
	mst_w_strb_o,
	mst_w_user_o,
	mst_w_last_o,
	mst_w_ready_i,
	mst_w_valid_o,
	mst_r_data_i,
	mst_r_resp_i,
	mst_r_last_i,
	mst_r_id_i,
	mst_r_user_i,
	mst_r_ready_o,
	mst_r_valid_i,
	mst_b_resp_i,
	mst_b_id_i,
	mst_b_user_i,
	mst_b_ready_o,
	mst_b_valid_i
);
	parameter [63:0] ADDR_BEGIN = 0;
	parameter [63:0] ADDR_END = 0;
	parameter [31:0] AXI_ADDR_WIDTH = 0;
	parameter [31:0] AXI_DATA_WIDTH = 0;
	parameter [31:0] AXI_ID_WIDTH = 0;
	parameter [31:0] AXI_USER_WIDTH = 0;
	localparam [31:0] AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
	input wire clk_i;
	input wire rst_ni;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_aw_addr_i;
	input wire [2:0] slv_aw_prot_i;
	input wire [3:0] slv_aw_region_i;
	input wire [5:0] slv_aw_atop_i;
	input wire [7:0] slv_aw_len_i;
	input wire [2:0] slv_aw_size_i;
	input wire [1:0] slv_aw_burst_i;
	input wire slv_aw_lock_i;
	input wire [3:0] slv_aw_cache_i;
	input wire [3:0] slv_aw_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_aw_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_aw_user_i;
	output reg slv_aw_ready_o;
	input wire slv_aw_valid_i;
	input wire [AXI_ADDR_WIDTH - 1:0] slv_ar_addr_i;
	input wire [2:0] slv_ar_prot_i;
	input wire [3:0] slv_ar_region_i;
	input wire [7:0] slv_ar_len_i;
	input wire [2:0] slv_ar_size_i;
	input wire [1:0] slv_ar_burst_i;
	input wire slv_ar_lock_i;
	input wire [3:0] slv_ar_cache_i;
	input wire [3:0] slv_ar_qos_i;
	input wire [AXI_ID_WIDTH - 1:0] slv_ar_id_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_ar_user_i;
	output reg slv_ar_ready_o;
	input wire slv_ar_valid_i;
	input wire [AXI_DATA_WIDTH - 1:0] slv_w_data_i;
	input wire [AXI_STRB_WIDTH - 1:0] slv_w_strb_i;
	input wire [AXI_USER_WIDTH - 1:0] slv_w_user_i;
	input wire slv_w_last_i;
	output reg slv_w_ready_o;
	input wire slv_w_valid_i;
	output wire [AXI_DATA_WIDTH - 1:0] slv_r_data_o;
	output reg [1:0] slv_r_resp_o;
	output wire slv_r_last_o;
	output wire [AXI_ID_WIDTH - 1:0] slv_r_id_o;
	output wire [AXI_USER_WIDTH - 1:0] slv_r_user_o;
	input wire slv_r_ready_i;
	output reg slv_r_valid_o;
	output reg [1:0] slv_b_resp_o;
	output reg [AXI_ID_WIDTH - 1:0] slv_b_id_o;
	output reg [AXI_USER_WIDTH - 1:0] slv_b_user_o;
	input wire slv_b_ready_i;
	output reg slv_b_valid_o;
	output wire [AXI_ADDR_WIDTH - 1:0] mst_aw_addr_o;
	output wire [2:0] mst_aw_prot_o;
	output wire [3:0] mst_aw_region_o;
	output wire [5:0] mst_aw_atop_o;
	output wire [7:0] mst_aw_len_o;
	output wire [2:0] mst_aw_size_o;
	output wire [1:0] mst_aw_burst_o;
	output wire mst_aw_lock_o;
	output wire [3:0] mst_aw_cache_o;
	output wire [3:0] mst_aw_qos_o;
	output wire [AXI_ID_WIDTH - 1:0] mst_aw_id_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_aw_user_o;
	input wire mst_aw_ready_i;
	output reg mst_aw_valid_o;
	output wire [AXI_ADDR_WIDTH - 1:0] mst_ar_addr_o;
	output wire [2:0] mst_ar_prot_o;
	output wire [3:0] mst_ar_region_o;
	output wire [7:0] mst_ar_len_o;
	output wire [2:0] mst_ar_size_o;
	output wire [1:0] mst_ar_burst_o;
	output wire mst_ar_lock_o;
	output wire [3:0] mst_ar_cache_o;
	output wire [3:0] mst_ar_qos_o;
	output wire [AXI_ID_WIDTH - 1:0] mst_ar_id_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_ar_user_o;
	input wire mst_ar_ready_i;
	output reg mst_ar_valid_o;
	output wire [AXI_DATA_WIDTH - 1:0] mst_w_data_o;
	output wire [AXI_STRB_WIDTH - 1:0] mst_w_strb_o;
	output wire [AXI_USER_WIDTH - 1:0] mst_w_user_o;
	output wire mst_w_last_o;
	input wire mst_w_ready_i;
	output reg mst_w_valid_o;
	input wire [AXI_DATA_WIDTH - 1:0] mst_r_data_i;
	input wire [1:0] mst_r_resp_i;
	input wire mst_r_last_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_r_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_r_user_i;
	output reg mst_r_ready_o;
	input wire mst_r_valid_i;
	input wire [1:0] mst_b_resp_i;
	input wire [AXI_ID_WIDTH - 1:0] mst_b_id_i;
	input wire [AXI_USER_WIDTH - 1:0] mst_b_user_i;
	output reg mst_b_ready_o;
	input wire mst_b_valid_i;
	reg [AXI_ID_WIDTH - 1:0] art_check_id;
	reg [AXI_ID_WIDTH - 1:0] art_set_id;
	reg [AXI_ID_WIDTH - 1:0] w_id_d;
	reg [AXI_ID_WIDTH - 1:0] w_id_q;
	reg [AXI_ADDR_WIDTH - 1:0] art_check_addr;
	wire [AXI_ADDR_WIDTH - 1:0] art_clr_addr;
	reg [AXI_ADDR_WIDTH - 1:0] art_set_addr;
	reg [AXI_ADDR_WIDTH - 1:0] rd_clr_addr;
	reg [AXI_ADDR_WIDTH - 1:0] wr_clr_addr;
	reg [AXI_ADDR_WIDTH - 1:0] w_addr_d;
	reg [AXI_ADDR_WIDTH - 1:0] w_addr_q;
	reg art_check_req;
	wire art_check_gnt;
	wire art_clr_req;
	wire art_clr_gnt;
	reg art_set_req;
	wire art_set_gnt;
	reg rd_clr_req;
	wire rd_clr_gnt;
	reg wr_clr_req;
	wire wr_clr_gnt;
	wire art_check_res;
	reg b_excl_d;
	reg b_excl_q;
	reg r_excl_d;
	reg r_excl_q;
	reg [1:0] r_state_d;
	reg [1:0] r_state_q;
	reg [2:0] w_state_d;
	reg [2:0] w_state_q;
	assign mst_ar_addr_o = slv_ar_addr_i;
	assign mst_ar_prot_o = slv_ar_prot_i;
	assign mst_ar_region_o = slv_ar_region_i;
	assign mst_ar_len_o = slv_ar_len_i;
	assign mst_ar_size_o = slv_ar_size_i;
	assign mst_ar_burst_o = slv_ar_burst_i;
	assign mst_ar_lock_o = 1'b0;
	assign mst_ar_cache_o = slv_ar_cache_i;
	assign mst_ar_qos_o = slv_ar_qos_i;
	assign mst_ar_id_o = slv_ar_id_i;
	assign mst_ar_user_o = slv_ar_user_i;
	assign slv_r_data_o = mst_r_data_i;
	assign slv_r_last_o = mst_r_last_i;
	assign slv_r_id_o = mst_r_id_i;
	assign slv_r_user_o = mst_r_user_i;
	always @(*) begin
		mst_ar_valid_o = 1'b0;
		slv_ar_ready_o = 1'b0;
		mst_r_ready_o = 1'b0;
		slv_r_valid_o = 1'b0;
		slv_r_resp_o = 1'sb0;
		art_set_addr = 1'sb0;
		art_set_id = 1'sb0;
		art_set_req = 1'b0;
		rd_clr_addr = 1'sb0;
		rd_clr_req = 1'b0;
		r_excl_d = r_excl_q;
		r_state_d = r_state_q;
		case (r_state_q)
			2'd0:
				if (slv_ar_valid_i) begin
					if ((((slv_ar_addr_i >= ADDR_BEGIN) && (slv_ar_addr_i <= ADDR_END)) && slv_ar_lock_i) && (slv_ar_len_i == 8'h00)) begin
						art_set_addr = slv_ar_addr_i;
						art_set_id = slv_ar_id_i;
						art_set_req = 1'b1;
						r_excl_d = 1'b1;
						if (art_set_gnt) begin
							mst_ar_valid_o = 1'b1;
							if (mst_ar_ready_i) begin
								slv_ar_ready_o = 1'b1;
								r_state_d = 2'd2;
							end
							else
								r_state_d = 2'd1;
						end
					end
					else begin
						r_excl_d = 1'b0;
						mst_ar_valid_o = 1'b1;
						if (mst_ar_ready_i) begin
							slv_ar_ready_o = 1'b1;
							r_state_d = 2'd2;
						end
						else
							r_state_d = 2'd1;
					end
				end
			2'd1: begin
				mst_ar_valid_o = slv_ar_valid_i;
				slv_ar_ready_o = mst_ar_ready_i;
				if (mst_ar_ready_i && mst_ar_valid_o)
					r_state_d = 2'd2;
			end
			2'd2: begin
				mst_r_ready_o = slv_r_ready_i;
				slv_r_valid_o = mst_r_valid_i;
				if (mst_r_resp_i[1] == 1'b0)
					slv_r_resp_o = {1'b0, r_excl_q};
				else
					slv_r_resp_o = mst_r_resp_i;
				if ((mst_r_valid_i && mst_r_ready_o) && mst_r_last_i) begin
					r_excl_d = 1'b0;
					r_state_d = 2'd0;
				end
			end
			default: r_state_d = 2'd0;
		endcase
	end
	assign mst_aw_addr_o = slv_aw_addr_i;
	assign mst_aw_prot_o = slv_aw_prot_i;
	assign mst_aw_region_o = slv_aw_region_i;
	assign mst_aw_atop_o = slv_aw_atop_i;
	assign mst_aw_len_o = slv_aw_len_i;
	assign mst_aw_size_o = slv_aw_size_i;
	assign mst_aw_burst_o = slv_aw_burst_i;
	assign mst_aw_lock_o = 1'b0;
	assign mst_aw_cache_o = slv_aw_cache_i;
	assign mst_aw_qos_o = slv_aw_qos_i;
	assign mst_aw_id_o = slv_aw_id_i;
	assign mst_aw_user_o = slv_aw_user_i;
	assign mst_w_data_o = slv_w_data_i;
	assign mst_w_strb_o = slv_w_strb_i;
	assign mst_w_user_o = slv_w_user_i;
	assign mst_w_last_o = slv_w_last_i;
	always @(*) begin
		w_addr_d = w_addr_q;
		w_id_d = w_id_q;
		if (slv_aw_valid_i && slv_aw_ready_o) begin
			w_addr_d = slv_aw_addr_i;
			w_id_d = slv_aw_id_i;
		end
	end
	always @(*) begin
		mst_aw_valid_o = 1'b0;
		slv_aw_ready_o = 1'b0;
		mst_w_valid_o = 1'b0;
		slv_w_ready_o = 1'b0;
		slv_b_valid_o = 1'b0;
		mst_b_ready_o = 1'b0;
		slv_b_resp_o = 1'sb0;
		slv_b_id_o = 1'sb0;
		slv_b_user_o = 1'sb0;
		art_check_addr = 1'sb0;
		art_check_id = 1'sb0;
		art_check_req = 1'b0;
		wr_clr_addr = 1'sb0;
		wr_clr_req = 1'b0;
		b_excl_d = b_excl_q;
		w_state_d = w_state_q;
		case (w_state_q)
			3'd0:
				if (slv_aw_valid_i) begin
					if ((slv_aw_addr_i >= ADDR_BEGIN) && (slv_aw_addr_i <= ADDR_END)) begin
						if (slv_aw_lock_i && (slv_aw_len_i == 8'h00)) begin
							art_check_addr = slv_aw_addr_i;
							art_check_id = slv_aw_id_i;
							art_check_req = 1'b1;
							if (art_check_gnt) begin
								if (art_check_res) begin
									mst_aw_valid_o = 1'b1;
									if (mst_aw_ready_i) begin
										slv_aw_ready_o = 1'b1;
										b_excl_d = 1'b1;
										w_state_d = 3'd1;
									end
								end
								else begin
									slv_aw_ready_o = 1'b1;
									w_state_d = 3'd4;
								end
							end
						end
						else begin
							mst_aw_valid_o = 1'b1;
							if (mst_aw_ready_i) begin
								slv_aw_ready_o = 1'b1;
								w_state_d = 3'd1;
							end
						end
					end
					else begin
						mst_aw_valid_o = 1'b1;
						slv_aw_ready_o = mst_aw_ready_i;
						if (slv_aw_ready_o)
							w_state_d = 3'd2;
					end
				end
			3'd1: begin
				mst_w_valid_o = slv_w_valid_i;
				slv_w_ready_o = mst_w_ready_i;
				if ((slv_w_valid_i && slv_w_ready_o) && slv_w_last_i) begin
					wr_clr_addr = w_addr_q;
					wr_clr_req = 1'b1;
					if (wr_clr_gnt)
						w_state_d = 3'd5;
					else
						w_state_d = 3'd3;
				end
			end
			3'd2: begin
				mst_w_valid_o = slv_w_valid_i;
				slv_w_ready_o = mst_w_ready_i;
				if ((slv_w_valid_i && slv_w_ready_o) && slv_w_last_i)
					w_state_d = 3'd5;
			end
			3'd3: begin
				wr_clr_addr = w_addr_q;
				wr_clr_req = 1'b1;
				if (wr_clr_gnt)
					w_state_d = 3'd5;
			end
			3'd4: begin
				slv_w_ready_o = 1'b1;
				if (slv_w_valid_i && slv_w_last_i)
					w_state_d = 3'd6;
			end
			3'd5: begin
				mst_b_ready_o = slv_b_ready_i;
				slv_b_valid_o = mst_b_valid_i;
				slv_b_resp_o[1] = mst_b_resp_i[1];
				slv_b_resp_o[0] = (mst_b_resp_i[1] == 1'b0 ? b_excl_q : mst_b_resp_i[0]);
				slv_b_user_o = mst_b_user_i;
				slv_b_id_o = mst_b_id_i;
				if (slv_b_valid_o && slv_b_ready_i) begin
					b_excl_d = 1'b0;
					w_state_d = 3'd0;
				end
			end
			3'd6: begin
				slv_b_id_o = w_id_q;
				slv_b_resp_o = 2'b00;
				slv_b_valid_o = 1'b1;
				if (slv_b_ready_i)
					w_state_d = 3'd0;
			end
			default: w_state_d = 3'd0;
		endcase
	end
	axi_res_tbl #(
		.AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
		.AXI_ID_WIDTH(AXI_ID_WIDTH)
	) i_art(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.clr_addr_i(art_clr_addr),
		.clr_req_i(art_clr_req),
		.clr_gnt_o(art_clr_gnt),
		.set_addr_i(art_set_addr),
		.set_id_i(art_set_id),
		.set_req_i(art_set_req),
		.set_gnt_o(art_set_gnt),
		.check_addr_i(art_check_addr),
		.check_id_i(art_check_id),
		.check_res_o(art_check_res),
		.check_req_i(art_check_req),
		.check_gnt_o(art_check_gnt)
	);
	stream_arbiter_22976_4AFBD #(
		.DATA_T_AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
		.N_INP(2)
	) i_non_excl_acc_arb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.inp_data_i({rd_clr_addr, wr_clr_addr}),
		.inp_valid_i({rd_clr_req, wr_clr_req}),
		.inp_ready_o({rd_clr_gnt, wr_clr_gnt}),
		.oup_data_o(art_clr_addr),
		.oup_valid_o(art_clr_req),
		.oup_ready_i(art_clr_gnt)
	);
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			b_excl_q <= 1'b0;
			r_excl_q <= 1'b0;
			r_state_q <= 2'd0;
			w_addr_q <= 1'sb0;
			w_id_q <= 1'sb0;
			w_state_q <= 3'd0;
		end
		else begin
			b_excl_q <= b_excl_d;
			r_excl_q <= r_excl_d;
			r_state_q <= r_state_d;
			w_addr_q <= w_addr_d;
			w_id_q <= w_id_d;
			w_state_q <= w_state_d;
		end
endmodule
module exp_backoff (
	clk_i,
	rst_ni,
	set_i,
	clr_i,
	is_zero_o
);
	parameter [31:0] Seed = 'hffff;
	parameter [31:0] MaxExp = 16;
	input wire clk_i;
	input wire rst_ni;
	input wire set_i;
	input wire clr_i;
	output wire is_zero_o;
	localparam WIDTH = 16;
	wire [15:0] lfsr_d;
	reg [15:0] lfsr_q;
	wire [15:0] cnt_d;
	reg [15:0] cnt_q;
	wire [15:0] mask_d;
	reg [15:0] mask_q;
	wire lfsr;
	assign lfsr = ((lfsr_q[0] ^ lfsr_q[2]) ^ lfsr_q[3]) ^ lfsr_q[5];
	assign lfsr_d = (set_i ? {lfsr, lfsr_q[15:1]} : lfsr_q);
	assign mask_d = (clr_i ? {16 {1'sb0}} : (set_i ? {{WIDTH - MaxExp {1'b0}}, mask_q[MaxExp - 2:0], 1'b1} : mask_q));
	assign cnt_d = (clr_i ? {16 {1'sb0}} : (set_i ? mask_q & lfsr_q : (!is_zero_o ? cnt_q - 1'b1 : {16 {1'sb0}})));
	assign is_zero_o = cnt_q == {16 {1'sb0}};
	function automatic [15:0] sv2v_cast_16;
		input reg [15:0] inp;
		sv2v_cast_16 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni) begin : p_regs
		if (!rst_ni) begin
			lfsr_q <= sv2v_cast_16(Seed);
			mask_q <= 1'sb0;
			cnt_q <= 1'sb0;
		end
		else begin
			lfsr_q <= lfsr_d;
			mask_q <= mask_d;
			cnt_q <= cnt_d;
		end
	end
endmodule
module sram (
	clk_i,
	rst_ni,
	req_i,
	we_i,
	addr_i,
	wdata_i,
	be_i,
	rdata_o
);
	parameter DATA_WIDTH = 64;
	parameter NUM_WORDS = 1024;
	parameter OUT_REGS = 0;
	parameter DROMAJO_RAM = 0;
	input wire clk_i;
	input wire rst_ni;
	input wire req_i;
	input wire we_i;
	input wire [$clog2(NUM_WORDS) - 1:0] addr_i;
	input wire [DATA_WIDTH - 1:0] wdata_i;
	input wire [((DATA_WIDTH + 7) / 8) - 1:0] be_i;
	output reg [DATA_WIDTH - 1:0] rdata_o;
	localparam DATA_WIDTH_ALIGNED = ((DATA_WIDTH + 63) / 64) * 64;
	localparam BE_WIDTH_ALIGNED = ((((DATA_WIDTH + 7) / 8) + 7) / 8) * 8;
	reg [DATA_WIDTH_ALIGNED - 1:0] wdata_aligned;
	reg [BE_WIDTH_ALIGNED - 1:0] be_aligned;
	wire [DATA_WIDTH_ALIGNED - 1:0] rdata_aligned;
	always @(*) begin : p_align
		wdata_aligned = 1'sb0;
		be_aligned = 1'sb0;
		wdata_aligned[DATA_WIDTH - 1:0] = wdata_i;
		be_aligned[BE_WIDTH_ALIGNED - 1:0] = be_i;
		rdata_o = rdata_aligned[DATA_WIDTH - 1:0];
	end
	genvar k;
	generate
		for (k = 0; k < ((DATA_WIDTH + 63) / 64); k = k + 1) begin : gen_cut
			if (DROMAJO_RAM) begin : gen_dromajo
				dromajo_ram #(
					.ADDR_WIDTH($clog2(NUM_WORDS)),
					.DATA_DEPTH(NUM_WORDS),
					.OUT_REGS(0)
				) i_ram(
					.Clk_CI(clk_i),
					.Rst_RBI(rst_ni),
					.CSel_SI(req_i),
					.WrEn_SI(we_i),
					.BEn_SI(be_aligned[k * 8+:8]),
					.WrData_DI(wdata_aligned[k * 64+:64]),
					.Addr_DI(addr_i),
					.RdData_DO(rdata_aligned[k * 64+:64])
				);
			end
			else begin : gen_mem
				SyncSpRamBeNx64 #(
					.ADDR_WIDTH($clog2(NUM_WORDS)),
					.DATA_DEPTH(NUM_WORDS),
					.OUT_REGS(0),
					.SIM_INIT(1)
				) i_ram(
					.Clk_CI(clk_i),
					.Rst_RBI(rst_ni),
					.CSel_SI(req_i),
					.WrEn_SI(we_i),
					.BEn_SI(be_aligned[k * 8+:8]),
					.WrData_DI(wdata_aligned[k * 64+:64]),
					.Addr_DI(addr_i),
					.RdData_DO(rdata_aligned[k * 64+:64])
				);
			end
		end
	endgenerate
endmodule
module SyncSpRamBeNx64 (
	Clk_CI,
	Rst_RBI,
	CSel_SI,
	WrEn_SI,
	BEn_SI,
	WrData_DI,
	Addr_DI,
	RdData_DO
);
	parameter ADDR_WIDTH = 10;
	parameter DATA_DEPTH = 1024;
	parameter OUT_REGS = 0;
	parameter SIM_INIT = 0;
	input wire Clk_CI;
	input wire Rst_RBI;
	input wire CSel_SI;
	input wire WrEn_SI;
	input wire [7:0] BEn_SI;
	input wire [63:0] WrData_DI;
	input wire [ADDR_WIDTH - 1:0] Addr_DI;
	output wire [63:0] RdData_DO;
	localparam DATA_BYTES = 8;
	reg [63:0] RdData_DN;
	reg [63:0] RdData_DP;
	reg [63:0] Mem_DP [DATA_DEPTH - 1:0];
	always @(posedge Clk_CI) begin : sv2v_autoblock_1
		reg [63:0] val;
		if ((Rst_RBI == 1'b0) && (SIM_INIT > 0)) begin : sv2v_autoblock_2
			reg signed [31:0] k;
			for (k = 0; k < DATA_DEPTH; k = k + 1)
				begin
					if (SIM_INIT == 1)
						val = 1'sb0;
					else
						val = 64'hdeadbeefdeadbeef;
					Mem_DP[k] = val;
				end
		end
		else if (CSel_SI) begin
			if (WrEn_SI) begin
				if (BEn_SI[0])
					Mem_DP[Addr_DI][7:0] <= WrData_DI[7:0];
				if (BEn_SI[1])
					Mem_DP[Addr_DI][15:8] <= WrData_DI[15:8];
				if (BEn_SI[2])
					Mem_DP[Addr_DI][23:16] <= WrData_DI[23:16];
				if (BEn_SI[3])
					Mem_DP[Addr_DI][31:24] <= WrData_DI[31:24];
				if (BEn_SI[4])
					Mem_DP[Addr_DI][39:32] <= WrData_DI[39:32];
				if (BEn_SI[5])
					Mem_DP[Addr_DI][47:40] <= WrData_DI[47:40];
				if (BEn_SI[6])
					Mem_DP[Addr_DI][55:48] <= WrData_DI[55:48];
				if (BEn_SI[7])
					Mem_DP[Addr_DI][63:56] <= WrData_DI[63:56];
			end
			RdData_DN <= Mem_DP[Addr_DI];
		end
	end
	generate
		if (OUT_REGS > 0) begin : g_outreg
			always @(posedge Clk_CI or negedge Rst_RBI)
				if (Rst_RBI == 1'b0)
					RdData_DP <= 0;
				else
					RdData_DP <= RdData_DN;
		end
		if (OUT_REGS == 0) begin : g_oureg_byp
			wire [64:1] sv2v_tmp_7FD8C;
			assign sv2v_tmp_7FD8C = RdData_DN;
			always @(*) RdData_DP = sv2v_tmp_7FD8C;
		end
	endgenerate
	assign RdData_DO = RdData_DP;
endmodule
module unread (d_i);
	input wire d_i;
endmodule
module stream_arbiter_22976_4AFBD (
	clk_i,
	rst_ni,
	inp_data_i,
	inp_valid_i,
	inp_ready_o,
	oup_data_o,
	oup_valid_o,
	oup_ready_i
);
	parameter [31:0] DATA_T_AXI_ADDR_WIDTH = 0;
	parameter integer N_INP = -1;
	parameter ARBITER = "rr";
	input wire clk_i;
	input wire rst_ni;
	input wire [(N_INP * DATA_T_AXI_ADDR_WIDTH) - 1:0] inp_data_i;
	input wire [N_INP - 1:0] inp_valid_i;
	output wire [N_INP - 1:0] inp_ready_o;
	output wire [DATA_T_AXI_ADDR_WIDTH - 1:0] oup_data_o;
	output wire oup_valid_o;
	input wire oup_ready_i;
	stream_arbiter_flushable_2A141_DBD2E #(
		.DATA_T_DATA_T_AXI_ADDR_WIDTH(DATA_T_AXI_ADDR_WIDTH),
		.N_INP(N_INP),
		.ARBITER(ARBITER)
	) i_arb(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.flush_i(1'b0),
		.inp_data_i(inp_data_i),
		.inp_valid_i(inp_valid_i),
		.inp_ready_o(inp_ready_o),
		.oup_data_o(oup_data_o),
		.oup_valid_o(oup_valid_o),
		.oup_ready_i(oup_ready_i)
	);
endmodule
module stream_arbiter_flushable_2A141_DBD2E (
	clk_i,
	rst_ni,
	flush_i,
	inp_data_i,
	inp_valid_i,
	inp_ready_o,
	oup_data_o,
	oup_valid_o,
	oup_ready_i
);
	parameter [31:0] DATA_T_DATA_T_AXI_ADDR_WIDTH = 0;
	parameter integer N_INP = -1;
	parameter ARBITER = "rr";
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [(N_INP * DATA_T_DATA_T_AXI_ADDR_WIDTH) - 1:0] inp_data_i;
	input wire [N_INP - 1:0] inp_valid_i;
	output wire [N_INP - 1:0] inp_ready_o;
	output wire [DATA_T_DATA_T_AXI_ADDR_WIDTH - 1:0] oup_data_o;
	output wire oup_valid_o;
	input wire oup_ready_i;
	generate
		if (ARBITER == "rr") begin : gen_rr_arb
			localparam [31:0] sv2v_uu_i_arbiter_NumIn = N_INP;
			localparam [$clog2(sv2v_uu_i_arbiter_NumIn) - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_E10E8_57195 #(
				.DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH(DATA_T_DATA_T_AXI_ADDR_WIDTH),
				.NumIn(N_INP),
				.ExtPrio(1'b0),
				.AxiVldRdy(1'b1),
				.LockIn(1'b1)
			) i_arbiter(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
				.req_i(inp_valid_i),
				.gnt_o(inp_ready_o),
				.data_i(inp_data_i),
				.gnt_i(oup_ready_i),
				.req_o(oup_valid_o),
				.data_o(oup_data_o),
				.idx_o()
			);
		end
		else if (ARBITER == "prio") begin : gen_prio_arb
			localparam [31:0] sv2v_uu_i_arbiter_NumIn = N_INP;
			localparam [$clog2(sv2v_uu_i_arbiter_NumIn) - 1:0] sv2v_uu_i_arbiter_ext_rr_i_0 = 1'sb0;
			rr_arb_tree_E10E8_57195 #(
				.DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH(DATA_T_DATA_T_AXI_ADDR_WIDTH),
				.NumIn(N_INP),
				.ExtPrio(1'b1),
				.AxiVldRdy(1'b1),
				.LockIn(1'b1)
			) i_arbiter(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(flush_i),
				.rr_i(sv2v_uu_i_arbiter_ext_rr_i_0),
				.req_i(inp_valid_i),
				.gnt_o(inp_ready_o),
				.data_i(inp_data_i),
				.gnt_i(oup_ready_i),
				.req_o(oup_valid_o),
				.data_o(oup_data_o),
				.idx_o()
			);
		end
		// else begin : gen_arb_error
		// 	$fatal(1, "Invalid value for parameter 'ARBITER'!");
		// end
	endgenerate
endmodule
module fifo_v3 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [DATA_WIDTH - 1:0] data_i;
	input wire push_i;
	output reg [DATA_WIDTH - 1:0] data_o;
	input wire pop_i;
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [(FIFO_DEPTH * DATA_WIDTH) - 1:0] mem_n;
	reg [(FIFO_DEPTH * DATA_WIDTH) - 1:0] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : genblk1
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : genblk1
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * DATA_WIDTH+:DATA_WIDTH]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[write_pointer_q * DATA_WIDTH+:DATA_WIDTH] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= 1'sb0;
		else if (!gate_clock)
			mem_q <= mem_n;
endmodule
module fifo_v3_4F30F_AEF03 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter signed [31:0] dtype_riscv_PLEN = 0;
	parameter signed [31:0] dtype_riscv_XLEN = 0;
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1:0] data_i;
	input wire push_i;
	output reg [((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1:0] data_o;
	input wire pop_i;
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? (FIFO_DEPTH * (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2)) - 1 : (FIFO_DEPTH * (1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1))) + (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 0)):((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? 0 : ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1)] mem_n;
	reg [((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? (FIFO_DEPTH * (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2)) - 1 : (FIFO_DEPTH * (1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1))) + (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 0)):((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? 0 : ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1)] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : genblk1
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : genblk1
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? 0 : ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) + (read_pointer_q * ((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2 : 1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1)))+:((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2 : 1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1))]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? 0 : ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) + (write_pointer_q * ((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2 : 1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1)))+:((((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1) >= 0 ? ((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 2 : 1 - (((4 + dtype_riscv_PLEN) + dtype_riscv_XLEN) + 1))] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= 1'sb0;
		else if (!gate_clock)
			mem_q <= mem_n;
endmodule
module fifo_v3_6C4C9_25B33 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter signed [31:0] dtype_i_icache_data_fifo_sv2v_pfunc_651B1 = 0;
	parameter signed [31:0] dtype_riscv_PLEN = 0;
	parameter signed [31:0] dtype_wt_cache_pkg_CACHE_ID_WIDTH = 0;
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [(((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) - 1:0] data_i;
	input wire push_i;
	output reg [(((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) - 1:0] data_o;
	input wire pop_i;
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [(FIFO_DEPTH * (((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH)) - 1:0] mem_n;
	reg [(FIFO_DEPTH * (((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH)) - 1:0] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : genblk1
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : genblk1
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * (((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH)+:((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[write_pointer_q * (((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH)+:((dtype_i_icache_data_fifo_sv2v_pfunc_651B1 + dtype_riscv_PLEN) + 1) + dtype_wt_cache_pkg_CACHE_ID_WIDTH] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= 1'sb0;
		else if (!gate_clock)
			mem_q <= mem_n;
endmodule
module fifo_v3_77734_A8EA3 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter signed [31:0] dtype_riscv_PLEN = 0;
	parameter signed [31:0] dtype_wt_cache_pkg_CACHE_ID_WIDTH = 0;
	parameter integer dtype_wt_cache_pkg_L1D_WAY_WIDTH = 0;
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3:0] data_i;
	input wire push_i;
	output reg [((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3:0] data_o;
	input wire pop_i;
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? (FIFO_DEPTH * (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4)) - 1 : (FIFO_DEPTH * (1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3))) + (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 2)):((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? 0 : ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3)] mem_n;
	reg [((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? (FIFO_DEPTH * (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4)) - 1 : (FIFO_DEPTH * (1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3))) + (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 2)):((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? 0 : ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3)] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : genblk1
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : genblk1
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? 0 : ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) + (read_pointer_q * ((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4 : 1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3)))+:((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4 : 1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3))]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? 0 : ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) + (write_pointer_q * ((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4 : 1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3)))+:((((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3) >= 0 ? ((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 4 : 1 - (((((5 + dtype_wt_cache_pkg_L1D_WAY_WIDTH) + dtype_riscv_PLEN) + 65) + dtype_wt_cache_pkg_CACHE_ID_WIDTH) + 3))] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= 1'sb0;
		else if (!gate_clock)
			mem_q <= mem_n;
endmodule
module fifo_v3_AECA2_3F763 (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter signed [31:0] dtype_riscv_VLEN = 0;
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [(37 + dtype_riscv_VLEN) - 1:0] data_i;
	input wire push_i;
	output reg [(37 + dtype_riscv_VLEN) - 1:0] data_o;
	input wire pop_i;
	localparam [31:0] FIFO_DEPTH = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [(FIFO_DEPTH * (37 + dtype_riscv_VLEN)) - 1:0] mem_n;
	reg [(FIFO_DEPTH * (37 + dtype_riscv_VLEN)) - 1:0] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : genblk1
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : genblk1
			assign full_o = status_cnt_q == FIFO_DEPTH[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[read_pointer_q * (37 + dtype_riscv_VLEN)+:37 + dtype_riscv_VLEN]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[write_pointer_q * (37 + dtype_riscv_VLEN)+:37 + dtype_riscv_VLEN] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FIFO_DEPTH[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= 1'sb0;
		else if (!gate_clock)
			mem_q <= mem_n;
endmodule
module lzc (
	in_i,
	cnt_o,
	empty_o
);
	parameter [31:0] WIDTH = 2;
	parameter [0:0] MODE = 1'b0;
	parameter [31:0] CNT_WIDTH = (WIDTH == 1 ? 1 : $clog2(WIDTH));
	input wire [WIDTH - 1:0] in_i;
	output wire [CNT_WIDTH - 1:0] cnt_o;
	output wire empty_o;
	generate
		if (WIDTH == 1) begin : gen_degenerate_lzc
			assign cnt_o[0] = !in_i[0];
			assign empty_o = !in_i[0];
		end
		else begin : gen_lzc
			localparam [31:0] NUM_LEVELS = $clog2(WIDTH);
			wire [(WIDTH * NUM_LEVELS) - 1:0] index_lut;
			wire [(2 ** NUM_LEVELS) - 1:0] sel_nodes;
			wire [((2 ** NUM_LEVELS) * NUM_LEVELS) - 1:0] index_nodes;
			reg [WIDTH - 1:0] in_tmp;
			always @(*) begin : flip_vector
				begin : sv2v_autoblock_1
					reg [31:0] i;
					for (i = 0; i < WIDTH; i = i + 1)
						in_tmp[i] = (MODE ? in_i[(WIDTH - 1) - i] : in_i[i]);
				end
			end
			genvar j;
			for (j = 0; $unsigned(j) < WIDTH; j = j + 1) begin : g_index_lut
				function automatic [NUM_LEVELS - 1:0] sv2v_cast_7179C;
					input reg [NUM_LEVELS - 1:0] inp;
					sv2v_cast_7179C = inp;
				endfunction
				assign index_lut[j * NUM_LEVELS+:NUM_LEVELS] = sv2v_cast_7179C($unsigned(j));
			end
			genvar level;
			for (level = 0; $unsigned(level) < NUM_LEVELS; level = level + 1) begin : g_levels
				if ($unsigned(level) == (NUM_LEVELS - 1)) begin : g_last_level
					genvar k;
					for (k = 0; k < (2 ** level); k = k + 1) begin : g_level
						if (($unsigned(k) * 2) < (WIDTH - 1)) begin : genblk1
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2] | in_tmp[(k * 2) + 1];
							assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = (in_tmp[k * 2] == 1'b1 ? index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS] : index_lut[((k * 2) + 1) * NUM_LEVELS+:NUM_LEVELS]);
						end
						if (($unsigned(k) * 2) == (WIDTH - 1)) begin : genblk2
							assign sel_nodes[((2 ** level) - 1) + k] = in_tmp[k * 2];
							assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = index_lut[(k * 2) * NUM_LEVELS+:NUM_LEVELS];
						end
						if (($unsigned(k) * 2) > (WIDTH - 1)) begin : genblk3
							assign sel_nodes[((2 ** level) - 1) + k] = 1'b0;
							assign index_nodes[(((2 ** level) - 1) + k) * NUM_LEVELS+:NUM_LEVELS] = 1'sb0;
						end
					end
				end
				else begin : genblk1
					genvar l;
					for (l = 0; l < (2 ** level); l = l + 1) begin : g_level
						assign sel_nodes[((2 ** level) - 1) + l] = sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] | sel_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) + 1];
						assign index_nodes[(((2 ** level) - 1) + l) * NUM_LEVELS+:NUM_LEVELS] = (sel_nodes[((2 ** (level + 1)) - 1) + (l * 2)] == 1'b1 ? index_nodes[(((2 ** (level + 1)) - 1) + (l * 2)) * NUM_LEVELS+:NUM_LEVELS] : index_nodes[((((2 ** (level + 1)) - 1) + (l * 2)) + 1) * NUM_LEVELS+:NUM_LEVELS]);
					end
				end
			end
			assign cnt_o = (NUM_LEVELS > $unsigned(0) ? index_nodes[0+:NUM_LEVELS] : {$clog2(WIDTH) {1'b0}});
			assign empty_o = (NUM_LEVELS > $unsigned(0) ? ~sel_nodes[0] : ~(|in_i));
		end
	endgenerate
endmodule
module popcount (
	data_i,
	popcount_o
);
	parameter [31:0] INPUT_WIDTH = 256;
	localparam POPCOUNT_WIDTH = $clog2(INPUT_WIDTH) + 1;
	input wire [INPUT_WIDTH - 1:0] data_i;
	output wire [POPCOUNT_WIDTH - 1:0] popcount_o;
	localparam [31:0] PADDED_WIDTH = 1 << $clog2(INPUT_WIDTH);
	reg [PADDED_WIDTH - 1:0] padded_input;
	wire [POPCOUNT_WIDTH - 2:0] left_child_result;
	wire [POPCOUNT_WIDTH - 2:0] right_child_result;
	always @(*) begin
		padded_input = 1'sb0;
		padded_input[INPUT_WIDTH - 1:0] = data_i;
	end
	generate
		if (INPUT_WIDTH == 1) begin : single_node
			assign left_child_result = 1'b0;
			assign right_child_result = padded_input[0];
		end
		else if (INPUT_WIDTH == 2) begin : leaf_node
			assign left_child_result = padded_input[1];
			assign right_child_result = padded_input[0];
		end
		else begin : non_leaf_node
			popcount #(.INPUT_WIDTH(PADDED_WIDTH / 2)) left_child(
				.data_i(padded_input[PADDED_WIDTH - 1:PADDED_WIDTH / 2]),
				.popcount_o(left_child_result)
			);
			popcount #(.INPUT_WIDTH(PADDED_WIDTH / 2)) right_child(
				.data_i(padded_input[(PADDED_WIDTH / 2) - 1:0]),
				.popcount_o(right_child_result)
			);
		end
	endgenerate
	assign popcount_o = left_child_result + right_child_result;
endmodule
module rr_arb_tree (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [(NumIn * DataWidth) - 1:0] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [DataWidth - 1:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	function automatic [DataWidth - 1:0] sv2v_cast_4AF59;
		input reg [DataWidth - 1:0] inp;
		sv2v_cast_4AF59 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[0+:DataWidth];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * DataWidth) - 1 : ((3 - (2 ** NumLevels)) * DataWidth) + ((((2 ** NumLevels) - 2) * DataWidth) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * DataWidth)] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * DataWidth+:DataWidth];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataWidth+:DataWidth] = (sel ? data_i[((l * 2) + 1) * DataWidth+:DataWidth] : data_i[(l * 2) * DataWidth+:DataWidth]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataWidth+:DataWidth] = data_i[(l * 2) * DataWidth+:DataWidth];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_4AF59(1'sb0);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataWidth+:DataWidth] = sv2v_cast_4AF59(1'sb0);
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataWidth+:DataWidth] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * DataWidth+:DataWidth] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * DataWidth+:DataWidth]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_866BD_14B99 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] DataType_ariane_pkg_DCACHE_INDEX_WIDTH = 0;
	parameter [31:0] DataType_ariane_pkg_DCACHE_SET_ASSOC = 0;
	parameter [31:0] DataType_ariane_pkg_DCACHE_TAG_WIDTH = 0;
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [(NumIn * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)) - 1:0] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [(((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC) - 1:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	function automatic [(((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC) - 1:0] sv2v_cast_ECD4F;
		input reg [(((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC) - 1:0] inp;
		sv2v_cast_ECD4F = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[0+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)) - 1 : ((3 - (2 ** NumLevels)) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)) + ((((2 ** NumLevels) - 2) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC))] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] = (sel ? data_i[((l * 2) + 1) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] : data_i[(l * 2) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] = data_i[(l * 2) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_ECD4F(1'sb0);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] = sv2v_cast_ECD4F(1'sb0);
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * (((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC)+:((DataType_ariane_pkg_DCACHE_INDEX_WIDTH + DataType_ariane_pkg_DCACHE_TAG_WIDTH) + 89) + DataType_ariane_pkg_DCACHE_SET_ASSOC]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_88014 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [(NumIn * 4) - 1:0] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [3:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[0+:4];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * 4) - 1 : ((3 - (2 ** NumLevels)) * 4) + ((((2 ** NumLevels) - 2) * 4) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * 4)] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * 4+:4];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * 4+:4] = (sel ? data_i[((l * 2) + 1) * 4+:4] : data_i[(l * 2) * 4+:4]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * 4+:4] = data_i[(l * 2) * 4+:4];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 4'b0000;
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * 4+:4] = 4'b0000;
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * 4+:4] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * 4+:4] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * 4+:4]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_36817_A990F (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] DataType_Width = 0;
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [((DataType_Width + 8) >= 0 ? (NumIn * (DataType_Width + 9)) - 1 : (NumIn * (1 - (DataType_Width + 8))) + (DataType_Width + 7)):((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8)] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [DataType_Width + 8:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	function automatic [((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)) - 1:0] sv2v_cast_A7B3D;
		input reg [((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)) - 1:0] inp;
		sv2v_cast_A7B3D = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + 0+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? ((DataType_Width + 8) >= 0 ? (((2 ** NumLevels) - 1) * (DataType_Width + 9)) - 1 : (((2 ** NumLevels) - 1) * (1 - (DataType_Width + 8))) + (DataType_Width + 7)) : ((DataType_Width + 8) >= 0 ? ((3 - (2 ** NumLevels)) * (DataType_Width + 9)) + ((((2 ** NumLevels) - 2) * (DataType_Width + 9)) - 1) : ((3 - (2 ** NumLevels)) * (1 - (DataType_Width + 8))) + (((DataType_Width + 8) + (((2 ** NumLevels) - 2) * (1 - (DataType_Width + 8)))) - 1))):(((2 ** NumLevels) - 2) >= 0 ? ((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) : ((DataType_Width + 8) >= 0 ? ((2 ** NumLevels) - 2) * (DataType_Width + 9) : (DataType_Width + 8) + (((2 ** NumLevels) - 2) * (1 - (DataType_Width + 8)))))] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] = (sel ? data_i[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + (((l * 2) + 1) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] : data_i[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((l * 2) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] = data_i[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((l * 2) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_A7B3D(1'sb0);
							assign data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] = sv2v_cast_A7B3D(1'sb0);
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] = (sel ? data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))] : data_nodes[((DataType_Width + 8) >= 0 ? 0 : DataType_Width + 8) + ((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * ((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8)))+:((DataType_Width + 8) >= 0 ? DataType_Width + 9 : 1 - (DataType_Width + 8))]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_E10E8_57195 (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH = 0;
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [(NumIn * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH) - 1:0] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH - 1:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	function automatic [DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH - 1:0] sv2v_cast_DD039;
		input reg [DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH - 1:0] inp;
		sv2v_cast_DD039 = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[0+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH) - 1 : ((3 - (2 ** NumLevels)) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH) + ((((2 ** NumLevels) - 2) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH)] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] = (sel ? data_i[((l * 2) + 1) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] : data_i[(l * 2) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] = data_i[(l * 2) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_DD039(1'sb0);
							assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] = sv2v_cast_DD039(1'sb0);
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] = (sel ? data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH] : data_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH+:DataType_DATA_T_DATA_T_AXI_ADDR_WIDTH]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module rr_arb_tree_79FBE_62ECB (
	clk_i,
	rst_ni,
	flush_i,
	rr_i,
	req_i,
	gnt_o,
	data_i,
	gnt_i,
	req_o,
	data_o,
	idx_o
);
	parameter [31:0] DataType_WIDTH = 0;
	parameter [31:0] NumIn = 64;
	parameter [31:0] DataWidth = 32;
	parameter [0:0] ExtPrio = 1'b0;
	parameter [0:0] AxiVldRdy = 1'b0;
	parameter [0:0] LockIn = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire [$clog2(NumIn) - 1:0] rr_i;
	input wire [NumIn - 1:0] req_i;
	output wire [NumIn - 1:0] gnt_o;
	input wire [((DataType_WIDTH + 7) >= 0 ? (NumIn * (DataType_WIDTH + 8)) - 1 : (NumIn * (1 - (DataType_WIDTH + 7))) + (DataType_WIDTH + 6)):((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7)] data_i;
	input wire gnt_i;
	output wire req_o;
	output wire [DataType_WIDTH + 7:0] data_o;
	output wire [$clog2(NumIn) - 1:0] idx_o;
	function automatic [((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)) - 1:0] sv2v_cast_BB0BC;
		input reg [((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)) - 1:0] inp;
		sv2v_cast_BB0BC = inp;
	endfunction
	generate
		if (NumIn == $unsigned(1)) begin : genblk1
			assign req_o = req_i[0];
			assign gnt_o[0] = gnt_i;
			assign data_o = data_i[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + 0+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))];
			assign idx_o = 1'sb0;
		end
		else begin : genblk1
			localparam [31:0] NumLevels = $clog2(NumIn);
			wire [(((2 ** NumLevels) - 2) >= 0 ? (((2 ** NumLevels) - 1) * NumLevels) - 1 : ((3 - (2 ** NumLevels)) * NumLevels) + ((((2 ** NumLevels) - 2) * NumLevels) - 1)):(((2 ** NumLevels) - 2) >= 0 ? 0 : ((2 ** NumLevels) - 2) * NumLevels)] index_nodes;
			wire [(((2 ** NumLevels) - 2) >= 0 ? ((DataType_WIDTH + 7) >= 0 ? (((2 ** NumLevels) - 1) * (DataType_WIDTH + 8)) - 1 : (((2 ** NumLevels) - 1) * (1 - (DataType_WIDTH + 7))) + (DataType_WIDTH + 6)) : ((DataType_WIDTH + 7) >= 0 ? ((3 - (2 ** NumLevels)) * (DataType_WIDTH + 8)) + ((((2 ** NumLevels) - 2) * (DataType_WIDTH + 8)) - 1) : ((3 - (2 ** NumLevels)) * (1 - (DataType_WIDTH + 7))) + (((DataType_WIDTH + 7) + (((2 ** NumLevels) - 2) * (1 - (DataType_WIDTH + 7)))) - 1))):(((2 ** NumLevels) - 2) >= 0 ? ((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) : ((DataType_WIDTH + 7) >= 0 ? ((2 ** NumLevels) - 2) * (DataType_WIDTH + 8) : (DataType_WIDTH + 7) + (((2 ** NumLevels) - 2) * (1 - (DataType_WIDTH + 7)))))] data_nodes;
			wire [(2 ** NumLevels) - 2:0] gnt_nodes;
			wire [(2 ** NumLevels) - 2:0] req_nodes;
			reg [NumLevels - 1:0] rr_q;
			wire [NumIn - 1:0] req_d;
			assign req_o = req_nodes[0];
			assign data_o = data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))];
			assign idx_o = index_nodes[(((2 ** NumLevels) - 2) >= 0 ? 0 : (2 ** NumLevels) - 2) * NumLevels+:NumLevels];
			if (ExtPrio) begin : gen_ext_rr
				wire [NumLevels:1] sv2v_tmp_4C2F0;
				assign sv2v_tmp_4C2F0 = rr_i;
				always @(*) rr_q = sv2v_tmp_4C2F0;
				assign req_d = req_i;
			end
			else begin : gen_int_rr
				wire [NumLevels - 1:0] rr_d;
				if (LockIn) begin : gen_lock
					wire lock_d;
					reg lock_q;
					reg [NumIn - 1:0] req_q;
					assign lock_d = req_o & ~gnt_i;
					assign req_d = (lock_q ? req_q : req_i);
					always @(posedge clk_i or negedge rst_ni) begin : p_lock_reg
						if (!rst_ni)
							lock_q <= 1'sb0;
						else if (flush_i)
							lock_q <= 1'sb0;
						else
							lock_q <= lock_d;
					end
					always @(posedge clk_i or negedge rst_ni) begin : p_req_regs
						if (!rst_ni)
							req_q <= 1'sb0;
						else if (flush_i)
							req_q <= 1'sb0;
						else
							req_q <= req_d;
					end
				end
				else begin : gen_no_lock
					assign req_d = req_i;
				end
				function automatic [NumLevels - 1:0] sv2v_cast_5699A;
					input reg [NumLevels - 1:0] inp;
					sv2v_cast_5699A = inp;
				endfunction
				assign rr_d = (gnt_i && req_o ? (rr_q == sv2v_cast_5699A(NumIn - 1) ? {NumLevels {1'sb0}} : rr_q + 1'b1) : rr_q);
				always @(posedge clk_i or negedge rst_ni) begin : p_rr_regs
					if (!rst_ni)
						rr_q <= 1'sb0;
					else if (flush_i)
						rr_q <= 1'sb0;
					else
						rr_q <= rr_d;
				end
			end
			assign gnt_nodes[0] = gnt_i;
			genvar level;
			for (level = 0; $unsigned(level) < NumLevels; level = level + 1) begin : gen_levels
				genvar l;
				for (l = 0; l < (2 ** level); l = l + 1) begin : gen_level
					wire sel;
					localparam [31:0] idx0 = ((2 ** level) - 1) + l;
					localparam [31:0] idx1 = ((2 ** (level + 1)) - 1) + (l * 2);
					if ($unsigned(level) == (NumLevels - 1)) begin : gen_first_level
						if (($unsigned(l) * 2) < (NumIn - 1)) begin : genblk1
							assign req_nodes[idx0] = req_d[l * 2] | req_d[(l * 2) + 1];
							assign sel = ~req_d[l * 2] | (req_d[(l * 2) + 1] & rr_q[(NumLevels - 1) - level]);
							function automatic [NumLevels - 1:0] sv2v_cast_5699A;
								input reg [NumLevels - 1:0] inp;
								sv2v_cast_5699A = inp;
							endfunction
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_5699A(sel);
							assign data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] = (sel ? data_i[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + (((l * 2) + 1) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] : data_i[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((l * 2) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))]);
							assign gnt_o[l * 2] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2])) & ~sel;
							assign gnt_o[(l * 2) + 1] = (gnt_nodes[idx0] & (AxiVldRdy | req_d[(l * 2) + 1])) & sel;
						end
						if (($unsigned(l) * 2) == (NumIn - 1)) begin : genblk2
							assign req_nodes[idx0] = req_d[l * 2];
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = 1'sb0;
							assign data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] = data_i[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((l * 2) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))];
							assign gnt_o[l * 2] = gnt_nodes[idx0] & (AxiVldRdy | req_d[l * 2]);
						end
						if (($unsigned(l) * 2) > (NumIn - 1)) begin : genblk3
							assign req_nodes[idx0] = 1'b0;
							assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = sv2v_cast_BB0BC(1'sb0);
							assign data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] = sv2v_cast_BB0BC(1'sb0);
						end
					end
					else begin : gen_other_levels
						assign req_nodes[idx0] = req_nodes[idx1] | req_nodes[idx1 + 1];
						assign sel = ~req_nodes[idx1] | (req_nodes[idx1 + 1] & rr_q[(NumLevels - 1) - level]);
						function automatic [NumLevels - 1:0] sv2v_cast_5699A;
							input reg [NumLevels - 1:0] inp;
							sv2v_cast_5699A = inp;
						endfunction
						assign index_nodes[(((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * NumLevels+:NumLevels] = (sel ? sv2v_cast_5699A({1'b1, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}) : sv2v_cast_5699A({1'b0, index_nodes[((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * NumLevels) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 2 : (((NumLevels - $unsigned(level)) - 2) + (((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))) - 1)-:(((NumLevels - $unsigned(level)) - 2) >= 0 ? (NumLevels - $unsigned(level)) - 1 : 3 - (NumLevels - $unsigned(level)))]}));
						assign data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx0 : ((2 ** NumLevels) - 2) - idx0) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] = (sel ? data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx1 + 1 : ((2 ** NumLevels) - 2) - (idx1 + 1)) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))] : data_nodes[((DataType_WIDTH + 7) >= 0 ? 0 : DataType_WIDTH + 7) + ((((2 ** NumLevels) - 2) >= 0 ? idx1 : ((2 ** NumLevels) - 2) - idx1) * ((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7)))+:((DataType_WIDTH + 7) >= 0 ? DataType_WIDTH + 8 : 1 - (DataType_WIDTH + 7))]);
						assign gnt_nodes[idx1] = gnt_nodes[idx0] & ~sel;
						assign gnt_nodes[idx1 + 1] = gnt_nodes[idx0] & sel;
					end
				end
			end
		end
	endgenerate
endmodule
module lfsr_8bit (
	clk_i,
	rst_ni,
	en_i,
	refill_way_oh,
	refill_way_bin
);
	parameter [7:0] SEED = 8'b00000000;
	parameter [31:0] WIDTH = 8;
	input wire clk_i;
	input wire rst_ni;
	input wire en_i;
	output reg [WIDTH - 1:0] refill_way_oh;
	output reg [$clog2(WIDTH) - 1:0] refill_way_bin;
	localparam [31:0] LOG_WIDTH = $clog2(WIDTH);
	reg [7:0] shift_d;
	reg [7:0] shift_q;
	always @(*) begin : sv2v_autoblock_1
		reg shift_in;
		shift_in = !(((shift_q[7] ^ shift_q[3]) ^ shift_q[2]) ^ shift_q[1]);
		shift_d = shift_q;
		if (en_i)
			shift_d = {shift_q[6:0], shift_in};
		refill_way_oh = 'b0;
		refill_way_oh[shift_q[LOG_WIDTH - 1:0]] = 1'b1;
		refill_way_bin = shift_q;
	end
	always @(posedge clk_i or negedge rst_ni) begin : proc_
		if (~rst_ni)
			shift_q <= SEED;
		else
			shift_q <= shift_d;
	end
endmodule
module shift_reg_1F3E0_50B1B (
	clk_i,
	rst_ni,
	d_i,
	d_o
);
	parameter signed [31:0] dtype_riscv_XLEN = 0;
	parameter [31:0] Depth = 1;
	input wire clk_i;
	input wire rst_ni;
	input wire [((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0))) - 1:0] d_i;
	output reg [((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0))) - 1:0] d_o;
	generate
		if (Depth == 0) begin : genblk1
			wire [(4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0)):1] sv2v_tmp_021F4;
			assign sv2v_tmp_021F4 = d_i;
			always @(*) d_o = sv2v_tmp_021F4;
		end
		else if (Depth == 1) begin : genblk1
			always @(posedge clk_i or negedge rst_ni)
				if (~rst_ni)
					d_o <= 1'sb0;
				else
					d_o <= d_i;
		end
		else if (Depth > 1) begin : genblk1
			wire [(Depth * ((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0)))) - 1:0] reg_d;
			reg [(Depth * ((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0)))) - 1:0] reg_q;
			wire [(4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0)):1] sv2v_tmp_6C962;
			assign sv2v_tmp_6C962 = reg_q[(Depth - 1) * ((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0)))+:(4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0))];
			always @(*) d_o = sv2v_tmp_6C962;
			assign reg_d = {reg_q[((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0))) * (((Depth - 2) >= 0 ? Depth - 2 : ((Depth - 2) + ((Depth - 2) >= 0 ? Depth - 1 : 3 - Depth)) - 1) - (((Depth - 2) >= 0 ? Depth - 1 : 3 - Depth) - 1))+:((4 + dtype_riscv_XLEN) + (((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0) >= 0 ? (dtype_riscv_XLEN + dtype_riscv_XLEN) + 1 : 1 - ((dtype_riscv_XLEN + dtype_riscv_XLEN) + 0))) * ((Depth - 2) >= 0 ? Depth - 1 : 3 - Depth)], d_i};
			always @(posedge clk_i or negedge rst_ni)
				if (~rst_ni)
					reg_q <= 1'sb0;
				else
					reg_q <= reg_d;
		end
	endgenerate
endmodule
module pmp (
	addr_i,
	access_type_i,
	priv_lvl_i,
	conf_addr_i,
	conf_i,
	allow_o
);
	parameter [31:0] PLEN = 34;
	parameter [31:0] PMP_LEN = 32;
	parameter [31:0] NR_ENTRIES = 4;
	input wire [PLEN - 1:0] addr_i;
	input wire [2:0] access_type_i;
	input wire [1:0] priv_lvl_i;
	input wire [(16 * PMP_LEN) - 1:0] conf_addr_i;
	input wire [127:0] conf_i;
	output reg allow_o;
	generate
		if (NR_ENTRIES > 0) begin : gen_pmp
			wire [NR_ENTRIES - 1:0] match;
			genvar i;
			for (i = 0; i < NR_ENTRIES; i = i + 1) begin : genblk1
				wire [PMP_LEN - 1:0] conf_addr_prev;
				assign conf_addr_prev = (i == 0 ? {PMP_LEN {1'sb0}} : conf_addr_i[(i - 1) * PMP_LEN+:PMP_LEN]);
				pmp_entry #(
					.PLEN(PLEN),
					.PMP_LEN(PMP_LEN)
				) i_pmp_entry(
					.addr_i(addr_i),
					.conf_addr_i(conf_addr_i[i * PMP_LEN+:PMP_LEN]),
					.conf_addr_prev_i(conf_addr_prev),
					.conf_addr_mode_i(conf_i[(i * 8) + 4-:2]),
					.match_o(match[i])
				);
			end
			always @(*) begin : sv2v_autoblock_1
				reg [0:1] _sv2v_jump;
				_sv2v_jump = 2'b00;
				begin : sv2v_autoblock_2
					reg signed [31:0] i;
					allow_o = 1'b0;
					begin : sv2v_autoblock_3
						reg signed [31:0] _sv2v_value_on_break;
						for (i = 0; i < NR_ENTRIES; i = i + 1)
							if (_sv2v_jump < 2'b10) begin
								_sv2v_jump = 2'b00;
								if ((priv_lvl_i != 2'b11) || conf_i[(i * 8) + 7]) begin
									if (match[i]) begin
										if ((access_type_i & conf_i[(i * 8) + 2-:3]) != access_type_i)
											allow_o = 1'b0;
										else
											allow_o = 1'b1;
										_sv2v_jump = 2'b10;
									end
								end
								_sv2v_value_on_break = i;
							end
						if (!(_sv2v_jump < 2'b10))
							i = _sv2v_value_on_break;
						if (_sv2v_jump != 2'b11)
							_sv2v_jump = 2'b00;
					end
					if (_sv2v_jump == 2'b00) begin
						if (i == NR_ENTRIES) begin
							if (priv_lvl_i == 2'b11)
								allow_o = 1'b1;
							else
								allow_o = 1'b0;
						end
					end
				end
			end
		end
		else begin : genblk1
			wire [1:1] sv2v_tmp_6821D;
			assign sv2v_tmp_6821D = 1'b1;
			always @(*) allow_o = sv2v_tmp_6821D;
		end
	endgenerate
endmodule
module pmp_entry (
	addr_i,
	conf_addr_i,
	conf_addr_prev_i,
	conf_addr_mode_i,
	match_o
);
	parameter [31:0] PLEN = 56;
	parameter [31:0] PMP_LEN = 54;
	input wire [PLEN - 1:0] addr_i;
	input wire [PMP_LEN - 1:0] conf_addr_i;
	input wire [PMP_LEN - 1:0] conf_addr_prev_i;
	input wire [1:0] conf_addr_mode_i;
	output reg match_o;
	wire [PLEN - 1:0] conf_addr_n;
	wire [$clog2(PLEN) - 1:0] trail_ones;
	assign conf_addr_n = ~conf_addr_i;
	lzc #(
		.WIDTH(PLEN),
		.MODE(1'b0)
	) i_lzc(
		.in_i(conf_addr_n),
		.cnt_o(trail_ones),
		.empty_o()
	);
	always @(*)
		case (conf_addr_mode_i)
			2'b01:
				if ((addr_i >= (conf_addr_prev_i << 2)) && (addr_i < (conf_addr_i << 2)))
					match_o = 1'b1;
				else
					match_o = 1'b0;
			2'b10, 2'b11: begin : sv2v_autoblock_1
				reg [PLEN - 1:0] base;
				reg [PLEN - 1:0] mask;
				reg [31:0] size;
				if (conf_addr_mode_i == 2'b10)
					size = 2;
				else
					size = trail_ones + 3;
				mask = 1'sb1 << size;
				base = (conf_addr_i << 2) & mask;
				match_o = ((addr_i & mask) == base ? 1'b1 : 1'b0);
			end
			2'b00: match_o = 1'b0;
			default: match_o = 0;
		endcase
endmodule
module CVA6CoreBlackbox (
	clk_i,
	rst_ni,
	boot_addr_i,
	hart_id_i,
	irq_i,
	ipi_i,
	time_irq_i,
	debug_req_i,
	trace_o,
	axi_resp_i_aw_ready,
	axi_req_o_aw_valid,
	axi_req_o_aw_bits_id,
	axi_req_o_aw_bits_addr,
	axi_req_o_aw_bits_len,
	axi_req_o_aw_bits_size,
	axi_req_o_aw_bits_burst,
	axi_req_o_aw_bits_lock,
	axi_req_o_aw_bits_cache,
	axi_req_o_aw_bits_prot,
	axi_req_o_aw_bits_qos,
	axi_req_o_aw_bits_region,
	axi_req_o_aw_bits_atop,
	axi_req_o_aw_bits_user,
	axi_resp_i_w_ready,
	axi_req_o_w_valid,
	axi_req_o_w_bits_data,
	axi_req_o_w_bits_strb,
	axi_req_o_w_bits_last,
	axi_req_o_w_bits_user,
	axi_resp_i_ar_ready,
	axi_req_o_ar_valid,
	axi_req_o_ar_bits_id,
	axi_req_o_ar_bits_addr,
	axi_req_o_ar_bits_len,
	axi_req_o_ar_bits_size,
	axi_req_o_ar_bits_burst,
	axi_req_o_ar_bits_lock,
	axi_req_o_ar_bits_cache,
	axi_req_o_ar_bits_prot,
	axi_req_o_ar_bits_qos,
	axi_req_o_ar_bits_region,
	axi_req_o_ar_bits_user,
	axi_req_o_b_ready,
	axi_resp_i_b_valid,
	axi_resp_i_b_bits_id,
	axi_resp_i_b_bits_resp,
	axi_resp_i_b_bits_user,
	axi_req_o_r_ready,
	axi_resp_i_r_valid,
	axi_resp_i_r_bits_id,
	axi_resp_i_r_bits_data,
	axi_resp_i_r_bits_resp,
	axi_resp_i_r_bits_last,
	axi_resp_i_r_bits_user
);
	parameter TRACEPORT_SZ = 0;
	parameter XLEN = 0;
	parameter RAS_ENTRIES = 0;
	parameter BTB_ENTRIES = 0;
	parameter BHT_ENTRIES = 0;
	parameter [63:0] EXEC_REG_CNT = 0;
	parameter [63:0] EXEC_REG_BASE_0 = 0;
	parameter [63:0] EXEC_REG_SZ_0 = 0;
	parameter [63:0] EXEC_REG_BASE_1 = 0;
	parameter [63:0] EXEC_REG_SZ_1 = 0;
	parameter [63:0] EXEC_REG_BASE_2 = 0;
	parameter [63:0] EXEC_REG_SZ_2 = 0;
	parameter [63:0] EXEC_REG_BASE_3 = 0;
	parameter [63:0] EXEC_REG_SZ_3 = 0;
	parameter [63:0] EXEC_REG_BASE_4 = 0;
	parameter [63:0] EXEC_REG_SZ_4 = 0;
	parameter [63:0] CACHE_REG_CNT = 0;
	parameter [63:0] CACHE_REG_BASE_0 = 0;
	parameter [63:0] CACHE_REG_SZ_0 = 0;
	parameter [63:0] CACHE_REG_BASE_1 = 0;
	parameter [63:0] CACHE_REG_SZ_1 = 0;
	parameter [63:0] CACHE_REG_BASE_2 = 0;
	parameter [63:0] CACHE_REG_SZ_2 = 0;
	parameter [63:0] CACHE_REG_BASE_3 = 0;
	parameter [63:0] CACHE_REG_SZ_3 = 0;
	parameter [63:0] CACHE_REG_BASE_4 = 0;
	parameter [63:0] CACHE_REG_SZ_4 = 0;
	parameter [63:0] DEBUG_BASE = 0;
	parameter AXI_ADDRESS_WIDTH = 0;
	parameter AXI_DATA_WIDTH = 0;
	parameter AXI_USER_WIDTH = 0;
	parameter AXI_ID_WIDTH = 0;
	parameter PMP_ENTRIES = 0;
	input clk_i;
	input rst_ni;
	input [XLEN - 1:0] boot_addr_i;
	input [63:0] hart_id_i;
	input [1:0] irq_i;
	input ipi_i;
	input time_irq_i;
	input debug_req_i;
	output wire [TRACEPORT_SZ - 1:0] trace_o;
	input axi_resp_i_aw_ready;
	output wire axi_req_o_aw_valid;
	output wire [AXI_ID_WIDTH - 1:0] axi_req_o_aw_bits_id;
	output wire [AXI_ADDRESS_WIDTH - 1:0] axi_req_o_aw_bits_addr;
	output wire [7:0] axi_req_o_aw_bits_len;
	output wire [2:0] axi_req_o_aw_bits_size;
	output wire [1:0] axi_req_o_aw_bits_burst;
	output wire axi_req_o_aw_bits_lock;
	output wire [3:0] axi_req_o_aw_bits_cache;
	output wire [2:0] axi_req_o_aw_bits_prot;
	output wire [3:0] axi_req_o_aw_bits_qos;
	output wire [3:0] axi_req_o_aw_bits_region;
	output wire [5:0] axi_req_o_aw_bits_atop;
	output wire [AXI_USER_WIDTH - 1:0] axi_req_o_aw_bits_user;
	input axi_resp_i_w_ready;
	output wire axi_req_o_w_valid;
	output wire [AXI_DATA_WIDTH - 1:0] axi_req_o_w_bits_data;
	output wire [(AXI_DATA_WIDTH / 8) - 1:0] axi_req_o_w_bits_strb;
	output wire axi_req_o_w_bits_last;
	output wire [AXI_USER_WIDTH - 1:0] axi_req_o_w_bits_user;
	input axi_resp_i_ar_ready;
	output wire axi_req_o_ar_valid;
	output wire [AXI_ID_WIDTH - 1:0] axi_req_o_ar_bits_id;
	output wire [AXI_ADDRESS_WIDTH - 1:0] axi_req_o_ar_bits_addr;
	output wire [7:0] axi_req_o_ar_bits_len;
	output wire [2:0] axi_req_o_ar_bits_size;
	output wire [1:0] axi_req_o_ar_bits_burst;
	output wire axi_req_o_ar_bits_lock;
	output wire [3:0] axi_req_o_ar_bits_cache;
	output wire [2:0] axi_req_o_ar_bits_prot;
	output wire [3:0] axi_req_o_ar_bits_qos;
	output wire [3:0] axi_req_o_ar_bits_region;
	output wire [AXI_USER_WIDTH - 1:0] axi_req_o_ar_bits_user;
	output wire axi_req_o_b_ready;
	input axi_resp_i_b_valid;
	input [AXI_ID_WIDTH - 1:0] axi_resp_i_b_bits_id;
	input [1:0] axi_resp_i_b_bits_resp;
	input [AXI_USER_WIDTH - 1:0] axi_resp_i_b_bits_user;
	output wire axi_req_o_r_ready;
	input axi_resp_i_r_valid;
	input [AXI_ID_WIDTH - 1:0] axi_resp_i_r_bits_id;
	input [AXI_DATA_WIDTH - 1:0] axi_resp_i_r_bits_data;
	input [1:0] axi_resp_i_r_bits_resp;
	input axi_resp_i_r_bits_last;
	input [AXI_USER_WIDTH - 1:0] axi_resp_i_r_bits_user;
	localparam ariane_pkg_NrMaxRules = 16;
	function automatic [31:0] sv2v_cast_32;
		input reg [31:0] inp;
		sv2v_cast_32 = inp;
	endfunction
	function automatic [1023:0] sv2v_cast_1024;
		input reg [1023:0] inp;
		sv2v_cast_1024 = inp;
	endfunction
	localparam [6433:0] CVA6SocCfg = {RAS_ENTRIES, BTB_ENTRIES, BHT_ENTRIES, 2080'h0, sv2v_cast_32(EXEC_REG_CNT), sv2v_cast_1024({EXEC_REG_BASE_4, EXEC_REG_BASE_3, EXEC_REG_BASE_2, EXEC_REG_BASE_1, EXEC_REG_BASE_0}), sv2v_cast_1024({EXEC_REG_SZ_4, EXEC_REG_SZ_3, EXEC_REG_SZ_2, EXEC_REG_SZ_1, EXEC_REG_SZ_0}), sv2v_cast_32(CACHE_REG_CNT), sv2v_cast_1024({CACHE_REG_BASE_4, CACHE_REG_BASE_3, CACHE_REG_BASE_2, CACHE_REG_BASE_1, CACHE_REG_BASE_0}), sv2v_cast_1024({CACHE_REG_SZ_4, CACHE_REG_SZ_3, CACHE_REG_SZ_2, CACHE_REG_SZ_1, CACHE_REG_SZ_0}), 2'b10, DEBUG_BASE, sv2v_cast_32(PMP_ENTRIES)};
	localparam ariane_axi_AddrWidth = 64;
	localparam ariane_axi_IdWidth = 4;
	localparam ariane_axi_UserWidth = 1;
	localparam ariane_axi_DataWidth = 64;
	localparam ariane_axi_StrbWidth = 8;
	wire [280:0] ariane_axi_req;
	wire [83:0] ariane_axi_resp;
	ariane #(.ArianeCfg(CVA6SocCfg)) i_ariane(
		.clk_i(clk_i),
		.rst_ni(rst_ni),
		.boot_addr_i(boot_addr_i),
		.hart_id_i(hart_id_i),
		.irq_i(irq_i),
		.ipi_i(ipi_i),
		.time_irq_i(time_irq_i),
		.debug_req_i(debug_req_i),
		.axi_req_o(ariane_axi_req),
		.axi_resp_i(ariane_axi_resp)
	);
	assign trace_o = 1'sb0;
	localparam _param_F9970_AXI_ADDR_WIDTH = AXI_ADDRESS_WIDTH;
	localparam _param_F9970_AXI_DATA_WIDTH = AXI_DATA_WIDTH;
	localparam _param_F9970_AXI_ID_WIDTH = AXI_ID_WIDTH;
	localparam _param_F9970_AXI_USER_WIDTH = AXI_USER_WIDTH;
	generate
		if (1) begin : axi_slave_bus
			localparam AXI_ADDR_WIDTH = _param_F9970_AXI_ADDR_WIDTH;
			localparam AXI_DATA_WIDTH = _param_F9970_AXI_DATA_WIDTH;
			localparam AXI_ID_WIDTH = _param_F9970_AXI_ID_WIDTH;
			localparam AXI_USER_WIDTH = _param_F9970_AXI_USER_WIDTH;
			localparam AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
			wire [AXI_ID_WIDTH - 1:0] aw_id;
			wire [AXI_ADDR_WIDTH - 1:0] aw_addr;
			wire [7:0] aw_len;
			wire [2:0] aw_size;
			wire [1:0] aw_burst;
			wire aw_lock;
			wire [3:0] aw_cache;
			wire [2:0] aw_prot;
			wire [3:0] aw_qos;
			wire [5:0] aw_atop;
			wire [3:0] aw_region;
			wire [AXI_USER_WIDTH - 1:0] aw_user;
			wire aw_valid;
			wire aw_ready;
			wire [AXI_DATA_WIDTH - 1:0] w_data;
			wire [AXI_STRB_WIDTH - 1:0] w_strb;
			wire w_last;
			wire [AXI_USER_WIDTH - 1:0] w_user;
			wire w_valid;
			wire w_ready;
			wire [AXI_ID_WIDTH - 1:0] b_id;
			wire [1:0] b_resp;
			wire [AXI_USER_WIDTH - 1:0] b_user;
			wire b_valid;
			wire b_ready;
			wire [AXI_ID_WIDTH - 1:0] ar_id;
			wire [AXI_ADDR_WIDTH - 1:0] ar_addr;
			wire [7:0] ar_len;
			wire [2:0] ar_size;
			wire [1:0] ar_burst;
			wire ar_lock;
			wire [3:0] ar_cache;
			wire [2:0] ar_prot;
			wire [3:0] ar_qos;
			wire [3:0] ar_region;
			wire [AXI_USER_WIDTH - 1:0] ar_user;
			wire ar_valid;
			wire ar_ready;
			wire [AXI_ID_WIDTH - 1:0] r_id;
			wire [AXI_DATA_WIDTH - 1:0] r_data;
			wire [1:0] r_resp;
			wire r_last;
			wire [AXI_USER_WIDTH - 1:0] r_user;
			wire r_valid;
			wire r_ready;
		end
		if (1) begin : i_axi_master_connect_ariane
			localparam ariane_axi_AddrWidth = 64;
			localparam ariane_axi_IdWidth = 4;
			localparam ariane_axi_UserWidth = 1;
			localparam ariane_axi_DataWidth = 64;
			localparam ariane_axi_StrbWidth = 8;
			wire [280:0] axi_req_i;
			wire [83:0] axi_resp_o;
			assign CVA6CoreBlackbox.axi_slave_bus.aw_id = axi_req_i[280-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_addr = axi_req_i[276-:64];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_len = axi_req_i[212-:8];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_size = axi_req_i[204-:3];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_burst = axi_req_i[201-:2];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_lock = axi_req_i[199];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_cache = axi_req_i[198-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_prot = axi_req_i[194-:3];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_qos = axi_req_i[191-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_atop = axi_req_i[183-:6];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_region = axi_req_i[187-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.aw_user = 1'sb0;
			assign CVA6CoreBlackbox.axi_slave_bus.aw_valid = axi_req_i[176];
			assign axi_resp_o[83] = CVA6CoreBlackbox.axi_slave_bus.aw_ready;
			assign CVA6CoreBlackbox.axi_slave_bus.w_data = axi_req_i[175-:64];
			assign CVA6CoreBlackbox.axi_slave_bus.w_strb = axi_req_i[111-:8];
			assign CVA6CoreBlackbox.axi_slave_bus.w_last = axi_req_i[103];
			assign CVA6CoreBlackbox.axi_slave_bus.w_user = 1'sb0;
			assign CVA6CoreBlackbox.axi_slave_bus.w_valid = axi_req_i[101];
			assign axi_resp_o[81] = CVA6CoreBlackbox.axi_slave_bus.w_ready;
			assign axi_resp_o[79-:4] = CVA6CoreBlackbox.axi_slave_bus.b_id;
			assign axi_resp_o[75-:2] = CVA6CoreBlackbox.axi_slave_bus.b_resp;
			assign axi_resp_o[80] = CVA6CoreBlackbox.axi_slave_bus.b_valid;
			assign CVA6CoreBlackbox.axi_slave_bus.b_ready = axi_req_i[100];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_id = axi_req_i[99-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_addr = axi_req_i[95-:64];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_len = axi_req_i[31-:8];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_size = axi_req_i[23-:3];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_burst = axi_req_i[20-:2];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_lock = axi_req_i[18];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_cache = axi_req_i[17-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_prot = axi_req_i[13-:3];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_qos = axi_req_i[10-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_region = axi_req_i[6-:4];
			assign CVA6CoreBlackbox.axi_slave_bus.ar_user = 1'sb0;
			assign CVA6CoreBlackbox.axi_slave_bus.ar_valid = axi_req_i[1];
			assign axi_resp_o[82] = CVA6CoreBlackbox.axi_slave_bus.ar_ready;
			assign axi_resp_o[71-:4] = CVA6CoreBlackbox.axi_slave_bus.r_id;
			assign axi_resp_o[67-:64] = CVA6CoreBlackbox.axi_slave_bus.r_data;
			assign axi_resp_o[3-:2] = CVA6CoreBlackbox.axi_slave_bus.r_resp;
			assign axi_resp_o[1] = CVA6CoreBlackbox.axi_slave_bus.r_last;
			assign axi_resp_o[72] = CVA6CoreBlackbox.axi_slave_bus.r_valid;
			assign CVA6CoreBlackbox.axi_slave_bus.r_ready = axi_req_i[0];
		end
	endgenerate
	assign i_axi_master_connect_ariane.axi_req_i = ariane_axi_req;
	assign ariane_axi_resp = i_axi_master_connect_ariane.axi_resp_o;
	localparam _param_71D8A_AXI_ADDR_WIDTH = AXI_ADDRESS_WIDTH;
	localparam _param_71D8A_AXI_DATA_WIDTH = AXI_DATA_WIDTH;
	localparam _param_71D8A_AXI_ID_WIDTH = AXI_ID_WIDTH;
	localparam _param_71D8A_AXI_USER_WIDTH = AXI_USER_WIDTH;
	generate
		if (1) begin : axi_master_bus
			localparam AXI_ADDR_WIDTH = _param_71D8A_AXI_ADDR_WIDTH;
			localparam AXI_DATA_WIDTH = _param_71D8A_AXI_DATA_WIDTH;
			localparam AXI_ID_WIDTH = _param_71D8A_AXI_ID_WIDTH;
			localparam AXI_USER_WIDTH = _param_71D8A_AXI_USER_WIDTH;
			localparam AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
			wire [AXI_ID_WIDTH - 1:0] aw_id;
			wire [AXI_ADDR_WIDTH - 1:0] aw_addr;
			wire [7:0] aw_len;
			wire [2:0] aw_size;
			wire [1:0] aw_burst;
			wire aw_lock;
			wire [3:0] aw_cache;
			wire [2:0] aw_prot;
			wire [3:0] aw_qos;
			wire [5:0] aw_atop;
			wire [3:0] aw_region;
			wire [AXI_USER_WIDTH - 1:0] aw_user;
			wire aw_valid;
			wire aw_ready;
			wire [AXI_DATA_WIDTH - 1:0] w_data;
			wire [AXI_STRB_WIDTH - 1:0] w_strb;
			wire w_last;
			wire [AXI_USER_WIDTH - 1:0] w_user;
			wire w_valid;
			wire w_ready;
			wire [AXI_ID_WIDTH - 1:0] b_id;
			wire [1:0] b_resp;
			wire [AXI_USER_WIDTH - 1:0] b_user;
			wire b_valid;
			wire b_ready;
			wire [AXI_ID_WIDTH - 1:0] ar_id;
			wire [AXI_ADDR_WIDTH - 1:0] ar_addr;
			wire [7:0] ar_len;
			wire [2:0] ar_size;
			wire [1:0] ar_burst;
			wire ar_lock;
			wire [3:0] ar_cache;
			wire [2:0] ar_prot;
			wire [3:0] ar_qos;
			wire [3:0] ar_region;
			wire [AXI_USER_WIDTH - 1:0] ar_user;
			wire ar_valid;
			wire ar_ready;
			wire [AXI_ID_WIDTH - 1:0] r_id;
			wire [AXI_DATA_WIDTH - 1:0] r_data;
			wire [1:0] r_resp;
			wire r_last;
			wire [AXI_USER_WIDTH - 1:0] r_user;
			wire r_valid;
			wire r_ready;
		end
	endgenerate
	localparam _param_F7A30_AXI_ADDR_WIDTH = AXI_ADDRESS_WIDTH;
	localparam _param_F7A30_AXI_DATA_WIDTH = AXI_DATA_WIDTH;
	localparam _param_F7A30_AXI_ID_WIDTH = AXI_ID_WIDTH;
	localparam _param_F7A30_AXI_USER_WIDTH = AXI_USER_WIDTH;
	localparam _param_F7A30_AXI_MAX_WRITE_TXNS = 1;
	localparam _param_F7A30_RISCV_WORD_WIDTH = XLEN;
	generate
		if (1) begin : i_axi_riscv_atomics
			localparam [31:0] AXI_ADDR_WIDTH = _param_F7A30_AXI_ADDR_WIDTH;
			localparam [31:0] AXI_DATA_WIDTH = _param_F7A30_AXI_DATA_WIDTH;
			localparam [31:0] AXI_ID_WIDTH = _param_F7A30_AXI_ID_WIDTH;
			localparam [31:0] AXI_USER_WIDTH = _param_F7A30_AXI_USER_WIDTH;
			localparam [31:0] AXI_MAX_WRITE_TXNS = _param_F7A30_AXI_MAX_WRITE_TXNS;
			localparam [31:0] RISCV_WORD_WIDTH = _param_F7A30_RISCV_WORD_WIDTH;
			localparam [31:0] AXI_STRB_WIDTH = AXI_DATA_WIDTH / 8;
			wire clk_i;
			wire rst_ni;
			axi_riscv_atomics #(
				.AXI_ADDR_WIDTH(AXI_ADDR_WIDTH),
				.AXI_DATA_WIDTH(AXI_DATA_WIDTH),
				.AXI_ID_WIDTH(AXI_ID_WIDTH),
				.AXI_USER_WIDTH(AXI_USER_WIDTH),
				.AXI_MAX_WRITE_TXNS(AXI_MAX_WRITE_TXNS),
				.RISCV_WORD_WIDTH(RISCV_WORD_WIDTH)
			) i_atomics(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.slv_aw_addr_i(CVA6CoreBlackbox.axi_slave_bus.aw_addr),
				.slv_aw_prot_i(CVA6CoreBlackbox.axi_slave_bus.aw_prot),
				.slv_aw_region_i(CVA6CoreBlackbox.axi_slave_bus.aw_region),
				.slv_aw_atop_i(CVA6CoreBlackbox.axi_slave_bus.aw_atop),
				.slv_aw_len_i(CVA6CoreBlackbox.axi_slave_bus.aw_len),
				.slv_aw_size_i(CVA6CoreBlackbox.axi_slave_bus.aw_size),
				.slv_aw_burst_i(CVA6CoreBlackbox.axi_slave_bus.aw_burst),
				.slv_aw_lock_i(CVA6CoreBlackbox.axi_slave_bus.aw_lock),
				.slv_aw_cache_i(CVA6CoreBlackbox.axi_slave_bus.aw_cache),
				.slv_aw_qos_i(CVA6CoreBlackbox.axi_slave_bus.aw_qos),
				.slv_aw_id_i(CVA6CoreBlackbox.axi_slave_bus.aw_id),
				.slv_aw_user_i(CVA6CoreBlackbox.axi_slave_bus.aw_user),
				.slv_aw_ready_o(CVA6CoreBlackbox.axi_slave_bus.aw_ready),
				.slv_aw_valid_i(CVA6CoreBlackbox.axi_slave_bus.aw_valid),
				.slv_ar_addr_i(CVA6CoreBlackbox.axi_slave_bus.ar_addr),
				.slv_ar_prot_i(CVA6CoreBlackbox.axi_slave_bus.ar_prot),
				.slv_ar_region_i(CVA6CoreBlackbox.axi_slave_bus.ar_region),
				.slv_ar_len_i(CVA6CoreBlackbox.axi_slave_bus.ar_len),
				.slv_ar_size_i(CVA6CoreBlackbox.axi_slave_bus.ar_size),
				.slv_ar_burst_i(CVA6CoreBlackbox.axi_slave_bus.ar_burst),
				.slv_ar_lock_i(CVA6CoreBlackbox.axi_slave_bus.ar_lock),
				.slv_ar_cache_i(CVA6CoreBlackbox.axi_slave_bus.ar_cache),
				.slv_ar_qos_i(CVA6CoreBlackbox.axi_slave_bus.ar_qos),
				.slv_ar_id_i(CVA6CoreBlackbox.axi_slave_bus.ar_id),
				.slv_ar_user_i(CVA6CoreBlackbox.axi_slave_bus.ar_user),
				.slv_ar_ready_o(CVA6CoreBlackbox.axi_slave_bus.ar_ready),
				.slv_ar_valid_i(CVA6CoreBlackbox.axi_slave_bus.ar_valid),
				.slv_w_data_i(CVA6CoreBlackbox.axi_slave_bus.w_data),
				.slv_w_strb_i(CVA6CoreBlackbox.axi_slave_bus.w_strb),
				.slv_w_user_i(CVA6CoreBlackbox.axi_slave_bus.w_user),
				.slv_w_last_i(CVA6CoreBlackbox.axi_slave_bus.w_last),
				.slv_w_ready_o(CVA6CoreBlackbox.axi_slave_bus.w_ready),
				.slv_w_valid_i(CVA6CoreBlackbox.axi_slave_bus.w_valid),
				.slv_r_data_o(CVA6CoreBlackbox.axi_slave_bus.r_data),
				.slv_r_resp_o(CVA6CoreBlackbox.axi_slave_bus.r_resp),
				.slv_r_last_o(CVA6CoreBlackbox.axi_slave_bus.r_last),
				.slv_r_id_o(CVA6CoreBlackbox.axi_slave_bus.r_id),
				.slv_r_user_o(CVA6CoreBlackbox.axi_slave_bus.r_user),
				.slv_r_ready_i(CVA6CoreBlackbox.axi_slave_bus.r_ready),
				.slv_r_valid_o(CVA6CoreBlackbox.axi_slave_bus.r_valid),
				.slv_b_resp_o(CVA6CoreBlackbox.axi_slave_bus.b_resp),
				.slv_b_id_o(CVA6CoreBlackbox.axi_slave_bus.b_id),
				.slv_b_user_o(CVA6CoreBlackbox.axi_slave_bus.b_user),
				.slv_b_ready_i(CVA6CoreBlackbox.axi_slave_bus.b_ready),
				.slv_b_valid_o(CVA6CoreBlackbox.axi_slave_bus.b_valid),
				.mst_aw_addr_o(CVA6CoreBlackbox.axi_master_bus.aw_addr),
				.mst_aw_prot_o(CVA6CoreBlackbox.axi_master_bus.aw_prot),
				.mst_aw_region_o(CVA6CoreBlackbox.axi_master_bus.aw_region),
				.mst_aw_atop_o(CVA6CoreBlackbox.axi_master_bus.aw_atop),
				.mst_aw_len_o(CVA6CoreBlackbox.axi_master_bus.aw_len),
				.mst_aw_size_o(CVA6CoreBlackbox.axi_master_bus.aw_size),
				.mst_aw_burst_o(CVA6CoreBlackbox.axi_master_bus.aw_burst),
				.mst_aw_lock_o(CVA6CoreBlackbox.axi_master_bus.aw_lock),
				.mst_aw_cache_o(CVA6CoreBlackbox.axi_master_bus.aw_cache),
				.mst_aw_qos_o(CVA6CoreBlackbox.axi_master_bus.aw_qos),
				.mst_aw_id_o(CVA6CoreBlackbox.axi_master_bus.aw_id),
				.mst_aw_user_o(CVA6CoreBlackbox.axi_master_bus.aw_user),
				.mst_aw_ready_i(CVA6CoreBlackbox.axi_master_bus.aw_ready),
				.mst_aw_valid_o(CVA6CoreBlackbox.axi_master_bus.aw_valid),
				.mst_ar_addr_o(CVA6CoreBlackbox.axi_master_bus.ar_addr),
				.mst_ar_prot_o(CVA6CoreBlackbox.axi_master_bus.ar_prot),
				.mst_ar_region_o(CVA6CoreBlackbox.axi_master_bus.ar_region),
				.mst_ar_len_o(CVA6CoreBlackbox.axi_master_bus.ar_len),
				.mst_ar_size_o(CVA6CoreBlackbox.axi_master_bus.ar_size),
				.mst_ar_burst_o(CVA6CoreBlackbox.axi_master_bus.ar_burst),
				.mst_ar_lock_o(CVA6CoreBlackbox.axi_master_bus.ar_lock),
				.mst_ar_cache_o(CVA6CoreBlackbox.axi_master_bus.ar_cache),
				.mst_ar_qos_o(CVA6CoreBlackbox.axi_master_bus.ar_qos),
				.mst_ar_id_o(CVA6CoreBlackbox.axi_master_bus.ar_id),
				.mst_ar_user_o(CVA6CoreBlackbox.axi_master_bus.ar_user),
				.mst_ar_ready_i(CVA6CoreBlackbox.axi_master_bus.ar_ready),
				.mst_ar_valid_o(CVA6CoreBlackbox.axi_master_bus.ar_valid),
				.mst_w_data_o(CVA6CoreBlackbox.axi_master_bus.w_data),
				.mst_w_strb_o(CVA6CoreBlackbox.axi_master_bus.w_strb),
				.mst_w_user_o(CVA6CoreBlackbox.axi_master_bus.w_user),
				.mst_w_last_o(CVA6CoreBlackbox.axi_master_bus.w_last),
				.mst_w_ready_i(CVA6CoreBlackbox.axi_master_bus.w_ready),
				.mst_w_valid_o(CVA6CoreBlackbox.axi_master_bus.w_valid),
				.mst_r_data_i(CVA6CoreBlackbox.axi_master_bus.r_data),
				.mst_r_resp_i(CVA6CoreBlackbox.axi_master_bus.r_resp),
				.mst_r_last_i(CVA6CoreBlackbox.axi_master_bus.r_last),
				.mst_r_id_i(CVA6CoreBlackbox.axi_master_bus.r_id),
				.mst_r_user_i(CVA6CoreBlackbox.axi_master_bus.r_user),
				.mst_r_ready_o(CVA6CoreBlackbox.axi_master_bus.r_ready),
				.mst_r_valid_i(CVA6CoreBlackbox.axi_master_bus.r_valid),
				.mst_b_resp_i(CVA6CoreBlackbox.axi_master_bus.b_resp),
				.mst_b_id_i(CVA6CoreBlackbox.axi_master_bus.b_id),
				.mst_b_user_i(CVA6CoreBlackbox.axi_master_bus.b_user),
				.mst_b_ready_o(CVA6CoreBlackbox.axi_master_bus.b_ready),
				.mst_b_valid_i(CVA6CoreBlackbox.axi_master_bus.b_valid)
			);
		end
	endgenerate
	assign i_axi_riscv_atomics.clk_i = clk_i;
	assign i_axi_riscv_atomics.rst_ni = rst_ni;
	assign axi_master_bus.aw_ready = axi_resp_i_aw_ready;
	assign axi_req_o_aw_valid = axi_master_bus.aw_valid;
	assign axi_req_o_aw_bits_id = axi_master_bus.aw_id;
	assign axi_req_o_aw_bits_addr = axi_master_bus.aw_addr;
	assign axi_req_o_aw_bits_len = axi_master_bus.aw_len;
	assign axi_req_o_aw_bits_size = axi_master_bus.aw_size;
	assign axi_req_o_aw_bits_burst = axi_master_bus.aw_burst;
	assign axi_req_o_aw_bits_lock = axi_master_bus.aw_lock;
	assign axi_req_o_aw_bits_cache = axi_master_bus.aw_cache;
	assign axi_req_o_aw_bits_prot = axi_master_bus.aw_prot;
	assign axi_req_o_aw_bits_qos = axi_master_bus.aw_qos;
	assign axi_req_o_aw_bits_region = axi_master_bus.aw_region;
	assign axi_req_o_aw_bits_atop = axi_master_bus.aw_atop;
	assign axi_req_o_aw_bits_user = axi_master_bus.aw_user;
	assign axi_master_bus.w_ready = axi_resp_i_w_ready;
	assign axi_req_o_w_valid = axi_master_bus.w_valid;
	assign axi_req_o_w_bits_data = axi_master_bus.w_data;
	assign axi_req_o_w_bits_strb = axi_master_bus.w_strb;
	assign axi_req_o_w_bits_last = axi_master_bus.w_last;
	assign axi_req_o_w_bits_user = axi_master_bus.w_user;
	assign axi_master_bus.ar_ready = axi_resp_i_ar_ready;
	assign axi_req_o_ar_valid = axi_master_bus.ar_valid;
	assign axi_req_o_ar_bits_id = axi_master_bus.ar_id;
	assign axi_req_o_ar_bits_addr = axi_master_bus.ar_addr;
	assign axi_req_o_ar_bits_len = axi_master_bus.ar_len;
	assign axi_req_o_ar_bits_size = axi_master_bus.ar_size;
	assign axi_req_o_ar_bits_burst = axi_master_bus.ar_burst;
	assign axi_req_o_ar_bits_lock = axi_master_bus.ar_lock;
	assign axi_req_o_ar_bits_cache = axi_master_bus.ar_cache;
	assign axi_req_o_ar_bits_prot = axi_master_bus.ar_prot;
	assign axi_req_o_ar_bits_qos = axi_master_bus.ar_qos;
	assign axi_req_o_ar_bits_region = axi_master_bus.ar_region;
	assign axi_req_o_ar_bits_user = axi_master_bus.ar_user;
	assign axi_req_o_b_ready = axi_master_bus.b_ready;
	assign axi_master_bus.b_valid = axi_resp_i_b_valid;
	assign axi_master_bus.b_id = axi_resp_i_b_bits_id;
	assign axi_master_bus.b_resp = axi_resp_i_b_bits_resp;
	assign axi_master_bus.b_user = axi_resp_i_b_bits_user;
	assign axi_req_o_r_ready = axi_master_bus.r_ready;
	assign axi_master_bus.r_valid = axi_resp_i_r_valid;
	assign axi_master_bus.r_id = axi_resp_i_r_bits_id;
	assign axi_master_bus.r_data = axi_resp_i_r_bits_data;
	assign axi_master_bus.r_resp = axi_resp_i_r_bits_resp;
	assign axi_master_bus.r_last = axi_resp_i_r_bits_last;
	assign axi_master_bus.r_user = axi_resp_i_r_bits_user;
endmodule