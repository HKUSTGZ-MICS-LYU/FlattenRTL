module wrapper #(
    parameter RTL___csr_regfile___f_reset_rsps___guarded=32'd1,
    parameter RTL___stage1_f_reset_reqs___guarded=32'd1,
    parameter RTL___stage1_f_reset_rsps___guarded=32'd1,
    parameter RTL___stage2_f_reset_reqs___guarded=32'd1,
    parameter RTL___stage2_f_reset_rsps___guarded=32'd1,
    parameter RTL___stage3_f_reset_reqs___guarded=32'd1,
    parameter RTL___stage3_f_reset_rsps___guarded=32'd1,
parameter RTL___f_reset_reqs___width=32'd1,
parameter RTL___f_reset_reqs___guarded=32'd1,
parameter RTL___f_reset_rsps___width=32'd1,
parameter RTL___f_reset_rsps___guarded=32'd1,
parameter RTL___gpr_regfile___f_reset_rsps___guarded=32'd1,
parameter RTL___gpr_regfile___regfile___addr_width=32'd5,
parameter RTL___gpr_regfile___regfile___data_width=32'd32,
parameter RTL___gpr_regfile___regfile___lo=5'h0,
parameter RTL___gpr_regfile___regfile___hi=5'd31,
parameter RTL___near_mem___dcache___dmem_not_imem=1'd1,
parameter RTL___near_mem___icache___dmem_not_imem=1'd0,
parameter RTL___near_mem___dcache___f_fabric_write_reqs___width=32'd99,
parameter RTL___near_mem___dcache___f_fabric_write_reqs___guarded=32'd1,
parameter RTL___near_mem___dcache___f_reset_reqs___width=32'd1,
parameter RTL___near_mem___dcache___f_reset_reqs___guarded=32'd1,
parameter RTL___near_mem___dcache___f_reset_rsps___width=32'd1,
parameter RTL___near_mem___dcache___f_reset_rsps___guarded=32'd1,
parameter RTL___near_mem___dcache___master_xactor_f_rd_addr___width=32'd97,
parameter RTL___near_mem___dcache___master_xactor_f_rd_addr___guarded=32'd1,
parameter RTL___near_mem___dcache___master_xactor_f_rd_data___width=32'd71,
parameter RTL___near_mem___dcache___master_xactor_f_rd_data___guarded=32'd1,
parameter RTL___near_mem___dcache___master_xactor_f_wr_addr___width=32'd97,
parameter RTL___near_mem___dcache___master_xactor_f_wr_addr___guarded=32'd1,
parameter RTL___near_mem___dcache___master_xactor_f_wr_data___width=32'd73,
parameter RTL___near_mem___dcache___master_xactor_f_wr_data___guarded=32'd1,
parameter RTL___near_mem___dcache___master_xactor_f_wr_resp___width=32'd6,
parameter RTL___near_mem___dcache___master_xactor_f_wr_resp___guarded=32'd1,
parameter RTL___near_mem___icache___f_fabric_write_reqs___width=32'd99,
parameter RTL___near_mem___icache___f_fabric_write_reqs___guarded=32'd1,
parameter RTL___near_mem___icache___f_reset_reqs___width=32'd1,
parameter RTL___near_mem___icache___f_reset_reqs___guarded=32'd1,
parameter RTL___near_mem___icache___f_reset_rsps___width=32'd1,
parameter RTL___near_mem___icache___f_reset_rsps___guarded=32'd1,
parameter RTL___near_mem___icache___master_xactor_f_rd_addr___width=32'd97,
parameter RTL___near_mem___icache___master_xactor_f_rd_addr___guarded=32'd1,
parameter RTL___near_mem___icache___master_xactor_f_rd_data___width=32'd71,
parameter RTL___near_mem___icache___master_xactor_f_rd_data___guarded=32'd1,
parameter RTL___near_mem___icache___master_xactor_f_wr_addr___width=32'd97,
parameter RTL___near_mem___icache___master_xactor_f_wr_addr___guarded=32'd1,
parameter RTL___near_mem___icache___master_xactor_f_wr_data___width=32'd73,
parameter RTL___near_mem___icache___master_xactor_f_wr_data___guarded=32'd1,
parameter RTL___near_mem___icache___master_xactor_f_wr_resp___width=32'd6,
parameter RTL___near_mem___icache___master_xactor_f_wr_resp___guarded=32'd1,
parameter RTL___near_mem___dcache___ram_state_and_ctag_cset___PIPELINED=1'd0,
parameter RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDR_WIDTH=32'd7,
parameter RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH=32'd23,
parameter RTL___near_mem___dcache___ram_state_and_ctag_cset___MEMSIZE=8'd128,
parameter RTL___near_mem___dcache___ram_word64_set___PIPELINED=1'd0,
parameter RTL___near_mem___dcache___ram_word64_set___ADDR_WIDTH=32'd9,
parameter RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH=32'd64,
parameter RTL___near_mem___dcache___ram_word64_set___MEMSIZE=10'd512,
parameter RTL___near_mem___icache___ram_state_and_ctag_cset___PIPELINED=1'd0,
parameter RTL___near_mem___icache___ram_state_and_ctag_cset___ADDR_WIDTH=32'd7,
parameter RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH=32'd23,
parameter RTL___near_mem___icache___ram_state_and_ctag_cset___MEMSIZE=8'd128,
parameter RTL___near_mem___icache___ram_word64_set___PIPELINED=1'd0,
parameter RTL___near_mem___icache___ram_word64_set___ADDR_WIDTH=32'd9,
parameter RTL___near_mem___icache___ram_word64_set___DATA_WIDTH=32'd64,
parameter RTL___near_mem___icache___ram_word64_set___MEMSIZE=10'd512,
parameter RTL___near_mem___f_reset_rsps___guarded=32'd1)(
__ILA_I_inst,
__ISSUE__,
__VLG_I_EN_hart0_server_reset_request_put,
__VLG_I_EN_hart0_server_reset_response_get,
__VLG_I_EN_set_verbosity,
__VLG_I_dmem_master_arready,
__VLG_I_dmem_master_awready,
__VLG_I_dmem_master_bid,
__VLG_I_dmem_master_bresp,
__VLG_I_dmem_master_bvalid,
__VLG_I_dmem_master_rdata,
__VLG_I_dmem_master_rid,
__VLG_I_dmem_master_rlast,
__VLG_I_dmem_master_rresp,
__VLG_I_dmem_master_rvalid,
__VLG_I_dmem_master_wready,
__VLG_I_hart0_server_reset_request_put,
__VLG_I_imem_master_arready,
__VLG_I_imem_master_awready,
__VLG_I_imem_master_bid,
__VLG_I_imem_master_bresp,
__VLG_I_imem_master_bvalid,
__VLG_I_imem_master_rdata,
__VLG_I_imem_master_rid,
__VLG_I_imem_master_rlast,
__VLG_I_imem_master_rresp,
__VLG_I_imem_master_rvalid,
__VLG_I_imem_master_wready,
__VLG_I_set_verbosity_logdelay,
__VLG_I_set_verbosity_verbosity,
____auxvar10__recorder_init__,
____auxvar11__recorder_init__,
____auxvar12__recorder_init__,
____auxvar13__recorder_init__,
____auxvar14__recorder_init__,
____auxvar15__recorder_init__,
____auxvar16__recorder_init__,
____auxvar17__recorder_init__,
____auxvar18__recorder_init__,
____auxvar19__recorder_init__,
____auxvar1__recorder_init__,
____auxvar20__recorder_init__,
____auxvar21__recorder_init__,
____auxvar22__recorder_init__,
____auxvar23__recorder_init__,
____auxvar24__recorder_init__,
____auxvar25__recorder_init__,
____auxvar26__recorder_init__,
____auxvar27__recorder_init__,
____auxvar28__recorder_init__,
____auxvar29__recorder_init__,
____auxvar2__recorder_init__,
____auxvar30__recorder_init__,
____auxvar31__recorder_init__,
____auxvar32__recorder_init__,
____auxvar33__recorder_init__,
____auxvar34__recorder_init__,
____auxvar35__recorder_init__,
____auxvar36__recorder_init__,
____auxvar37__recorder_init__,
____auxvar38__recorder_init__,
____auxvar3__recorder_init__,
____auxvar4__recorder_init__,
____auxvar5__recorder_init__,
____auxvar6__recorder_init__,
____auxvar7__recorder_init__,
____auxvar8__recorder_init__,
____auxvar9__recorder_init__,
clk,
dummy_reset,
rst,
RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__csr_regfile__DOT__rg_nmi,
RTL__DOT__csr_regfile__DOT__rg_state,
RTL__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_,
RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_,
RTL__DOT__near_mem$EN_dmem_req,
RTL__DOT__near_mem$dmem_exc,
RTL__DOT__near_mem$dmem_req_addr,
RTL__DOT__near_mem$dmem_req_f3,
RTL__DOT__near_mem$dmem_req_op,
RTL__DOT__near_mem$dmem_req_store_value,
RTL__DOT__near_mem$dmem_word64,
RTL__DOT__near_mem$imem_instr,
RTL__DOT__near_mem$imem_pc,
RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg,
RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr,
RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa,
RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg,
RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg,
RTL__DOT__rg_cur_priv,
RTL__DOT__rg_retiring$EN,
RTL__DOT__rg_run_on_reset,
RTL__DOT__rg_state,
RTL__DOT__rg_trap_instr,
RTL__DOT__s1_to_s2$D_IN,
RTL__DOT__s1_to_s2$EN,
RTL__DOT__s2_to_s3$D_IN,
RTL__DOT__s2_to_s3$EN,
RTL__DOT__s3_deq$D_IN,
RTL__DOT__s3_deq$EN,
RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage1_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage1_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage1_rg_full,
RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage2_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage2_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage2_rg_full,
RTL__DOT__stage2_rg_stage2,
RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg,
RTL__DOT__stage3_f_reset_reqs__DOT__full_reg,
RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg,
RTL__DOT__stage3_f_reset_rsps__DOT__full_reg,
RTL__DOT__stage3_rg_full,
__EDCOND__,
__IEND__,
__ILA_SO_load_addr,
__ILA_SO_load_data,
__ILA_SO_load_en,
__ILA_SO_load_size,
__ILA_SO_pc,
__ILA_SO_store_addr,
__ILA_SO_store_data,
__ILA_SO_store_en,
__ILA_SO_store_size,
__ILA_SO_x0,
__ILA_SO_x1,
__ILA_SO_x10,
__ILA_SO_x11,
__ILA_SO_x12,
__ILA_SO_x13,
__ILA_SO_x14,
__ILA_SO_x15,
__ILA_SO_x16,
__ILA_SO_x17,
__ILA_SO_x18,
__ILA_SO_x19,
__ILA_SO_x2,
__ILA_SO_x20,
__ILA_SO_x21,
__ILA_SO_x22,
__ILA_SO_x23,
__ILA_SO_x24,
__ILA_SO_x25,
__ILA_SO_x26,
__ILA_SO_x27,
__ILA_SO_x28,
__ILA_SO_x29,
__ILA_SO_x3,
__ILA_SO_x30,
__ILA_SO_x31,
__ILA_SO_x4,
__ILA_SO_x5,
__ILA_SO_x6,
__ILA_SO_x7,
__ILA_SO_x8,
__ILA_SO_x9,
__VLG_II_m_external_interrupt_req_set_not_clear,
__VLG_II_nmi_req_set_not_clear,
__VLG_II_s_external_interrupt_req_set_not_clear,
__VLG_II_software_interrupt_req_set_not_clear,
__VLG_II_timer_interrupt_req_set_not_clear,
__VLG_O_RDY_hart0_server_reset_request_put,
__VLG_O_RDY_hart0_server_reset_response_get,
__VLG_O_RDY_set_verbosity,
__VLG_O_dmem_master_araddr,
__VLG_O_dmem_master_arburst,
__VLG_O_dmem_master_arcache,
__VLG_O_dmem_master_arid,
__VLG_O_dmem_master_arlen,
__VLG_O_dmem_master_arlock,
__VLG_O_dmem_master_arprot,
__VLG_O_dmem_master_arqos,
__VLG_O_dmem_master_arregion,
__VLG_O_dmem_master_arsize,
__VLG_O_dmem_master_arvalid,
__VLG_O_dmem_master_awaddr,
__VLG_O_dmem_master_awburst,
__VLG_O_dmem_master_awcache,
__VLG_O_dmem_master_awid,
__VLG_O_dmem_master_awlen,
__VLG_O_dmem_master_awlock,
__VLG_O_dmem_master_awprot,
__VLG_O_dmem_master_awqos,
__VLG_O_dmem_master_awregion,
__VLG_O_dmem_master_awsize,
__VLG_O_dmem_master_awvalid,
__VLG_O_dmem_master_bready,
__VLG_O_dmem_master_rready,
__VLG_O_dmem_master_wdata,
__VLG_O_dmem_master_wlast,
__VLG_O_dmem_master_wstrb,
__VLG_O_dmem_master_wvalid,
__VLG_O_hart0_server_reset_response_get,
__VLG_O_imem_master_araddr,
__VLG_O_imem_master_arburst,
__VLG_O_imem_master_arcache,
__VLG_O_imem_master_arid,
__VLG_O_imem_master_arlen,
__VLG_O_imem_master_arlock,
__VLG_O_imem_master_arprot,
__VLG_O_imem_master_arqos,
__VLG_O_imem_master_arregion,
__VLG_O_imem_master_arsize,
__VLG_O_imem_master_arvalid,
__VLG_O_imem_master_awaddr,
__VLG_O_imem_master_awburst,
__VLG_O_imem_master_awcache,
__VLG_O_imem_master_awid,
__VLG_O_imem_master_awlen,
__VLG_O_imem_master_awlock,
__VLG_O_imem_master_awprot,
__VLG_O_imem_master_awqos,
__VLG_O_imem_master_awregion,
__VLG_O_imem_master_awsize,
__VLG_O_imem_master_awvalid,
__VLG_O_imem_master_bready,
__VLG_O_imem_master_rready,
__VLG_O_imem_master_wdata,
__VLG_O_imem_master_wlast,
__VLG_O_imem_master_wstrb,
__VLG_O_imem_master_wvalid,
__all_assert_wire__,
__all_assume_wire__,
__auxvar0__delay_d_0,
__sanitycheck_wire__,
end_of_pipeline,
input_map_assume___p0__,
invariant_assume__p10__,
invariant_assume__p11__,
invariant_assume__p12__,
invariant_assume__p13__,
invariant_assume__p14__,
invariant_assume__p15__,
invariant_assume__p16__,
invariant_assume__p17__,
invariant_assume__p18__,
invariant_assume__p19__,
invariant_assume__p1__,
invariant_assume__p20__,
invariant_assume__p21__,
invariant_assume__p22__,
invariant_assume__p23__,
invariant_assume__p24__,
invariant_assume__p25__,
invariant_assume__p26__,
invariant_assume__p27__,
invariant_assume__p28__,
invariant_assume__p29__,
invariant_assume__p2__,
invariant_assume__p30__,
invariant_assume__p31__,
invariant_assume__p32__,
invariant_assume__p3__,
invariant_assume__p4__,
invariant_assume__p5__,
invariant_assume__p6__,
invariant_assume__p7__,
invariant_assume__p8__,
invariant_assume__p9__,
issue_decode__p33__,
issue_valid__p34__,
mem_req_addr,
mem_req_en,
mem_req_funct3,
mem_req_op,
mem_req_rd_data,
mem_req_wd_data,
monitor_s1,
monitor_s1_already_enter_cond,
monitor_s1_already_exit_cond,
monitor_s2_enter_cond,
monitor_s2_exit_cond,
monitor_s3_enter_cond,
monitor_s3_exit_cond,
monitor_s4_enter_cond,
monitor_s4_exit_cond,
noreset__p35__,
post_value_holder__p36__,
post_value_holder__p37__,
post_value_holder__p38__,
post_value_holder__p39__,
post_value_holder__p40__,
post_value_holder__p41__,
post_value_holder__p42__,
post_value_holder__p43__,
post_value_holder__p44__,
post_value_holder__p45__,
post_value_holder__p46__,
post_value_holder__p47__,
post_value_holder__p48__,
post_value_holder__p49__,
post_value_holder__p50__,
post_value_holder__p51__,
post_value_holder__p52__,
post_value_holder__p53__,
post_value_holder__p54__,
post_value_holder__p55__,
post_value_holder__p56__,
post_value_holder__p57__,
post_value_holder__p58__,
post_value_holder__p59__,
post_value_holder__p60__,
post_value_holder__p61__,
post_value_holder__p62__,
post_value_holder__p63__,
post_value_holder__p64__,
post_value_holder__p65__,
post_value_holder__p66__,
post_value_holder__p67__,
post_value_holder__p68__,
post_value_holder__p69__,
post_value_holder__p70__,
post_value_holder__p71__,
post_value_holder__p72__,
post_value_holder__p73__,
post_value_holder_overly_constrained__p153__,
post_value_holder_overly_constrained__p154__,
post_value_holder_overly_constrained__p155__,
post_value_holder_overly_constrained__p156__,
post_value_holder_overly_constrained__p157__,
post_value_holder_overly_constrained__p158__,
post_value_holder_overly_constrained__p159__,
post_value_holder_overly_constrained__p160__,
post_value_holder_overly_constrained__p161__,
post_value_holder_overly_constrained__p162__,
post_value_holder_overly_constrained__p163__,
post_value_holder_overly_constrained__p164__,
post_value_holder_overly_constrained__p165__,
post_value_holder_overly_constrained__p166__,
post_value_holder_overly_constrained__p167__,
post_value_holder_overly_constrained__p168__,
post_value_holder_overly_constrained__p169__,
post_value_holder_overly_constrained__p170__,
post_value_holder_overly_constrained__p171__,
post_value_holder_overly_constrained__p172__,
post_value_holder_overly_constrained__p173__,
post_value_holder_overly_constrained__p174__,
post_value_holder_overly_constrained__p175__,
post_value_holder_overly_constrained__p176__,
post_value_holder_overly_constrained__p177__,
post_value_holder_overly_constrained__p178__,
post_value_holder_overly_constrained__p179__,
post_value_holder_overly_constrained__p180__,
post_value_holder_overly_constrained__p181__,
post_value_holder_overly_constrained__p182__,
post_value_holder_overly_constrained__p183__,
post_value_holder_overly_constrained__p184__,
post_value_holder_overly_constrained__p185__,
post_value_holder_overly_constrained__p186__,
post_value_holder_overly_constrained__p187__,
post_value_holder_overly_constrained__p188__,
post_value_holder_overly_constrained__p189__,
post_value_holder_overly_constrained__p190__,
post_value_holder_triggered__p191__,
post_value_holder_triggered__p192__,
post_value_holder_triggered__p193__,
post_value_holder_triggered__p194__,
post_value_holder_triggered__p195__,
post_value_holder_triggered__p196__,
post_value_holder_triggered__p197__,
post_value_holder_triggered__p198__,
post_value_holder_triggered__p199__,
post_value_holder_triggered__p200__,
post_value_holder_triggered__p201__,
post_value_holder_triggered__p202__,
post_value_holder_triggered__p203__,
post_value_holder_triggered__p204__,
post_value_holder_triggered__p205__,
post_value_holder_triggered__p206__,
post_value_holder_triggered__p207__,
post_value_holder_triggered__p208__,
post_value_holder_triggered__p209__,
post_value_holder_triggered__p210__,
post_value_holder_triggered__p211__,
post_value_holder_triggered__p212__,
post_value_holder_triggered__p213__,
post_value_holder_triggered__p214__,
post_value_holder_triggered__p215__,
post_value_holder_triggered__p216__,
post_value_holder_triggered__p217__,
post_value_holder_triggered__p218__,
post_value_holder_triggered__p219__,
post_value_holder_triggered__p220__,
post_value_holder_triggered__p221__,
post_value_holder_triggered__p222__,
post_value_holder_triggered__p223__,
post_value_holder_triggered__p224__,
post_value_holder_triggered__p225__,
post_value_holder_triggered__p226__,
post_value_holder_triggered__p227__,
post_value_holder_triggered__p228__,
rfassumptions__p74__,
rfassumptions__p75__,
rfassumptions__p76__,
s2_enter,
s2_exit,
s3_enter,
s3_exit,
s4_enter,
variable_map_assert__p118__,
variable_map_assert__p119__,
variable_map_assert__p120__,
variable_map_assert__p121__,
variable_map_assert__p122__,
variable_map_assert__p123__,
variable_map_assert__p124__,
variable_map_assert__p125__,
variable_map_assert__p126__,
variable_map_assert__p127__,
variable_map_assert__p128__,
variable_map_assert__p129__,
variable_map_assert__p130__,
variable_map_assert__p131__,
variable_map_assert__p132__,
variable_map_assert__p133__,
variable_map_assert__p134__,
variable_map_assert__p135__,
variable_map_assert__p136__,
variable_map_assert__p137__,
variable_map_assert__p138__,
variable_map_assert__p139__,
variable_map_assert__p140__,
variable_map_assert__p141__,
variable_map_assert__p142__,
variable_map_assert__p143__,
variable_map_assert__p144__,
variable_map_assert__p145__,
variable_map_assert__p146__,
variable_map_assert__p147__,
variable_map_assert__p148__,
variable_map_assert__p149__,
variable_map_assert__p150__,
variable_map_assert__p151__,
variable_map_assert__p152__,
variable_map_assume___p100__,
variable_map_assume___p101__,
variable_map_assume___p102__,
variable_map_assume___p103__,
variable_map_assume___p104__,
variable_map_assume___p105__,
variable_map_assume___p106__,
variable_map_assume___p107__,
variable_map_assume___p108__,
variable_map_assume___p109__,
variable_map_assume___p110__,
variable_map_assume___p111__,
variable_map_assume___p112__,
variable_map_assume___p113__,
variable_map_assume___p114__,
variable_map_assume___p115__,
variable_map_assume___p116__,
variable_map_assume___p117__,
variable_map_assume___p77__,
variable_map_assume___p78__,
variable_map_assume___p79__,
variable_map_assume___p80__,
variable_map_assume___p81__,
variable_map_assume___p82__,
variable_map_assume___p83__,
variable_map_assume___p84__,
variable_map_assume___p85__,
variable_map_assume___p86__,
variable_map_assume___p87__,
variable_map_assume___p88__,
variable_map_assume___p89__,
variable_map_assume___p90__,
variable_map_assume___p91__,
variable_map_assume___p92__,
variable_map_assume___p93__,
variable_map_assume___p94__,
variable_map_assume___p95__,
variable_map_assume___p96__,
variable_map_assume___p97__,
variable_map_assume___p98__,
variable_map_assume___p99__,
__CYCLE_CNT__,
__START__,
__STARTED__,
__ENDED__,
__2ndENDED__,
__RESETED__,
__auxvar10__recorder,
__auxvar10__recorder_sn_vhold,
__auxvar10__recorder_sn_condmet,
__auxvar11__recorder,
__auxvar11__recorder_sn_vhold,
__auxvar11__recorder_sn_condmet,
__auxvar12__recorder,
__auxvar12__recorder_sn_vhold,
__auxvar12__recorder_sn_condmet,
__auxvar13__recorder,
__auxvar13__recorder_sn_vhold,
__auxvar13__recorder_sn_condmet,
__auxvar14__recorder,
__auxvar14__recorder_sn_vhold,
__auxvar14__recorder_sn_condmet,
__auxvar15__recorder,
__auxvar15__recorder_sn_vhold,
__auxvar15__recorder_sn_condmet,
__auxvar16__recorder,
__auxvar16__recorder_sn_vhold,
__auxvar16__recorder_sn_condmet,
__auxvar17__recorder,
__auxvar17__recorder_sn_vhold,
__auxvar17__recorder_sn_condmet,
__auxvar18__recorder,
__auxvar18__recorder_sn_vhold,
__auxvar18__recorder_sn_condmet,
__auxvar19__recorder,
__auxvar19__recorder_sn_vhold,
__auxvar19__recorder_sn_condmet,
__auxvar1__recorder,
__auxvar1__recorder_sn_vhold,
__auxvar1__recorder_sn_condmet,
__auxvar20__recorder,
__auxvar20__recorder_sn_vhold,
__auxvar20__recorder_sn_condmet,
__auxvar21__recorder,
__auxvar21__recorder_sn_vhold,
__auxvar21__recorder_sn_condmet,
__auxvar22__recorder,
__auxvar22__recorder_sn_vhold,
__auxvar22__recorder_sn_condmet,
__auxvar23__recorder,
__auxvar23__recorder_sn_vhold,
__auxvar23__recorder_sn_condmet,
__auxvar24__recorder,
__auxvar24__recorder_sn_vhold,
__auxvar24__recorder_sn_condmet,
__auxvar25__recorder,
__auxvar25__recorder_sn_vhold,
__auxvar25__recorder_sn_condmet,
__auxvar26__recorder,
__auxvar26__recorder_sn_vhold,
__auxvar26__recorder_sn_condmet,
__auxvar27__recorder,
__auxvar27__recorder_sn_vhold,
__auxvar27__recorder_sn_condmet,
__auxvar28__recorder,
__auxvar28__recorder_sn_vhold,
__auxvar28__recorder_sn_condmet,
__auxvar29__recorder,
__auxvar29__recorder_sn_vhold,
__auxvar29__recorder_sn_condmet,
__auxvar2__recorder,
__auxvar2__recorder_sn_vhold,
__auxvar2__recorder_sn_condmet,
__auxvar30__recorder,
__auxvar30__recorder_sn_vhold,
__auxvar30__recorder_sn_condmet,
__auxvar31__recorder,
__auxvar31__recorder_sn_vhold,
__auxvar31__recorder_sn_condmet,
__auxvar32__recorder,
__auxvar32__recorder_sn_vhold,
__auxvar32__recorder_sn_condmet,
__auxvar33__recorder,
__auxvar33__recorder_sn_vhold,
__auxvar33__recorder_sn_condmet,
__auxvar34__recorder,
__auxvar34__recorder_sn_vhold,
__auxvar34__recorder_sn_condmet,
__auxvar35__recorder,
__auxvar35__recorder_sn_vhold,
__auxvar35__recorder_sn_condmet,
__auxvar36__recorder,
__auxvar36__recorder_sn_vhold,
__auxvar36__recorder_sn_condmet,
__auxvar37__recorder,
__auxvar37__recorder_sn_vhold,
__auxvar37__recorder_sn_condmet,
__auxvar38__recorder,
__auxvar38__recorder_sn_vhold,
__auxvar38__recorder_sn_condmet,
__auxvar3__recorder,
__auxvar3__recorder_sn_vhold,
__auxvar3__recorder_sn_condmet,
__auxvar4__recorder,
__auxvar4__recorder_sn_vhold,
__auxvar4__recorder_sn_condmet,
__auxvar5__recorder,
__auxvar5__recorder_sn_vhold,
__auxvar5__recorder_sn_condmet,
__auxvar6__recorder,
__auxvar6__recorder_sn_vhold,
__auxvar6__recorder_sn_condmet,
__auxvar7__recorder,
__auxvar7__recorder_sn_vhold,
__auxvar7__recorder_sn_condmet,
__auxvar8__recorder,
__auxvar8__recorder_sn_vhold,
__auxvar8__recorder_sn_condmet,
__auxvar9__recorder,
__auxvar9__recorder_sn_vhold,
__auxvar9__recorder_sn_condmet,
__auxvar0__delay_d_1,
monitor_s1_already,
monitor_s2,
monitor_s3,
monitor_s4
);
input     [31:0] __ILA_I_inst;
input            __ISSUE__;
input            __VLG_I_EN_hart0_server_reset_request_put;
input            __VLG_I_EN_hart0_server_reset_response_get;
input            __VLG_I_EN_set_verbosity;
input            __VLG_I_dmem_master_arready;
input            __VLG_I_dmem_master_awready;
input      [3:0] __VLG_I_dmem_master_bid;
input      [1:0] __VLG_I_dmem_master_bresp;
input            __VLG_I_dmem_master_bvalid;
input     [63:0] __VLG_I_dmem_master_rdata;
input      [3:0] __VLG_I_dmem_master_rid;
input            __VLG_I_dmem_master_rlast;
input      [1:0] __VLG_I_dmem_master_rresp;
input            __VLG_I_dmem_master_rvalid;
input            __VLG_I_dmem_master_wready;
input            __VLG_I_hart0_server_reset_request_put;
input            __VLG_I_imem_master_arready;
input            __VLG_I_imem_master_awready;
input      [3:0] __VLG_I_imem_master_bid;
input      [1:0] __VLG_I_imem_master_bresp;
input            __VLG_I_imem_master_bvalid;
input     [63:0] __VLG_I_imem_master_rdata;
input      [3:0] __VLG_I_imem_master_rid;
input            __VLG_I_imem_master_rlast;
input      [1:0] __VLG_I_imem_master_rresp;
input            __VLG_I_imem_master_rvalid;
input            __VLG_I_imem_master_wready;
input     [63:0] __VLG_I_set_verbosity_logdelay;
input      [3:0] __VLG_I_set_verbosity_verbosity;
input     [31:0] ____auxvar10__recorder_init__;
input     [31:0] ____auxvar11__recorder_init__;
input     [31:0] ____auxvar12__recorder_init__;
input     [31:0] ____auxvar13__recorder_init__;
input     [31:0] ____auxvar14__recorder_init__;
input     [31:0] ____auxvar15__recorder_init__;
input     [31:0] ____auxvar16__recorder_init__;
input     [31:0] ____auxvar17__recorder_init__;
input     [31:0] ____auxvar18__recorder_init__;
input     [31:0] ____auxvar19__recorder_init__;
input     [31:0] ____auxvar1__recorder_init__;
input     [31:0] ____auxvar20__recorder_init__;
input     [31:0] ____auxvar21__recorder_init__;
input     [31:0] ____auxvar22__recorder_init__;
input     [31:0] ____auxvar23__recorder_init__;
input     [31:0] ____auxvar24__recorder_init__;
input     [31:0] ____auxvar25__recorder_init__;
input     [31:0] ____auxvar26__recorder_init__;
input     [31:0] ____auxvar27__recorder_init__;
input     [31:0] ____auxvar28__recorder_init__;
input     [31:0] ____auxvar29__recorder_init__;
input     [31:0] ____auxvar2__recorder_init__;
input     [31:0] ____auxvar30__recorder_init__;
input     [31:0] ____auxvar31__recorder_init__;
input     [31:0] ____auxvar32__recorder_init__;
input     [31:0] ____auxvar33__recorder_init__;
input            ____auxvar34__recorder_init__;
input      [2:0] ____auxvar35__recorder_init__;
input            ____auxvar36__recorder_init__;
input     [31:0] ____auxvar37__recorder_init__;
input     [31:0] ____auxvar38__recorder_init__;
input     [31:0] ____auxvar3__recorder_init__;
input     [31:0] ____auxvar4__recorder_init__;
input     [31:0] ____auxvar5__recorder_init__;
input     [31:0] ____auxvar6__recorder_init__;
input     [31:0] ____auxvar7__recorder_init__;
input     [31:0] ____auxvar8__recorder_init__;
input     [31:0] ____auxvar9__recorder_init__;
input            clk;
input            dummy_reset;
input            rst;
output            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__csr_regfile__DOT__rg_nmi;
output            RTL__DOT__csr_regfile__DOT__rg_state;
output            RTL__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
output     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
output            RTL__DOT__near_mem$EN_dmem_req;
output            RTL__DOT__near_mem$dmem_exc;
output     [31:0] RTL__DOT__near_mem$dmem_req_addr;
output      [2:0] RTL__DOT__near_mem$dmem_req_f3;
output            RTL__DOT__near_mem$dmem_req_op;
output     [63:0] RTL__DOT__near_mem$dmem_req_store_value;
output     [63:0] RTL__DOT__near_mem$dmem_word64;
output     [31:0] RTL__DOT__near_mem$imem_instr;
output     [31:0] RTL__DOT__near_mem$imem_pc;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
output     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
output     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
output            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
output            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
output      [1:0] RTL__DOT__rg_cur_priv;
output            RTL__DOT__rg_retiring$EN;
output            RTL__DOT__rg_run_on_reset;
output      [3:0] RTL__DOT__rg_state;
output     [31:0] RTL__DOT__rg_trap_instr;
output            RTL__DOT__s1_to_s2$D_IN;
output            RTL__DOT__s1_to_s2$EN;
output            RTL__DOT__s2_to_s3$D_IN;
output            RTL__DOT__s2_to_s3$EN;
output            RTL__DOT__s3_deq$D_IN;
output            RTL__DOT__s3_deq$EN;
output            RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage1_rg_full;
output            RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage2_rg_full;
output    [168:0] RTL__DOT__stage2_rg_stage2;
output            RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
output            RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
output            RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
output            RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
output            RTL__DOT__stage3_rg_full;
output            __EDCOND__;
output            __IEND__;
output     [31:0] __ILA_SO_load_addr;
output     [31:0] __ILA_SO_load_data;
output            __ILA_SO_load_en;
output      [2:0] __ILA_SO_load_size;
output     [31:0] __ILA_SO_pc;
output     [31:0] __ILA_SO_store_addr;
output     [31:0] __ILA_SO_store_data;
output            __ILA_SO_store_en;
output      [2:0] __ILA_SO_store_size;
output     [31:0] __ILA_SO_x0;
output     [31:0] __ILA_SO_x1;
output     [31:0] __ILA_SO_x10;
output     [31:0] __ILA_SO_x11;
output     [31:0] __ILA_SO_x12;
output     [31:0] __ILA_SO_x13;
output     [31:0] __ILA_SO_x14;
output     [31:0] __ILA_SO_x15;
output     [31:0] __ILA_SO_x16;
output     [31:0] __ILA_SO_x17;
output     [31:0] __ILA_SO_x18;
output     [31:0] __ILA_SO_x19;
output     [31:0] __ILA_SO_x2;
output     [31:0] __ILA_SO_x20;
output     [31:0] __ILA_SO_x21;
output     [31:0] __ILA_SO_x22;
output     [31:0] __ILA_SO_x23;
output     [31:0] __ILA_SO_x24;
output     [31:0] __ILA_SO_x25;
output     [31:0] __ILA_SO_x26;
output     [31:0] __ILA_SO_x27;
output     [31:0] __ILA_SO_x28;
output     [31:0] __ILA_SO_x29;
output     [31:0] __ILA_SO_x3;
output     [31:0] __ILA_SO_x30;
output     [31:0] __ILA_SO_x31;
output     [31:0] __ILA_SO_x4;
output     [31:0] __ILA_SO_x5;
output     [31:0] __ILA_SO_x6;
output     [31:0] __ILA_SO_x7;
output     [31:0] __ILA_SO_x8;
output     [31:0] __ILA_SO_x9;
output            __VLG_II_m_external_interrupt_req_set_not_clear;
output            __VLG_II_nmi_req_set_not_clear;
output            __VLG_II_s_external_interrupt_req_set_not_clear;
output            __VLG_II_software_interrupt_req_set_not_clear;
output            __VLG_II_timer_interrupt_req_set_not_clear;
output            __VLG_O_RDY_hart0_server_reset_request_put;
output            __VLG_O_RDY_hart0_server_reset_response_get;
output            __VLG_O_RDY_set_verbosity;
output     [63:0] __VLG_O_dmem_master_araddr;
output      [1:0] __VLG_O_dmem_master_arburst;
output      [3:0] __VLG_O_dmem_master_arcache;
output      [3:0] __VLG_O_dmem_master_arid;
output      [7:0] __VLG_O_dmem_master_arlen;
output            __VLG_O_dmem_master_arlock;
output      [2:0] __VLG_O_dmem_master_arprot;
output      [3:0] __VLG_O_dmem_master_arqos;
output      [3:0] __VLG_O_dmem_master_arregion;
output      [2:0] __VLG_O_dmem_master_arsize;
output            __VLG_O_dmem_master_arvalid;
output     [63:0] __VLG_O_dmem_master_awaddr;
output      [1:0] __VLG_O_dmem_master_awburst;
output      [3:0] __VLG_O_dmem_master_awcache;
output      [3:0] __VLG_O_dmem_master_awid;
output      [7:0] __VLG_O_dmem_master_awlen;
output            __VLG_O_dmem_master_awlock;
output      [2:0] __VLG_O_dmem_master_awprot;
output      [3:0] __VLG_O_dmem_master_awqos;
output      [3:0] __VLG_O_dmem_master_awregion;
output      [2:0] __VLG_O_dmem_master_awsize;
output            __VLG_O_dmem_master_awvalid;
output            __VLG_O_dmem_master_bready;
output            __VLG_O_dmem_master_rready;
output     [63:0] __VLG_O_dmem_master_wdata;
output            __VLG_O_dmem_master_wlast;
output      [7:0] __VLG_O_dmem_master_wstrb;
output            __VLG_O_dmem_master_wvalid;
output            __VLG_O_hart0_server_reset_response_get;
output     [63:0] __VLG_O_imem_master_araddr;
output      [1:0] __VLG_O_imem_master_arburst;
output      [3:0] __VLG_O_imem_master_arcache;
output      [3:0] __VLG_O_imem_master_arid;
output      [7:0] __VLG_O_imem_master_arlen;
output            __VLG_O_imem_master_arlock;
output      [2:0] __VLG_O_imem_master_arprot;
output      [3:0] __VLG_O_imem_master_arqos;
output      [3:0] __VLG_O_imem_master_arregion;
output      [2:0] __VLG_O_imem_master_arsize;
output            __VLG_O_imem_master_arvalid;
output     [63:0] __VLG_O_imem_master_awaddr;
output      [1:0] __VLG_O_imem_master_awburst;
output      [3:0] __VLG_O_imem_master_awcache;
output      [3:0] __VLG_O_imem_master_awid;
output      [7:0] __VLG_O_imem_master_awlen;
output            __VLG_O_imem_master_awlock;
output      [2:0] __VLG_O_imem_master_awprot;
output      [3:0] __VLG_O_imem_master_awqos;
output      [3:0] __VLG_O_imem_master_awregion;
output      [2:0] __VLG_O_imem_master_awsize;
output            __VLG_O_imem_master_awvalid;
output            __VLG_O_imem_master_bready;
output            __VLG_O_imem_master_rready;
output     [63:0] __VLG_O_imem_master_wdata;
output            __VLG_O_imem_master_wlast;
output      [7:0] __VLG_O_imem_master_wstrb;
output            __VLG_O_imem_master_wvalid;
output            __all_assert_wire__;
output            __all_assume_wire__;
output            __auxvar0__delay_d_0;
output            __sanitycheck_wire__;
output            end_of_pipeline;
output            input_map_assume___p0__;
output            invariant_assume__p10__;
output            invariant_assume__p11__;
output            invariant_assume__p12__;
output            invariant_assume__p13__;
output            invariant_assume__p14__;
output            invariant_assume__p15__;
output            invariant_assume__p16__;
output            invariant_assume__p17__;
output            invariant_assume__p18__;
output            invariant_assume__p19__;
output            invariant_assume__p1__;
output            invariant_assume__p20__;
output            invariant_assume__p21__;
output            invariant_assume__p22__;
output            invariant_assume__p23__;
output            invariant_assume__p24__;
output            invariant_assume__p25__;
output            invariant_assume__p26__;
output            invariant_assume__p27__;
output            invariant_assume__p28__;
output            invariant_assume__p29__;
output            invariant_assume__p2__;
output            invariant_assume__p30__;
output            invariant_assume__p31__;
output            invariant_assume__p32__;
output            invariant_assume__p3__;
output            invariant_assume__p4__;
output            invariant_assume__p5__;
output            invariant_assume__p6__;
output            invariant_assume__p7__;
output            invariant_assume__p8__;
output            invariant_assume__p9__;
output            issue_decode__p33__;
output            issue_valid__p34__;
output     [31:0] mem_req_addr;
output            mem_req_en;
output      [2:0] mem_req_funct3;
output            mem_req_op;
output     [31:0] mem_req_rd_data;
output     [31:0] mem_req_wd_data;
output            monitor_s1;
output            monitor_s1_already_enter_cond;
output            monitor_s1_already_exit_cond;
output            monitor_s2_enter_cond;
output            monitor_s2_exit_cond;
output            monitor_s3_enter_cond;
output            monitor_s3_exit_cond;
output            monitor_s4_enter_cond;
output            monitor_s4_exit_cond;
output            noreset__p35__;
output            post_value_holder__p36__;
output            post_value_holder__p37__;
output            post_value_holder__p38__;
output            post_value_holder__p39__;
output            post_value_holder__p40__;
output            post_value_holder__p41__;
output            post_value_holder__p42__;
output            post_value_holder__p43__;
output            post_value_holder__p44__;
output            post_value_holder__p45__;
output            post_value_holder__p46__;
output            post_value_holder__p47__;
output            post_value_holder__p48__;
output            post_value_holder__p49__;
output            post_value_holder__p50__;
output            post_value_holder__p51__;
output            post_value_holder__p52__;
output            post_value_holder__p53__;
output            post_value_holder__p54__;
output            post_value_holder__p55__;
output            post_value_holder__p56__;
output            post_value_holder__p57__;
output            post_value_holder__p58__;
output            post_value_holder__p59__;
output            post_value_holder__p60__;
output            post_value_holder__p61__;
output            post_value_holder__p62__;
output            post_value_holder__p63__;
output            post_value_holder__p64__;
output            post_value_holder__p65__;
output            post_value_holder__p66__;
output            post_value_holder__p67__;
output            post_value_holder__p68__;
output            post_value_holder__p69__;
output            post_value_holder__p70__;
output            post_value_holder__p71__;
output            post_value_holder__p72__;
output            post_value_holder__p73__;
output            post_value_holder_overly_constrained__p153__;
output            post_value_holder_overly_constrained__p154__;
output            post_value_holder_overly_constrained__p155__;
output            post_value_holder_overly_constrained__p156__;
output            post_value_holder_overly_constrained__p157__;
output            post_value_holder_overly_constrained__p158__;
output            post_value_holder_overly_constrained__p159__;
output            post_value_holder_overly_constrained__p160__;
output            post_value_holder_overly_constrained__p161__;
output            post_value_holder_overly_constrained__p162__;
output            post_value_holder_overly_constrained__p163__;
output            post_value_holder_overly_constrained__p164__;
output            post_value_holder_overly_constrained__p165__;
output            post_value_holder_overly_constrained__p166__;
output            post_value_holder_overly_constrained__p167__;
output            post_value_holder_overly_constrained__p168__;
output            post_value_holder_overly_constrained__p169__;
output            post_value_holder_overly_constrained__p170__;
output            post_value_holder_overly_constrained__p171__;
output            post_value_holder_overly_constrained__p172__;
output            post_value_holder_overly_constrained__p173__;
output            post_value_holder_overly_constrained__p174__;
output            post_value_holder_overly_constrained__p175__;
output            post_value_holder_overly_constrained__p176__;
output            post_value_holder_overly_constrained__p177__;
output            post_value_holder_overly_constrained__p178__;
output            post_value_holder_overly_constrained__p179__;
output            post_value_holder_overly_constrained__p180__;
output            post_value_holder_overly_constrained__p181__;
output            post_value_holder_overly_constrained__p182__;
output            post_value_holder_overly_constrained__p183__;
output            post_value_holder_overly_constrained__p184__;
output            post_value_holder_overly_constrained__p185__;
output            post_value_holder_overly_constrained__p186__;
output            post_value_holder_overly_constrained__p187__;
output            post_value_holder_overly_constrained__p188__;
output            post_value_holder_overly_constrained__p189__;
output            post_value_holder_overly_constrained__p190__;
output            post_value_holder_triggered__p191__;
output            post_value_holder_triggered__p192__;
output            post_value_holder_triggered__p193__;
output            post_value_holder_triggered__p194__;
output            post_value_holder_triggered__p195__;
output            post_value_holder_triggered__p196__;
output            post_value_holder_triggered__p197__;
output            post_value_holder_triggered__p198__;
output            post_value_holder_triggered__p199__;
output            post_value_holder_triggered__p200__;
output            post_value_holder_triggered__p201__;
output            post_value_holder_triggered__p202__;
output            post_value_holder_triggered__p203__;
output            post_value_holder_triggered__p204__;
output            post_value_holder_triggered__p205__;
output            post_value_holder_triggered__p206__;
output            post_value_holder_triggered__p207__;
output            post_value_holder_triggered__p208__;
output            post_value_holder_triggered__p209__;
output            post_value_holder_triggered__p210__;
output            post_value_holder_triggered__p211__;
output            post_value_holder_triggered__p212__;
output            post_value_holder_triggered__p213__;
output            post_value_holder_triggered__p214__;
output            post_value_holder_triggered__p215__;
output            post_value_holder_triggered__p216__;
output            post_value_holder_triggered__p217__;
output            post_value_holder_triggered__p218__;
output            post_value_holder_triggered__p219__;
output            post_value_holder_triggered__p220__;
output            post_value_holder_triggered__p221__;
output            post_value_holder_triggered__p222__;
output            post_value_holder_triggered__p223__;
output            post_value_holder_triggered__p224__;
output            post_value_holder_triggered__p225__;
output            post_value_holder_triggered__p226__;
output            post_value_holder_triggered__p227__;
output            post_value_holder_triggered__p228__;
output            rfassumptions__p74__;
output            rfassumptions__p75__;
output            rfassumptions__p76__;
output            s2_enter;
output            s2_exit;
output            s3_enter;
output            s3_exit;
output            s4_enter;
output            variable_map_assert__p118__;
output            variable_map_assert__p119__;
output            variable_map_assert__p120__;
output            variable_map_assert__p121__;
output            variable_map_assert__p122__;
output            variable_map_assert__p123__;
output            variable_map_assert__p124__;
output            variable_map_assert__p125__;
output            variable_map_assert__p126__;
output            variable_map_assert__p127__;
output            variable_map_assert__p128__;
output            variable_map_assert__p129__;
output            variable_map_assert__p130__;
output            variable_map_assert__p131__;
output            variable_map_assert__p132__;
output            variable_map_assert__p133__;
output            variable_map_assert__p134__;
output            variable_map_assert__p135__;
output            variable_map_assert__p136__;
output            variable_map_assert__p137__;
output            variable_map_assert__p138__;
output            variable_map_assert__p139__;
output            variable_map_assert__p140__;
output            variable_map_assert__p141__;
output            variable_map_assert__p142__;
output            variable_map_assert__p143__;
output            variable_map_assert__p144__;
output            variable_map_assert__p145__;
output            variable_map_assert__p146__;
output            variable_map_assert__p147__;
output            variable_map_assert__p148__;
output            variable_map_assert__p149__;
output            variable_map_assert__p150__;
output            variable_map_assert__p151__;
output            variable_map_assert__p152__;
output            variable_map_assume___p100__;
output            variable_map_assume___p101__;
output            variable_map_assume___p102__;
output            variable_map_assume___p103__;
output            variable_map_assume___p104__;
output            variable_map_assume___p105__;
output            variable_map_assume___p106__;
output            variable_map_assume___p107__;
output            variable_map_assume___p108__;
output            variable_map_assume___p109__;
output            variable_map_assume___p110__;
output            variable_map_assume___p111__;
output            variable_map_assume___p112__;
output            variable_map_assume___p113__;
output            variable_map_assume___p114__;
output            variable_map_assume___p115__;
output            variable_map_assume___p116__;
output            variable_map_assume___p117__;
output            variable_map_assume___p77__;
output            variable_map_assume___p78__;
output            variable_map_assume___p79__;
output            variable_map_assume___p80__;
output            variable_map_assume___p81__;
output            variable_map_assume___p82__;
output            variable_map_assume___p83__;
output            variable_map_assume___p84__;
output            variable_map_assume___p85__;
output            variable_map_assume___p86__;
output            variable_map_assume___p87__;
output            variable_map_assume___p88__;
output            variable_map_assume___p89__;
output            variable_map_assume___p90__;
output            variable_map_assume___p91__;
output            variable_map_assume___p92__;
output            variable_map_assume___p93__;
output            variable_map_assume___p94__;
output            variable_map_assume___p95__;
output            variable_map_assume___p96__;
output            variable_map_assume___p97__;
output            variable_map_assume___p98__;
output            variable_map_assume___p99__;
output reg      [7:0] __CYCLE_CNT__;
output reg            __START__;
output reg            __STARTED__;
output reg            __ENDED__;
output reg            __2ndENDED__;
output reg            __RESETED__;
output reg     [31:0] __auxvar10__recorder;
output reg     [31:0] __auxvar10__recorder_sn_vhold;
output reg            __auxvar10__recorder_sn_condmet;
output reg     [31:0] __auxvar11__recorder;
output reg     [31:0] __auxvar11__recorder_sn_vhold;
output reg            __auxvar11__recorder_sn_condmet;
output reg     [31:0] __auxvar12__recorder;
output reg     [31:0] __auxvar12__recorder_sn_vhold;
output reg            __auxvar12__recorder_sn_condmet;
output reg     [31:0] __auxvar13__recorder;
output reg     [31:0] __auxvar13__recorder_sn_vhold;
output reg            __auxvar13__recorder_sn_condmet;
output reg     [31:0] __auxvar14__recorder;
output reg     [31:0] __auxvar14__recorder_sn_vhold;
output reg            __auxvar14__recorder_sn_condmet;
output reg     [31:0] __auxvar15__recorder;
output reg     [31:0] __auxvar15__recorder_sn_vhold;
output reg            __auxvar15__recorder_sn_condmet;
output reg     [31:0] __auxvar16__recorder;
output reg     [31:0] __auxvar16__recorder_sn_vhold;
output reg            __auxvar16__recorder_sn_condmet;
output reg     [31:0] __auxvar17__recorder;
output reg     [31:0] __auxvar17__recorder_sn_vhold;
output reg            __auxvar17__recorder_sn_condmet;
output reg     [31:0] __auxvar18__recorder;
output reg     [31:0] __auxvar18__recorder_sn_vhold;
output reg            __auxvar18__recorder_sn_condmet;
output reg     [31:0] __auxvar19__recorder;
output reg     [31:0] __auxvar19__recorder_sn_vhold;
output reg            __auxvar19__recorder_sn_condmet;
output reg     [31:0] __auxvar1__recorder;
output reg     [31:0] __auxvar1__recorder_sn_vhold;
output reg            __auxvar1__recorder_sn_condmet;
output reg     [31:0] __auxvar20__recorder;
output reg     [31:0] __auxvar20__recorder_sn_vhold;
output reg            __auxvar20__recorder_sn_condmet;
output reg     [31:0] __auxvar21__recorder;
output reg     [31:0] __auxvar21__recorder_sn_vhold;
output reg            __auxvar21__recorder_sn_condmet;
output reg     [31:0] __auxvar22__recorder;
output reg     [31:0] __auxvar22__recorder_sn_vhold;
output reg            __auxvar22__recorder_sn_condmet;
output reg     [31:0] __auxvar23__recorder;
output reg     [31:0] __auxvar23__recorder_sn_vhold;
output reg            __auxvar23__recorder_sn_condmet;
output reg     [31:0] __auxvar24__recorder;
output reg     [31:0] __auxvar24__recorder_sn_vhold;
output reg            __auxvar24__recorder_sn_condmet;
output reg     [31:0] __auxvar25__recorder;
output reg     [31:0] __auxvar25__recorder_sn_vhold;
output reg            __auxvar25__recorder_sn_condmet;
output reg     [31:0] __auxvar26__recorder;
output reg     [31:0] __auxvar26__recorder_sn_vhold;
output reg            __auxvar26__recorder_sn_condmet;
output reg     [31:0] __auxvar27__recorder;
output reg     [31:0] __auxvar27__recorder_sn_vhold;
output reg            __auxvar27__recorder_sn_condmet;
output reg     [31:0] __auxvar28__recorder;
output reg     [31:0] __auxvar28__recorder_sn_vhold;
output reg            __auxvar28__recorder_sn_condmet;
output reg     [31:0] __auxvar29__recorder;
output reg     [31:0] __auxvar29__recorder_sn_vhold;
output reg            __auxvar29__recorder_sn_condmet;
output reg     [31:0] __auxvar2__recorder;
output reg     [31:0] __auxvar2__recorder_sn_vhold;
output reg            __auxvar2__recorder_sn_condmet;
output reg     [31:0] __auxvar30__recorder;
output reg     [31:0] __auxvar30__recorder_sn_vhold;
output reg            __auxvar30__recorder_sn_condmet;
output reg     [31:0] __auxvar31__recorder;
output reg     [31:0] __auxvar31__recorder_sn_vhold;
output reg            __auxvar31__recorder_sn_condmet;
output reg     [31:0] __auxvar32__recorder;
output reg     [31:0] __auxvar32__recorder_sn_vhold;
output reg            __auxvar32__recorder_sn_condmet;
output reg     [31:0] __auxvar33__recorder;
output reg     [31:0] __auxvar33__recorder_sn_vhold;
output reg            __auxvar33__recorder_sn_condmet;
output reg            __auxvar34__recorder;
output reg            __auxvar34__recorder_sn_vhold;
output reg            __auxvar34__recorder_sn_condmet;
output reg      [2:0] __auxvar35__recorder;
output reg      [2:0] __auxvar35__recorder_sn_vhold;
output reg            __auxvar35__recorder_sn_condmet;
output reg            __auxvar36__recorder;
output reg            __auxvar36__recorder_sn_vhold;
output reg            __auxvar36__recorder_sn_condmet;
output reg     [31:0] __auxvar37__recorder;
output reg     [31:0] __auxvar37__recorder_sn_vhold;
output reg            __auxvar37__recorder_sn_condmet;
output reg     [31:0] __auxvar38__recorder;
output reg     [31:0] __auxvar38__recorder_sn_vhold;
output reg            __auxvar38__recorder_sn_condmet;
output reg     [31:0] __auxvar3__recorder;
output reg     [31:0] __auxvar3__recorder_sn_vhold;
output reg            __auxvar3__recorder_sn_condmet;
output reg     [31:0] __auxvar4__recorder;
output reg     [31:0] __auxvar4__recorder_sn_vhold;
output reg            __auxvar4__recorder_sn_condmet;
output reg     [31:0] __auxvar5__recorder;
output reg     [31:0] __auxvar5__recorder_sn_vhold;
output reg            __auxvar5__recorder_sn_condmet;
output reg     [31:0] __auxvar6__recorder;
output reg     [31:0] __auxvar6__recorder_sn_vhold;
output reg            __auxvar6__recorder_sn_condmet;
output reg     [31:0] __auxvar7__recorder;
output reg     [31:0] __auxvar7__recorder_sn_vhold;
output reg            __auxvar7__recorder_sn_condmet;
output reg     [31:0] __auxvar8__recorder;
output reg     [31:0] __auxvar8__recorder_sn_vhold;
output reg            __auxvar8__recorder_sn_condmet;
output reg     [31:0] __auxvar9__recorder;
output reg     [31:0] __auxvar9__recorder_sn_vhold;
output reg            __auxvar9__recorder_sn_condmet;
output reg            __auxvar0__delay_d_1;
output reg            monitor_s1_already;
output reg            monitor_s2;
output reg            monitor_s3;
output reg            monitor_s4;
 wire            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__csr_regfile__DOT__rg_nmi;
 wire            RTL__DOT__csr_regfile__DOT__rg_state;
 wire            RTL__DOT__f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
 wire     [31:0] RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
 wire            RTL__DOT__near_mem$EN_dmem_req;
 wire            RTL__DOT__near_mem$dmem_exc;
 wire     [31:0] RTL__DOT__near_mem$dmem_req_addr;
 wire      [2:0] RTL__DOT__near_mem$dmem_req_f3;
 wire            RTL__DOT__near_mem$dmem_req_op;
 wire     [63:0] RTL__DOT__near_mem$dmem_req_store_value;
 wire     [63:0] RTL__DOT__near_mem$dmem_word64;
 wire     [31:0] RTL__DOT__near_mem$imem_instr;
 wire     [31:0] RTL__DOT__near_mem$imem_pc;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
 wire     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
 wire     [31:0] RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
 wire            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
 wire            RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
 wire      [1:0] RTL__DOT__rg_cur_priv;
 wire            RTL__DOT__rg_retiring$EN;
 wire            RTL__DOT__rg_run_on_reset;
 wire      [3:0] RTL__DOT__rg_state;
 wire     [31:0] RTL__DOT__rg_trap_instr;
 wire            RTL__DOT__s1_to_s2$D_IN;
 wire            RTL__DOT__s1_to_s2$EN;
 wire            RTL__DOT__s2_to_s3$D_IN;
 wire            RTL__DOT__s2_to_s3$EN;
 wire            RTL__DOT__s3_deq$D_IN;
 wire            RTL__DOT__s3_deq$EN;
 wire            RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__stage1_rg_full;
 wire            RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__stage2_rg_full;
 wire    [168:0] RTL__DOT__stage2_rg_stage2;
 wire            RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
 wire            RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
 wire            RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
 wire            RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
 wire            RTL__DOT__stage3_rg_full;
wire            __2ndIEND__;
 wire            __EDCOND__;
 wire            __IEND__;
 wire     [31:0] __ILA_I_inst;
 wire     [31:0] __ILA_SO_load_addr;
 wire     [31:0] __ILA_SO_load_data;
 wire            __ILA_SO_load_en;
 wire      [2:0] __ILA_SO_load_size;
 wire     [31:0] __ILA_SO_pc;
 wire     [31:0] __ILA_SO_store_addr;
 wire     [31:0] __ILA_SO_store_data;
 wire            __ILA_SO_store_en;
 wire      [2:0] __ILA_SO_store_size;
 wire     [31:0] __ILA_SO_x0;
 wire     [31:0] __ILA_SO_x1;
 wire     [31:0] __ILA_SO_x10;
 wire     [31:0] __ILA_SO_x11;
 wire     [31:0] __ILA_SO_x12;
 wire     [31:0] __ILA_SO_x13;
 wire     [31:0] __ILA_SO_x14;
 wire     [31:0] __ILA_SO_x15;
 wire     [31:0] __ILA_SO_x16;
 wire     [31:0] __ILA_SO_x17;
 wire     [31:0] __ILA_SO_x18;
 wire     [31:0] __ILA_SO_x19;
 wire     [31:0] __ILA_SO_x2;
 wire     [31:0] __ILA_SO_x20;
 wire     [31:0] __ILA_SO_x21;
 wire     [31:0] __ILA_SO_x22;
 wire     [31:0] __ILA_SO_x23;
 wire     [31:0] __ILA_SO_x24;
 wire     [31:0] __ILA_SO_x25;
 wire     [31:0] __ILA_SO_x26;
 wire     [31:0] __ILA_SO_x27;
 wire     [31:0] __ILA_SO_x28;
 wire     [31:0] __ILA_SO_x29;
 wire     [31:0] __ILA_SO_x3;
 wire     [31:0] __ILA_SO_x30;
 wire     [31:0] __ILA_SO_x31;
 wire     [31:0] __ILA_SO_x4;
 wire     [31:0] __ILA_SO_x5;
 wire     [31:0] __ILA_SO_x6;
 wire     [31:0] __ILA_SO_x7;
 wire     [31:0] __ILA_SO_x8;
 wire     [31:0] __ILA_SO_x9;
 wire            __ILA_riscv_decode_of_ADD__;
 wire            __ILA_riscv_valid__;
 wire            __ISSUE__;
 wire            __VLG_II_m_external_interrupt_req_set_not_clear;
 wire            __VLG_II_nmi_req_set_not_clear;
 wire            __VLG_II_s_external_interrupt_req_set_not_clear;
 wire            __VLG_II_software_interrupt_req_set_not_clear;
 wire            __VLG_II_timer_interrupt_req_set_not_clear;
 wire            __VLG_I_EN_hart0_server_reset_request_put;
 wire            __VLG_I_EN_hart0_server_reset_response_get;
 wire            __VLG_I_EN_set_verbosity;
 wire            __VLG_I_dmem_master_arready;
 wire            __VLG_I_dmem_master_awready;
 wire      [3:0] __VLG_I_dmem_master_bid;
 wire      [1:0] __VLG_I_dmem_master_bresp;
 wire            __VLG_I_dmem_master_bvalid;
 wire     [63:0] __VLG_I_dmem_master_rdata;
 wire      [3:0] __VLG_I_dmem_master_rid;
 wire            __VLG_I_dmem_master_rlast;
 wire      [1:0] __VLG_I_dmem_master_rresp;
 wire            __VLG_I_dmem_master_rvalid;
 wire            __VLG_I_dmem_master_wready;
 wire            __VLG_I_hart0_server_reset_request_put;
 wire            __VLG_I_imem_master_arready;
 wire            __VLG_I_imem_master_awready;
 wire      [3:0] __VLG_I_imem_master_bid;
 wire      [1:0] __VLG_I_imem_master_bresp;
 wire            __VLG_I_imem_master_bvalid;
 wire     [63:0] __VLG_I_imem_master_rdata;
 wire      [3:0] __VLG_I_imem_master_rid;
 wire            __VLG_I_imem_master_rlast;
 wire      [1:0] __VLG_I_imem_master_rresp;
 wire            __VLG_I_imem_master_rvalid;
 wire            __VLG_I_imem_master_wready;
 wire     [63:0] __VLG_I_set_verbosity_logdelay;
 wire      [3:0] __VLG_I_set_verbosity_verbosity;
 wire            __VLG_O_RDY_hart0_server_reset_request_put;
 wire            __VLG_O_RDY_hart0_server_reset_response_get;
 wire            __VLG_O_RDY_set_verbosity;
 wire     [63:0] __VLG_O_dmem_master_araddr;
 wire      [1:0] __VLG_O_dmem_master_arburst;
 wire      [3:0] __VLG_O_dmem_master_arcache;
 wire      [3:0] __VLG_O_dmem_master_arid;
 wire      [7:0] __VLG_O_dmem_master_arlen;
 wire            __VLG_O_dmem_master_arlock;
 wire      [2:0] __VLG_O_dmem_master_arprot;
 wire      [3:0] __VLG_O_dmem_master_arqos;
 wire      [3:0] __VLG_O_dmem_master_arregion;
 wire      [2:0] __VLG_O_dmem_master_arsize;
 wire            __VLG_O_dmem_master_arvalid;
 wire     [63:0] __VLG_O_dmem_master_awaddr;
 wire      [1:0] __VLG_O_dmem_master_awburst;
 wire      [3:0] __VLG_O_dmem_master_awcache;
 wire      [3:0] __VLG_O_dmem_master_awid;
 wire      [7:0] __VLG_O_dmem_master_awlen;
 wire            __VLG_O_dmem_master_awlock;
 wire      [2:0] __VLG_O_dmem_master_awprot;
 wire      [3:0] __VLG_O_dmem_master_awqos;
 wire      [3:0] __VLG_O_dmem_master_awregion;
 wire      [2:0] __VLG_O_dmem_master_awsize;
 wire            __VLG_O_dmem_master_awvalid;
 wire            __VLG_O_dmem_master_bready;
 wire            __VLG_O_dmem_master_rready;
 wire     [63:0] __VLG_O_dmem_master_wdata;
 wire            __VLG_O_dmem_master_wlast;
 wire      [7:0] __VLG_O_dmem_master_wstrb;
 wire            __VLG_O_dmem_master_wvalid;
 wire            __VLG_O_hart0_server_reset_response_get;
 wire     [63:0] __VLG_O_imem_master_araddr;
 wire      [1:0] __VLG_O_imem_master_arburst;
 wire      [3:0] __VLG_O_imem_master_arcache;
 wire      [3:0] __VLG_O_imem_master_arid;
 wire      [7:0] __VLG_O_imem_master_arlen;
 wire            __VLG_O_imem_master_arlock;
 wire      [2:0] __VLG_O_imem_master_arprot;
 wire      [3:0] __VLG_O_imem_master_arqos;
 wire      [3:0] __VLG_O_imem_master_arregion;
 wire      [2:0] __VLG_O_imem_master_arsize;
 wire            __VLG_O_imem_master_arvalid;
 wire     [63:0] __VLG_O_imem_master_awaddr;
 wire      [1:0] __VLG_O_imem_master_awburst;
 wire      [3:0] __VLG_O_imem_master_awcache;
 wire      [3:0] __VLG_O_imem_master_awid;
 wire      [7:0] __VLG_O_imem_master_awlen;
 wire            __VLG_O_imem_master_awlock;
 wire      [2:0] __VLG_O_imem_master_awprot;
 wire      [3:0] __VLG_O_imem_master_awqos;
 wire      [3:0] __VLG_O_imem_master_awregion;
 wire      [2:0] __VLG_O_imem_master_awsize;
 wire            __VLG_O_imem_master_awvalid;
 wire            __VLG_O_imem_master_bready;
 wire            __VLG_O_imem_master_rready;
 wire     [63:0] __VLG_O_imem_master_wdata;
 wire            __VLG_O_imem_master_wlast;
 wire      [7:0] __VLG_O_imem_master_wstrb;
 wire            __VLG_O_imem_master_wvalid;
wire     [31:0] ____auxvar10__recorder_init__;
wire     [31:0] ____auxvar11__recorder_init__;
wire     [31:0] ____auxvar12__recorder_init__;
wire     [31:0] ____auxvar13__recorder_init__;
wire     [31:0] ____auxvar14__recorder_init__;
wire     [31:0] ____auxvar15__recorder_init__;
wire     [31:0] ____auxvar16__recorder_init__;
wire     [31:0] ____auxvar17__recorder_init__;
wire     [31:0] ____auxvar18__recorder_init__;
wire     [31:0] ____auxvar19__recorder_init__;
wire     [31:0] ____auxvar1__recorder_init__;
wire     [31:0] ____auxvar20__recorder_init__;
wire     [31:0] ____auxvar21__recorder_init__;
wire     [31:0] ____auxvar22__recorder_init__;
wire     [31:0] ____auxvar23__recorder_init__;
wire     [31:0] ____auxvar24__recorder_init__;
wire     [31:0] ____auxvar25__recorder_init__;
wire     [31:0] ____auxvar26__recorder_init__;
wire     [31:0] ____auxvar27__recorder_init__;
wire     [31:0] ____auxvar28__recorder_init__;
wire     [31:0] ____auxvar29__recorder_init__;
wire     [31:0] ____auxvar2__recorder_init__;
wire     [31:0] ____auxvar30__recorder_init__;
wire     [31:0] ____auxvar31__recorder_init__;
wire     [31:0] ____auxvar32__recorder_init__;
wire     [31:0] ____auxvar33__recorder_init__;
wire            ____auxvar34__recorder_init__;
wire      [2:0] ____auxvar35__recorder_init__;
wire            ____auxvar36__recorder_init__;
wire     [31:0] ____auxvar37__recorder_init__;
wire     [31:0] ____auxvar38__recorder_init__;
wire     [31:0] ____auxvar3__recorder_init__;
wire     [31:0] ____auxvar4__recorder_init__;
wire     [31:0] ____auxvar5__recorder_init__;
wire     [31:0] ____auxvar6__recorder_init__;
wire     [31:0] ____auxvar7__recorder_init__;
wire     [31:0] ____auxvar8__recorder_init__;
wire     [31:0] ____auxvar9__recorder_init__;
 wire            __all_assert_wire__;
 wire            __all_assume_wire__;
wire            __auxvar0__delay;
 wire            __auxvar0__delay_d_0;
wire            __auxvar10__recorder_sn_cond;
wire     [31:0] __auxvar10__recorder_sn_value;
wire            __auxvar11__recorder_sn_cond;
wire     [31:0] __auxvar11__recorder_sn_value;
wire            __auxvar12__recorder_sn_cond;
wire     [31:0] __auxvar12__recorder_sn_value;
wire            __auxvar13__recorder_sn_cond;
wire     [31:0] __auxvar13__recorder_sn_value;
wire            __auxvar14__recorder_sn_cond;
wire     [31:0] __auxvar14__recorder_sn_value;
wire            __auxvar15__recorder_sn_cond;
wire     [31:0] __auxvar15__recorder_sn_value;
wire            __auxvar16__recorder_sn_cond;
wire     [31:0] __auxvar16__recorder_sn_value;
wire            __auxvar17__recorder_sn_cond;
wire     [31:0] __auxvar17__recorder_sn_value;
wire            __auxvar18__recorder_sn_cond;
wire     [31:0] __auxvar18__recorder_sn_value;
wire            __auxvar19__recorder_sn_cond;
wire     [31:0] __auxvar19__recorder_sn_value;
wire            __auxvar1__recorder_sn_cond;
wire     [31:0] __auxvar1__recorder_sn_value;
wire            __auxvar20__recorder_sn_cond;
wire     [31:0] __auxvar20__recorder_sn_value;
wire            __auxvar21__recorder_sn_cond;
wire     [31:0] __auxvar21__recorder_sn_value;
wire            __auxvar22__recorder_sn_cond;
wire     [31:0] __auxvar22__recorder_sn_value;
wire            __auxvar23__recorder_sn_cond;
wire     [31:0] __auxvar23__recorder_sn_value;
wire            __auxvar24__recorder_sn_cond;
wire     [31:0] __auxvar24__recorder_sn_value;
wire            __auxvar25__recorder_sn_cond;
wire     [31:0] __auxvar25__recorder_sn_value;
wire            __auxvar26__recorder_sn_cond;
wire     [31:0] __auxvar26__recorder_sn_value;
wire            __auxvar27__recorder_sn_cond;
wire     [31:0] __auxvar27__recorder_sn_value;
wire            __auxvar28__recorder_sn_cond;
wire     [31:0] __auxvar28__recorder_sn_value;
wire            __auxvar29__recorder_sn_cond;
wire     [31:0] __auxvar29__recorder_sn_value;
wire            __auxvar2__recorder_sn_cond;
wire     [31:0] __auxvar2__recorder_sn_value;
wire            __auxvar30__recorder_sn_cond;
wire     [31:0] __auxvar30__recorder_sn_value;
wire            __auxvar31__recorder_sn_cond;
wire     [31:0] __auxvar31__recorder_sn_value;
wire            __auxvar32__recorder_sn_cond;
wire     [31:0] __auxvar32__recorder_sn_value;
wire            __auxvar33__recorder_sn_cond;
wire     [31:0] __auxvar33__recorder_sn_value;
wire            __auxvar34__recorder_sn_cond;
wire            __auxvar34__recorder_sn_value;
wire            __auxvar35__recorder_sn_cond;
wire      [2:0] __auxvar35__recorder_sn_value;
wire            __auxvar36__recorder_sn_cond;
wire            __auxvar36__recorder_sn_value;
wire            __auxvar37__recorder_sn_cond;
wire     [31:0] __auxvar37__recorder_sn_value;
wire            __auxvar38__recorder_sn_cond;
wire     [31:0] __auxvar38__recorder_sn_value;
wire            __auxvar3__recorder_sn_cond;
wire     [31:0] __auxvar3__recorder_sn_value;
wire            __auxvar4__recorder_sn_cond;
wire     [31:0] __auxvar4__recorder_sn_value;
wire            __auxvar5__recorder_sn_cond;
wire     [31:0] __auxvar5__recorder_sn_value;
wire            __auxvar6__recorder_sn_cond;
wire     [31:0] __auxvar6__recorder_sn_value;
wire            __auxvar7__recorder_sn_cond;
wire     [31:0] __auxvar7__recorder_sn_value;
wire            __auxvar8__recorder_sn_cond;
wire     [31:0] __auxvar8__recorder_sn_value;
wire            __auxvar9__recorder_sn_cond;
wire     [31:0] __auxvar9__recorder_sn_value;
 wire            __sanitycheck_wire__;
wire            clk;
 wire            dummy_reset;
wire            end_of_pipeline;
wire            input_map_assume___p0__;
wire            invariant_assume__p10__;
wire            invariant_assume__p11__;
wire            invariant_assume__p12__;
wire            invariant_assume__p13__;
wire            invariant_assume__p14__;
wire            invariant_assume__p15__;
wire            invariant_assume__p16__;
wire            invariant_assume__p17__;
wire            invariant_assume__p18__;
wire            invariant_assume__p19__;
wire            invariant_assume__p1__;
wire            invariant_assume__p20__;
wire            invariant_assume__p21__;
wire            invariant_assume__p22__;
wire            invariant_assume__p23__;
wire            invariant_assume__p24__;
wire            invariant_assume__p25__;
wire            invariant_assume__p26__;
wire            invariant_assume__p27__;
wire            invariant_assume__p28__;
wire            invariant_assume__p29__;
wire            invariant_assume__p2__;
wire            invariant_assume__p30__;
wire            invariant_assume__p31__;
wire            invariant_assume__p32__;
wire            invariant_assume__p3__;
wire            invariant_assume__p4__;
wire            invariant_assume__p5__;
wire            invariant_assume__p6__;
wire            invariant_assume__p7__;
wire            invariant_assume__p8__;
wire            invariant_assume__p9__;
wire            issue_decode__p33__;
wire            issue_valid__p34__;
 wire     [31:0] mem_req_addr;
 wire            mem_req_en;
 wire      [2:0] mem_req_funct3;
 wire            mem_req_op;
 wire     [31:0] mem_req_rd_data;
 wire     [31:0] mem_req_wd_data;
wire            monitor_s1;
 wire            monitor_s1_already_enter_cond;
 wire            monitor_s1_already_exit_cond;
 wire            monitor_s2_enter_cond;
 wire            monitor_s2_exit_cond;
 wire            monitor_s3_enter_cond;
 wire            monitor_s3_exit_cond;
 wire            monitor_s4_enter_cond;
 wire            monitor_s4_exit_cond;
wire            noreset__p35__;
wire            post_value_holder__p36__;
wire            post_value_holder__p37__;
wire            post_value_holder__p38__;
wire            post_value_holder__p39__;
wire            post_value_holder__p40__;
wire            post_value_holder__p41__;
wire            post_value_holder__p42__;
wire            post_value_holder__p43__;
wire            post_value_holder__p44__;
wire            post_value_holder__p45__;
wire            post_value_holder__p46__;
wire            post_value_holder__p47__;
wire            post_value_holder__p48__;
wire            post_value_holder__p49__;
wire            post_value_holder__p50__;
wire            post_value_holder__p51__;
wire            post_value_holder__p52__;
wire            post_value_holder__p53__;
wire            post_value_holder__p54__;
wire            post_value_holder__p55__;
wire            post_value_holder__p56__;
wire            post_value_holder__p57__;
wire            post_value_holder__p58__;
wire            post_value_holder__p59__;
wire            post_value_holder__p60__;
wire            post_value_holder__p61__;
wire            post_value_holder__p62__;
wire            post_value_holder__p63__;
wire            post_value_holder__p64__;
wire            post_value_holder__p65__;
wire            post_value_holder__p66__;
wire            post_value_holder__p67__;
wire            post_value_holder__p68__;
wire            post_value_holder__p69__;
wire            post_value_holder__p70__;
wire            post_value_holder__p71__;
wire            post_value_holder__p72__;
wire            post_value_holder__p73__;
wire            post_value_holder_overly_constrained__p153__;
wire            post_value_holder_overly_constrained__p154__;
wire            post_value_holder_overly_constrained__p155__;
wire            post_value_holder_overly_constrained__p156__;
wire            post_value_holder_overly_constrained__p157__;
wire            post_value_holder_overly_constrained__p158__;
wire            post_value_holder_overly_constrained__p159__;
wire            post_value_holder_overly_constrained__p160__;
wire            post_value_holder_overly_constrained__p161__;
wire            post_value_holder_overly_constrained__p162__;
wire            post_value_holder_overly_constrained__p163__;
wire            post_value_holder_overly_constrained__p164__;
wire            post_value_holder_overly_constrained__p165__;
wire            post_value_holder_overly_constrained__p166__;
wire            post_value_holder_overly_constrained__p167__;
wire            post_value_holder_overly_constrained__p168__;
wire            post_value_holder_overly_constrained__p169__;
wire            post_value_holder_overly_constrained__p170__;
wire            post_value_holder_overly_constrained__p171__;
wire            post_value_holder_overly_constrained__p172__;
wire            post_value_holder_overly_constrained__p173__;
wire            post_value_holder_overly_constrained__p174__;
wire            post_value_holder_overly_constrained__p175__;
wire            post_value_holder_overly_constrained__p176__;
wire            post_value_holder_overly_constrained__p177__;
wire            post_value_holder_overly_constrained__p178__;
wire            post_value_holder_overly_constrained__p179__;
wire            post_value_holder_overly_constrained__p180__;
wire            post_value_holder_overly_constrained__p181__;
wire            post_value_holder_overly_constrained__p182__;
wire            post_value_holder_overly_constrained__p183__;
wire            post_value_holder_overly_constrained__p184__;
wire            post_value_holder_overly_constrained__p185__;
wire            post_value_holder_overly_constrained__p186__;
wire            post_value_holder_overly_constrained__p187__;
wire            post_value_holder_overly_constrained__p188__;
wire            post_value_holder_overly_constrained__p189__;
wire            post_value_holder_overly_constrained__p190__;
wire            post_value_holder_triggered__p191__;
wire            post_value_holder_triggered__p192__;
wire            post_value_holder_triggered__p193__;
wire            post_value_holder_triggered__p194__;
wire            post_value_holder_triggered__p195__;
wire            post_value_holder_triggered__p196__;
wire            post_value_holder_triggered__p197__;
wire            post_value_holder_triggered__p198__;
wire            post_value_holder_triggered__p199__;
wire            post_value_holder_triggered__p200__;
wire            post_value_holder_triggered__p201__;
wire            post_value_holder_triggered__p202__;
wire            post_value_holder_triggered__p203__;
wire            post_value_holder_triggered__p204__;
wire            post_value_holder_triggered__p205__;
wire            post_value_holder_triggered__p206__;
wire            post_value_holder_triggered__p207__;
wire            post_value_holder_triggered__p208__;
wire            post_value_holder_triggered__p209__;
wire            post_value_holder_triggered__p210__;
wire            post_value_holder_triggered__p211__;
wire            post_value_holder_triggered__p212__;
wire            post_value_holder_triggered__p213__;
wire            post_value_holder_triggered__p214__;
wire            post_value_holder_triggered__p215__;
wire            post_value_holder_triggered__p216__;
wire            post_value_holder_triggered__p217__;
wire            post_value_holder_triggered__p218__;
wire            post_value_holder_triggered__p219__;
wire            post_value_holder_triggered__p220__;
wire            post_value_holder_triggered__p221__;
wire            post_value_holder_triggered__p222__;
wire            post_value_holder_triggered__p223__;
wire            post_value_holder_triggered__p224__;
wire            post_value_holder_triggered__p225__;
wire            post_value_holder_triggered__p226__;
wire            post_value_holder_triggered__p227__;
wire            post_value_holder_triggered__p228__;
wire            rfassumptions__p74__;
wire            rfassumptions__p75__;
wire            rfassumptions__p76__;
wire            rst;
wire            s2_enter;
wire            s2_exit;
wire            s3_enter;
wire            s3_exit;
wire            s4_enter;
wire            variable_map_assert__p118__;
wire            variable_map_assert__p119__;
wire            variable_map_assert__p120__;
wire            variable_map_assert__p121__;
wire            variable_map_assert__p122__;
wire            variable_map_assert__p123__;
wire            variable_map_assert__p124__;
wire            variable_map_assert__p125__;
wire            variable_map_assert__p126__;
wire            variable_map_assert__p127__;
wire            variable_map_assert__p128__;
wire            variable_map_assert__p129__;
wire            variable_map_assert__p130__;
wire            variable_map_assert__p131__;
wire            variable_map_assert__p132__;
wire            variable_map_assert__p133__;
wire            variable_map_assert__p134__;
wire            variable_map_assert__p135__;
wire            variable_map_assert__p136__;
wire            variable_map_assert__p137__;
wire            variable_map_assert__p138__;
wire            variable_map_assert__p139__;
wire            variable_map_assert__p140__;
wire            variable_map_assert__p141__;
wire            variable_map_assert__p142__;
wire            variable_map_assert__p143__;
wire            variable_map_assert__p144__;
wire            variable_map_assert__p145__;
wire            variable_map_assert__p146__;
wire            variable_map_assert__p147__;
wire            variable_map_assert__p148__;
wire            variable_map_assert__p149__;
wire            variable_map_assert__p150__;
wire            variable_map_assert__p151__;
wire            variable_map_assert__p152__;
wire            variable_map_assume___p100__;
wire            variable_map_assume___p101__;
wire            variable_map_assume___p102__;
wire            variable_map_assume___p103__;
wire            variable_map_assume___p104__;
wire            variable_map_assume___p105__;
wire            variable_map_assume___p106__;
wire            variable_map_assume___p107__;
wire            variable_map_assume___p108__;
wire            variable_map_assume___p109__;
wire            variable_map_assume___p110__;
wire            variable_map_assume___p111__;
wire            variable_map_assume___p112__;
wire            variable_map_assume___p113__;
wire            variable_map_assume___p114__;
wire            variable_map_assume___p115__;
wire            variable_map_assume___p116__;
wire            variable_map_assume___p117__;
wire            variable_map_assume___p77__;
wire            variable_map_assume___p78__;
wire            variable_map_assume___p79__;
wire            variable_map_assume___p80__;
wire            variable_map_assume___p81__;
wire            variable_map_assume___p82__;
wire            variable_map_assume___p83__;
wire            variable_map_assume___p84__;
wire            variable_map_assume___p85__;
wire            variable_map_assume___p86__;
wire            variable_map_assume___p87__;
wire            variable_map_assume___p88__;
wire            variable_map_assume___p89__;
wire            variable_map_assume___p90__;
wire            variable_map_assume___p91__;
wire            variable_map_assume___p92__;
wire            variable_map_assume___p93__;
wire            variable_map_assume___p94__;
wire            variable_map_assume___p95__;
wire            variable_map_assume___p96__;
wire            variable_map_assume___p97__;
wire            variable_map_assume___p98__;
wire            variable_map_assume___p99__;
always @(posedge clk) begin
if (rst) __CYCLE_CNT__ <= 0;
else if ( ( __START__ || __STARTED__ ) &&  __CYCLE_CNT__ < 137) __CYCLE_CNT__ <= __CYCLE_CNT__ + 1;
end
always @(posedge clk) begin
if (__ISSUE__ && !__START__ && !__STARTED__) __START__ <= 1;
else if (__START__ || __STARTED__) __START__ <= 0;
end
always @(posedge clk) begin
if (rst) __STARTED__ <= 0;
else if (__START__) __STARTED__ <= 1;
end
always @(posedge clk) begin
if (rst) __ENDED__ <= 0;
else if (__IEND__) __ENDED__ <= 1;
end
always @(posedge clk) begin
if (rst) __2ndENDED__ <= 1'b0;
else if (__ENDED__ && __EDCOND__ && ~__2ndENDED__)  __2ndENDED__ <= 1'b1; end
assign __2ndIEND__ = __ENDED__ && __EDCOND__ && ~__2ndENDED__ ;
always @(posedge clk) begin
if (rst) __RESETED__ <= 1;
end
assign __auxvar0__delay = __auxvar0__delay_d_1 ;
assign monitor_s1_already_exit_cond = 1'b0 ;
assign monitor_s4_exit_cond = 1'b0 ;
    reg[31:0] ILA___pc;
    reg ILA___load_en;
    reg[31:0] ILA___load_addr;
    reg[2:0] ILA___load_size;
    reg[31:0] ILA___load_data;
    reg ILA___store_en;
    reg[31:0] ILA___store_addr;
    reg[2:0] ILA___store_size;
    reg[31:0] ILA___store_data;
    reg[31:0] ILA___x0;
    reg[31:0] ILA___x1;
    reg[31:0] ILA___x2;
    reg[31:0] ILA___x3;
    reg[31:0] ILA___x4;
    reg[31:0] ILA___x5;
    reg[31:0] ILA___x6;
    reg[31:0] ILA___x7;
    reg[31:0] ILA___x8;
    reg[31:0] ILA___x9;
    reg[31:0] ILA___x10;
    reg[31:0] ILA___x11;
    reg[31:0] ILA___x12;
    reg[31:0] ILA___x13;
    reg[31:0] ILA___x14;
    reg[31:0] ILA___x15;
    reg[31:0] ILA___x16;
    reg[31:0] ILA___x17;
    reg[31:0] ILA___x18;
    reg[31:0] ILA___x19;
    reg[31:0] ILA___x20;
    reg[31:0] ILA___x21;
    reg[31:0] ILA___x22;
    reg[31:0] ILA___x23;
    reg[31:0] ILA___x24;
    reg[31:0] ILA___x25;
    reg[31:0] ILA___x26;
    reg[31:0] ILA___x27;
    reg[31:0] ILA___x28;
    reg[31:0] ILA___x29;
    reg[31:0] ILA___x30;
    reg[31:0] ILA___x31;
    reg[7:0] ILA_____COUNTER_start__n11;

    wire ILA_____ILA_riscv_decode_of_ADD__ ; 
    wire ILA_____ILA_riscv_valid__ ; 
    wire ILA_____START__ ; 
    wire ILA___bv_1_0_n14 ; 
    wire[31:0] ILA___bv_32_0_n15 ; 
    wire[31:0] ILA___bv_32_4_n12 ; 
    wire[2:0] ILA___bv_3_0_n4 ; 
    wire[4:0] ILA___bv_5_10_n62 ; 
    wire[4:0] ILA___bv_5_11_n60 ; 
    wire[4:0] ILA___bv_5_12_n58 ; 
    wire[4:0] ILA___bv_5_13_n56 ; 
    wire[4:0] ILA___bv_5_14_n54 ; 
    wire[4:0] ILA___bv_5_15_n52 ; 
    wire[4:0] ILA___bv_5_16_n50 ; 
    wire[4:0] ILA___bv_5_17_n48 ; 
    wire[4:0] ILA___bv_5_18_n46 ; 
    wire[4:0] ILA___bv_5_19_n44 ; 
    wire[4:0] ILA___bv_5_1_n17 ; 
    wire[4:0] ILA___bv_5_20_n42 ; 
    wire[4:0] ILA___bv_5_21_n40 ; 
    wire[4:0] ILA___bv_5_22_n38 ; 
    wire[4:0] ILA___bv_5_23_n36 ; 
    wire[4:0] ILA___bv_5_24_n34 ; 
    wire[4:0] ILA___bv_5_25_n32 ; 
    wire[4:0] ILA___bv_5_26_n30 ; 
    wire[4:0] ILA___bv_5_27_n28 ; 
    wire[4:0] ILA___bv_5_28_n26 ; 
    wire[4:0] ILA___bv_5_29_n24 ; 
    wire[4:0] ILA___bv_5_2_n78 ; 
    wire[4:0] ILA___bv_5_30_n22 ; 
    wire[4:0] ILA___bv_5_31_n20 ; 
    wire[4:0] ILA___bv_5_3_n76 ; 
    wire[4:0] ILA___bv_5_4_n74 ; 
    wire[4:0] ILA___bv_5_5_n72 ; 
    wire[4:0] ILA___bv_5_6_n70 ; 
    wire[4:0] ILA___bv_5_7_n68 ; 
    wire[4:0] ILA___bv_5_8_n66 ; 
    wire[4:0] ILA___bv_5_9_n64 ; 
    wire[6:0] ILA___bv_7_0_n8 ; 
    wire[6:0] ILA___bv_7_51_n1 ; 
    wire ILA___clk ; 
    wire[31:0] ILA___inst ; 
    wire[31:0] ILA___load_addr_randinit ; 
    wire[31:0] ILA___load_data_randinit ; 
    wire ILA___load_en_randinit ; 
    wire[2:0] ILA___load_size_randinit ; 
    wire[6:0] ILA___n0 ; 
    wire ILA___n10 ; 
    wire[31:0] ILA___n100 ; 
    wire[31:0] ILA___n101 ; 
    wire[31:0] ILA___n102 ; 
    wire[31:0] ILA___n103 ; 
    wire[31:0] ILA___n104 ; 
    wire[31:0] ILA___n105 ; 
    wire[31:0] ILA___n106 ; 
    wire[31:0] ILA___n107 ; 
    wire[31:0] ILA___n108 ; 
    wire[31:0] ILA___n109 ; 
    wire[31:0] ILA___n110 ; 
    wire[31:0] ILA___n111 ; 
    wire[4:0] ILA___n112 ; 
    wire ILA___n113 ; 
    wire ILA___n114 ; 
    wire ILA___n115 ; 
    wire ILA___n116 ; 
    wire ILA___n117 ; 
    wire ILA___n118 ; 
    wire ILA___n119 ; 
    wire ILA___n120 ; 
    wire ILA___n121 ; 
    wire ILA___n122 ; 
    wire ILA___n123 ; 
    wire ILA___n124 ; 
    wire ILA___n125 ; 
    wire ILA___n126 ; 
    wire ILA___n127 ; 
    wire ILA___n128 ; 
    wire ILA___n129 ; 
    wire[31:0] ILA___n13 ; 
    wire ILA___n130 ; 
    wire ILA___n131 ; 
    wire ILA___n132 ; 
    wire ILA___n133 ; 
    wire ILA___n134 ; 
    wire ILA___n135 ; 
    wire ILA___n136 ; 
    wire ILA___n137 ; 
    wire ILA___n138 ; 
    wire ILA___n139 ; 
    wire ILA___n140 ; 
    wire ILA___n141 ; 
    wire ILA___n142 ; 
    wire ILA___n143 ; 
    wire[31:0] ILA___n144 ; 
    wire[31:0] ILA___n145 ; 
    wire[31:0] ILA___n146 ; 
    wire[31:0] ILA___n147 ; 
    wire[31:0] ILA___n148 ; 
    wire[31:0] ILA___n149 ; 
    wire[31:0] ILA___n150 ; 
    wire[31:0] ILA___n151 ; 
    wire[31:0] ILA___n152 ; 
    wire[31:0] ILA___n153 ; 
    wire[31:0] ILA___n154 ; 
    wire[31:0] ILA___n155 ; 
    wire[31:0] ILA___n156 ; 
    wire[31:0] ILA___n157 ; 
    wire[31:0] ILA___n158 ; 
    wire[31:0] ILA___n159 ; 
    wire[4:0] ILA___n16 ; 
    wire[31:0] ILA___n160 ; 
    wire[31:0] ILA___n161 ; 
    wire[31:0] ILA___n162 ; 
    wire[31:0] ILA___n163 ; 
    wire[31:0] ILA___n164 ; 
    wire[31:0] ILA___n165 ; 
    wire[31:0] ILA___n166 ; 
    wire[31:0] ILA___n167 ; 
    wire[31:0] ILA___n168 ; 
    wire[31:0] ILA___n169 ; 
    wire[31:0] ILA___n170 ; 
    wire[31:0] ILA___n171 ; 
    wire[31:0] ILA___n172 ; 
    wire[31:0] ILA___n173 ; 
    wire[31:0] ILA___n174 ; 
    wire[31:0] ILA___n175 ; 
    wire[31:0] ILA___n176 ; 
    wire ILA___n177 ; 
    wire[31:0] ILA___n178 ; 
    wire ILA___n179 ; 
    wire ILA___n18 ; 
    wire[31:0] ILA___n180 ; 
    wire ILA___n181 ; 
    wire[31:0] ILA___n182 ; 
    wire ILA___n183 ; 
    wire[31:0] ILA___n184 ; 
    wire ILA___n185 ; 
    wire[31:0] ILA___n186 ; 
    wire ILA___n187 ; 
    wire[31:0] ILA___n188 ; 
    wire ILA___n189 ; 
    wire[4:0] ILA___n19 ; 
    wire[31:0] ILA___n190 ; 
    wire ILA___n191 ; 
    wire[31:0] ILA___n192 ; 
    wire ILA___n193 ; 
    wire[31:0] ILA___n194 ; 
    wire ILA___n195 ; 
    wire[31:0] ILA___n196 ; 
    wire ILA___n197 ; 
    wire[31:0] ILA___n198 ; 
    wire ILA___n199 ; 
    wire ILA___n2 ; 
    wire[31:0] ILA___n200 ; 
    wire ILA___n201 ; 
    wire[31:0] ILA___n202 ; 
    wire ILA___n203 ; 
    wire[31:0] ILA___n204 ; 
    wire ILA___n205 ; 
    wire[31:0] ILA___n206 ; 
    wire ILA___n207 ; 
    wire[31:0] ILA___n208 ; 
    wire ILA___n209 ; 
    wire ILA___n21 ; 
    wire[31:0] ILA___n210 ; 
    wire ILA___n211 ; 
    wire[31:0] ILA___n212 ; 
    wire ILA___n213 ; 
    wire[31:0] ILA___n214 ; 
    wire ILA___n215 ; 
    wire[31:0] ILA___n216 ; 
    wire ILA___n217 ; 
    wire[31:0] ILA___n218 ; 
    wire ILA___n219 ; 
    wire[31:0] ILA___n220 ; 
    wire ILA___n221 ; 
    wire[31:0] ILA___n222 ; 
    wire ILA___n223 ; 
    wire[31:0] ILA___n224 ; 
    wire ILA___n225 ; 
    wire[31:0] ILA___n226 ; 
    wire ILA___n227 ; 
    wire[31:0] ILA___n228 ; 
    wire ILA___n229 ; 
    wire ILA___n23 ; 
    wire[31:0] ILA___n230 ; 
    wire ILA___n231 ; 
    wire[31:0] ILA___n232 ; 
    wire ILA___n233 ; 
    wire[31:0] ILA___n234 ; 
    wire ILA___n235 ; 
    wire[31:0] ILA___n236 ; 
    wire ILA___n25 ; 
    wire ILA___n27 ; 
    wire ILA___n29 ; 
    wire[2:0] ILA___n3 ; 
    wire ILA___n31 ; 
    wire ILA___n33 ; 
    wire ILA___n35 ; 
    wire ILA___n37 ; 
    wire ILA___n39 ; 
    wire ILA___n41 ; 
    wire ILA___n43 ; 
    wire ILA___n45 ; 
    wire ILA___n47 ; 
    wire ILA___n49 ; 
    wire ILA___n5 ; 
    wire ILA___n51 ; 
    wire ILA___n53 ; 
    wire ILA___n55 ; 
    wire ILA___n57 ; 
    wire ILA___n59 ; 
    wire ILA___n6 ; 
    wire ILA___n61 ; 
    wire ILA___n63 ; 
    wire ILA___n65 ; 
    wire ILA___n67 ; 
    wire ILA___n69 ; 
    wire[6:0] ILA___n7 ; 
    wire ILA___n71 ; 
    wire ILA___n73 ; 
    wire ILA___n75 ; 
    wire ILA___n77 ; 
    wire ILA___n79 ; 
    wire ILA___n80 ; 
    wire[31:0] ILA___n81 ; 
    wire[31:0] ILA___n82 ; 
    wire[31:0] ILA___n83 ; 
    wire[31:0] ILA___n84 ; 
    wire[31:0] ILA___n85 ; 
    wire[31:0] ILA___n86 ; 
    wire[31:0] ILA___n87 ; 
    wire[31:0] ILA___n88 ; 
    wire[31:0] ILA___n89 ; 
    wire ILA___n9 ; 
    wire[31:0] ILA___n90 ; 
    wire[31:0] ILA___n91 ; 
    wire[31:0] ILA___n92 ; 
    wire[31:0] ILA___n93 ; 
    wire[31:0] ILA___n94 ; 
    wire[31:0] ILA___n95 ; 
    wire[31:0] ILA___n96 ; 
    wire[31:0] ILA___n97 ; 
    wire[31:0] ILA___n98 ; 
    wire[31:0] ILA___n99 ; 
    wire[31:0] ILA___pc_randinit ; 
    wire ILA___rst ; 
    wire[31:0] ILA___store_addr_randinit ; 
    wire[31:0] ILA___store_data_randinit ; 
    wire ILA___store_en_randinit ; 
    wire[2:0] ILA___store_size_randinit ; 
    wire[31:0] ILA___x0_randinit ; 
    wire[31:0] ILA___x10_randinit ; 
    wire[31:0] ILA___x11_randinit ; 
    wire[31:0] ILA___x12_randinit ; 
    wire[31:0] ILA___x13_randinit ; 
    wire[31:0] ILA___x14_randinit ; 
    wire[31:0] ILA___x15_randinit ; 
    wire[31:0] ILA___x16_randinit ; 
    wire[31:0] ILA___x17_randinit ; 
    wire[31:0] ILA___x18_randinit ; 
    wire[31:0] ILA___x19_randinit ; 
    wire[31:0] ILA___x1_randinit ; 
    wire[31:0] ILA___x20_randinit ; 
    wire[31:0] ILA___x21_randinit ; 
    wire[31:0] ILA___x22_randinit ; 
    wire[31:0] ILA___x23_randinit ; 
    wire[31:0] ILA___x24_randinit ; 
    wire[31:0] ILA___x25_randinit ; 
    wire[31:0] ILA___x26_randinit ; 
    wire[31:0] ILA___x27_randinit ; 
    wire[31:0] ILA___x28_randinit ; 
    wire[31:0] ILA___x29_randinit ; 
    wire[31:0] ILA___x2_randinit ; 
    wire[31:0] ILA___x30_randinit ; 
    wire[31:0] ILA___x31_randinit ; 
    wire[31:0] ILA___x3_randinit ; 
    wire[31:0] ILA___x4_randinit ; 
    wire[31:0] ILA___x5_randinit ; 
    wire[31:0] ILA___x6_randinit ; 
    wire[31:0] ILA___x7_randinit ; 
    wire[31:0] ILA___x8_randinit ; 
    wire[31:0] ILA___x9_randinit ; 
  assign  ILA_____ILA_riscv_valid__ =1'b1; 
  assign  ILA___n0 = ILA___inst [6:0]; 
  assign  ILA___bv_7_51_n1 =7'h33; 
  assign  ILA___n2 =( ILA___n0 )==( ILA___bv_7_51_n1 ); 
  assign  ILA___n3 = ILA___inst [14:12]; 
  assign  ILA___bv_3_0_n4 =3'h0; 
  assign  ILA___n5 =( ILA___n3 )==( ILA___bv_3_0_n4 ); 
  assign  ILA___n6 =( ILA___n2 )&( ILA___n5 ); 
  assign  ILA___n7 = ILA___inst [31:25]; 
  assign  ILA___bv_7_0_n8 =7'h0; 
  assign  ILA___n9 =( ILA___n7 )==( ILA___bv_7_0_n8 ); 
  assign  ILA___n10 =( ILA___n6 )&( ILA___n9 ); 
  assign  ILA_____ILA_riscv_decode_of_ADD__ = ILA___n10 ; 
  assign  ILA___bv_32_4_n12 =32'h4; 
  assign  ILA___n13 =( ILA___pc )+( ILA___bv_32_4_n12 ); 
  assign  ILA___bv_1_0_n14 =1'h0; 
  assign  ILA___bv_32_0_n15 =32'h0; 
  assign  ILA___n16 = ILA___inst [11:7]; 
  assign  ILA___bv_5_1_n17 =5'h1; 
  assign  ILA___n18 =( ILA___n16 )==( ILA___bv_5_1_n17 ); 
  assign  ILA___n19 = ILA___inst [19:15]; 
  assign  ILA___bv_5_31_n20 =5'h1f; 
  assign  ILA___n21 =( ILA___n19 )==( ILA___bv_5_31_n20 ); 
  assign  ILA___bv_5_30_n22 =5'h1e; 
  assign  ILA___n23 =( ILA___n19 )==( ILA___bv_5_30_n22 ); 
  assign  ILA___bv_5_29_n24 =5'h1d; 
  assign  ILA___n25 =( ILA___n19 )==( ILA___bv_5_29_n24 ); 
  assign  ILA___bv_5_28_n26 =5'h1c; 
  assign  ILA___n27 =( ILA___n19 )==( ILA___bv_5_28_n26 ); 
  assign  ILA___bv_5_27_n28 =5'h1b; 
  assign  ILA___n29 =( ILA___n19 )==( ILA___bv_5_27_n28 ); 
  assign  ILA___bv_5_26_n30 =5'h1a; 
  assign  ILA___n31 =( ILA___n19 )==( ILA___bv_5_26_n30 ); 
  assign  ILA___bv_5_25_n32 =5'h19; 
  assign  ILA___n33 =( ILA___n19 )==( ILA___bv_5_25_n32 ); 
  assign  ILA___bv_5_24_n34 =5'h18; 
  assign  ILA___n35 =( ILA___n19 )==( ILA___bv_5_24_n34 ); 
  assign  ILA___bv_5_23_n36 =5'h17; 
  assign  ILA___n37 =( ILA___n19 )==( ILA___bv_5_23_n36 ); 
  assign  ILA___bv_5_22_n38 =5'h16; 
  assign  ILA___n39 =( ILA___n19 )==( ILA___bv_5_22_n38 ); 
  assign  ILA___bv_5_21_n40 =5'h15; 
  assign  ILA___n41 =( ILA___n19 )==( ILA___bv_5_21_n40 ); 
  assign  ILA___bv_5_20_n42 =5'h14; 
  assign  ILA___n43 =( ILA___n19 )==( ILA___bv_5_20_n42 ); 
  assign  ILA___bv_5_19_n44 =5'h13; 
  assign  ILA___n45 =( ILA___n19 )==( ILA___bv_5_19_n44 ); 
  assign  ILA___bv_5_18_n46 =5'h12; 
  assign  ILA___n47 =( ILA___n19 )==( ILA___bv_5_18_n46 ); 
  assign  ILA___bv_5_17_n48 =5'h11; 
  assign  ILA___n49 =( ILA___n19 )==( ILA___bv_5_17_n48 ); 
  assign  ILA___bv_5_16_n50 =5'h10; 
  assign  ILA___n51 =( ILA___n19 )==( ILA___bv_5_16_n50 ); 
  assign  ILA___bv_5_15_n52 =5'hf; 
  assign  ILA___n53 =( ILA___n19 )==( ILA___bv_5_15_n52 ); 
  assign  ILA___bv_5_14_n54 =5'he; 
  assign  ILA___n55 =( ILA___n19 )==( ILA___bv_5_14_n54 ); 
  assign  ILA___bv_5_13_n56 =5'hd; 
  assign  ILA___n57 =( ILA___n19 )==( ILA___bv_5_13_n56 ); 
  assign  ILA___bv_5_12_n58 =5'hc; 
  assign  ILA___n59 =( ILA___n19 )==( ILA___bv_5_12_n58 ); 
  assign  ILA___bv_5_11_n60 =5'hb; 
  assign  ILA___n61 =( ILA___n19 )==( ILA___bv_5_11_n60 ); 
  assign  ILA___bv_5_10_n62 =5'ha; 
  assign  ILA___n63 =( ILA___n19 )==( ILA___bv_5_10_n62 ); 
  assign  ILA___bv_5_9_n64 =5'h9; 
  assign  ILA___n65 =( ILA___n19 )==( ILA___bv_5_9_n64 ); 
  assign  ILA___bv_5_8_n66 =5'h8; 
  assign  ILA___n67 =( ILA___n19 )==( ILA___bv_5_8_n66 ); 
  assign  ILA___bv_5_7_n68 =5'h7; 
  assign  ILA___n69 =( ILA___n19 )==( ILA___bv_5_7_n68 ); 
  assign  ILA___bv_5_6_n70 =5'h6; 
  assign  ILA___n71 =( ILA___n19 )==( ILA___bv_5_6_n70 ); 
  assign  ILA___bv_5_5_n72 =5'h5; 
  assign  ILA___n73 =( ILA___n19 )==( ILA___bv_5_5_n72 ); 
  assign  ILA___bv_5_4_n74 =5'h4; 
  assign  ILA___n75 =( ILA___n19 )==( ILA___bv_5_4_n74 ); 
  assign  ILA___bv_5_3_n76 =5'h3; 
  assign  ILA___n77 =( ILA___n19 )==( ILA___bv_5_3_n76 ); 
  assign  ILA___bv_5_2_n78 =5'h2; 
  assign  ILA___n79 =( ILA___n19 )==( ILA___bv_5_2_n78 ); 
  assign  ILA___n80 =( ILA___n19 )==( ILA___bv_5_1_n17 ); 
  assign  ILA___n81 =( ILA___n80 ) ? ( ILA___x1 ):( ILA___bv_32_0_n15 ); 
  assign  ILA___n82 =( ILA___n79 ) ? ( ILA___x2 ):( ILA___n81 ); 
  assign  ILA___n83 =( ILA___n77 ) ? ( ILA___x3 ):( ILA___n82 ); 
  assign  ILA___n84 =( ILA___n75 ) ? ( ILA___x4 ):( ILA___n83 ); 
  assign  ILA___n85 =( ILA___n73 ) ? ( ILA___x5 ):( ILA___n84 ); 
  assign  ILA___n86 =( ILA___n71 ) ? ( ILA___x6 ):( ILA___n85 ); 
  assign  ILA___n87 =( ILA___n69 ) ? ( ILA___x7 ):( ILA___n86 ); 
  assign  ILA___n88 =( ILA___n67 ) ? ( ILA___x8 ):( ILA___n87 ); 
  assign  ILA___n89 =( ILA___n65 ) ? ( ILA___x9 ):( ILA___n88 ); 
  assign  ILA___n90 =( ILA___n63 ) ? ( ILA___x10 ):( ILA___n89 ); 
  assign  ILA___n91 =( ILA___n61 ) ? ( ILA___x11 ):( ILA___n90 ); 
  assign  ILA___n92 =( ILA___n59 ) ? ( ILA___x12 ):( ILA___n91 ); 
  assign  ILA___n93 =( ILA___n57 ) ? ( ILA___x13 ):( ILA___n92 ); 
  assign  ILA___n94 =( ILA___n55 ) ? ( ILA___x14 ):( ILA___n93 ); 
  assign  ILA___n95 =( ILA___n53 ) ? ( ILA___x15 ):( ILA___n94 ); 
  assign  ILA___n96 =( ILA___n51 ) ? ( ILA___x16 ):( ILA___n95 ); 
  assign  ILA___n97 =( ILA___n49 ) ? ( ILA___x17 ):( ILA___n96 ); 
  assign  ILA___n98 =( ILA___n47 ) ? ( ILA___x18 ):( ILA___n97 ); 
  assign  ILA___n99 =( ILA___n45 ) ? ( ILA___x19 ):( ILA___n98 ); 
  assign  ILA___n100 =( ILA___n43 ) ? ( ILA___x20 ):( ILA___n99 ); 
  assign  ILA___n101 =( ILA___n41 ) ? ( ILA___x21 ):( ILA___n100 ); 
  assign  ILA___n102 =( ILA___n39 ) ? ( ILA___x22 ):( ILA___n101 ); 
  assign  ILA___n103 =( ILA___n37 ) ? ( ILA___x23 ):( ILA___n102 ); 
  assign  ILA___n104 =( ILA___n35 ) ? ( ILA___x24 ):( ILA___n103 ); 
  assign  ILA___n105 =( ILA___n33 ) ? ( ILA___x25 ):( ILA___n104 ); 
  assign  ILA___n106 =( ILA___n31 ) ? ( ILA___x26 ):( ILA___n105 ); 
  assign  ILA___n107 =( ILA___n29 ) ? ( ILA___x27 ):( ILA___n106 ); 
  assign  ILA___n108 =( ILA___n27 ) ? ( ILA___x28 ):( ILA___n107 ); 
  assign  ILA___n109 =( ILA___n25 ) ? ( ILA___x29 ):( ILA___n108 ); 
  assign  ILA___n110 =( ILA___n23 ) ? ( ILA___x30 ):( ILA___n109 ); 
  assign  ILA___n111 =( ILA___n21 ) ? ( ILA___x31 ):( ILA___n110 ); 
  assign  ILA___n112 = ILA___inst [24:20]; 
  assign  ILA___n113 =( ILA___n112 )==( ILA___bv_5_31_n20 ); 
  assign  ILA___n114 =( ILA___n112 )==( ILA___bv_5_30_n22 ); 
  assign  ILA___n115 =( ILA___n112 )==( ILA___bv_5_29_n24 ); 
  assign  ILA___n116 =( ILA___n112 )==( ILA___bv_5_28_n26 ); 
  assign  ILA___n117 =( ILA___n112 )==( ILA___bv_5_27_n28 ); 
  assign  ILA___n118 =( ILA___n112 )==( ILA___bv_5_26_n30 ); 
  assign  ILA___n119 =( ILA___n112 )==( ILA___bv_5_25_n32 ); 
  assign  ILA___n120 =( ILA___n112 )==( ILA___bv_5_24_n34 ); 
  assign  ILA___n121 =( ILA___n112 )==( ILA___bv_5_23_n36 ); 
  assign  ILA___n122 =( ILA___n112 )==( ILA___bv_5_22_n38 ); 
  assign  ILA___n123 =( ILA___n112 )==( ILA___bv_5_21_n40 ); 
  assign  ILA___n124 =( ILA___n112 )==( ILA___bv_5_20_n42 ); 
  assign  ILA___n125 =( ILA___n112 )==( ILA___bv_5_19_n44 ); 
  assign  ILA___n126 =( ILA___n112 )==( ILA___bv_5_18_n46 ); 
  assign  ILA___n127 =( ILA___n112 )==( ILA___bv_5_17_n48 ); 
  assign  ILA___n128 =( ILA___n112 )==( ILA___bv_5_16_n50 ); 
  assign  ILA___n129 =( ILA___n112 )==( ILA___bv_5_15_n52 ); 
  assign  ILA___n130 =( ILA___n112 )==( ILA___bv_5_14_n54 ); 
  assign  ILA___n131 =( ILA___n112 )==( ILA___bv_5_13_n56 ); 
  assign  ILA___n132 =( ILA___n112 )==( ILA___bv_5_12_n58 ); 
  assign  ILA___n133 =( ILA___n112 )==( ILA___bv_5_11_n60 ); 
  assign  ILA___n134 =( ILA___n112 )==( ILA___bv_5_10_n62 ); 
  assign  ILA___n135 =( ILA___n112 )==( ILA___bv_5_9_n64 ); 
  assign  ILA___n136 =( ILA___n112 )==( ILA___bv_5_8_n66 ); 
  assign  ILA___n137 =( ILA___n112 )==( ILA___bv_5_7_n68 ); 
  assign  ILA___n138 =( ILA___n112 )==( ILA___bv_5_6_n70 ); 
  assign  ILA___n139 =( ILA___n112 )==( ILA___bv_5_5_n72 ); 
  assign  ILA___n140 =( ILA___n112 )==( ILA___bv_5_4_n74 ); 
  assign  ILA___n141 =( ILA___n112 )==( ILA___bv_5_3_n76 ); 
  assign  ILA___n142 =( ILA___n112 )==( ILA___bv_5_2_n78 ); 
  assign  ILA___n143 =( ILA___n112 )==( ILA___bv_5_1_n17 ); 
  assign  ILA___n144 =( ILA___n143 ) ? ( ILA___x1 ):( ILA___bv_32_0_n15 ); 
  assign  ILA___n145 =( ILA___n142 ) ? ( ILA___x2 ):( ILA___n144 ); 
  assign  ILA___n146 =( ILA___n141 ) ? ( ILA___x3 ):( ILA___n145 ); 
  assign  ILA___n147 =( ILA___n140 ) ? ( ILA___x4 ):( ILA___n146 ); 
  assign  ILA___n148 =( ILA___n139 ) ? ( ILA___x5 ):( ILA___n147 ); 
  assign  ILA___n149 =( ILA___n138 ) ? ( ILA___x6 ):( ILA___n148 ); 
  assign  ILA___n150 =( ILA___n137 ) ? ( ILA___x7 ):( ILA___n149 ); 
  assign  ILA___n151 =( ILA___n136 ) ? ( ILA___x8 ):( ILA___n150 ); 
  assign  ILA___n152 =( ILA___n135 ) ? ( ILA___x9 ):( ILA___n151 ); 
  assign  ILA___n153 =( ILA___n134 ) ? ( ILA___x10 ):( ILA___n152 ); 
  assign  ILA___n154 =( ILA___n133 ) ? ( ILA___x11 ):( ILA___n153 ); 
  assign  ILA___n155 =( ILA___n132 ) ? ( ILA___x12 ):( ILA___n154 ); 
  assign  ILA___n156 =( ILA___n131 ) ? ( ILA___x13 ):( ILA___n155 ); 
  assign  ILA___n157 =( ILA___n130 ) ? ( ILA___x14 ):( ILA___n156 ); 
  assign  ILA___n158 =( ILA___n129 ) ? ( ILA___x15 ):( ILA___n157 ); 
  assign  ILA___n159 =( ILA___n128 ) ? ( ILA___x16 ):( ILA___n158 ); 
  assign  ILA___n160 =( ILA___n127 ) ? ( ILA___x17 ):( ILA___n159 ); 
  assign  ILA___n161 =( ILA___n126 ) ? ( ILA___x18 ):( ILA___n160 ); 
  assign  ILA___n162 =( ILA___n125 ) ? ( ILA___x19 ):( ILA___n161 ); 
  assign  ILA___n163 =( ILA___n124 ) ? ( ILA___x20 ):( ILA___n162 ); 
  assign  ILA___n164 =( ILA___n123 ) ? ( ILA___x21 ):( ILA___n163 ); 
  assign  ILA___n165 =( ILA___n122 ) ? ( ILA___x22 ):( ILA___n164 ); 
  assign  ILA___n166 =( ILA___n121 ) ? ( ILA___x23 ):( ILA___n165 ); 
  assign  ILA___n167 =( ILA___n120 ) ? ( ILA___x24 ):( ILA___n166 ); 
  assign  ILA___n168 =( ILA___n119 ) ? ( ILA___x25 ):( ILA___n167 ); 
  assign  ILA___n169 =( ILA___n118 ) ? ( ILA___x26 ):( ILA___n168 ); 
  assign  ILA___n170 =( ILA___n117 ) ? ( ILA___x27 ):( ILA___n169 ); 
  assign  ILA___n171 =( ILA___n116 ) ? ( ILA___x28 ):( ILA___n170 ); 
  assign  ILA___n172 =( ILA___n115 ) ? ( ILA___x29 ):( ILA___n171 ); 
  assign  ILA___n173 =( ILA___n114 ) ? ( ILA___x30 ):( ILA___n172 ); 
  assign  ILA___n174 =( ILA___n113 ) ? ( ILA___x31 ):( ILA___n173 ); 
  assign  ILA___n175 =( ILA___n111 )+( ILA___n174 ); 
  assign  ILA___n176 =( ILA___n18 ) ? ( ILA___n175 ):( ILA___x1 ); 
  assign  ILA___n177 =( ILA___n16 )==( ILA___bv_5_2_n78 ); 
  assign  ILA___n178 =( ILA___n177 ) ? ( ILA___n175 ):( ILA___x2 ); 
  assign  ILA___n179 =( ILA___n16 )==( ILA___bv_5_3_n76 ); 
  assign  ILA___n180 =( ILA___n179 ) ? ( ILA___n175 ):( ILA___x3 ); 
  assign  ILA___n181 =( ILA___n16 )==( ILA___bv_5_4_n74 ); 
  assign  ILA___n182 =( ILA___n181 ) ? ( ILA___n175 ):( ILA___x4 ); 
  assign  ILA___n183 =( ILA___n16 )==( ILA___bv_5_5_n72 ); 
  assign  ILA___n184 =( ILA___n183 ) ? ( ILA___n175 ):( ILA___x5 ); 
  assign  ILA___n185 =( ILA___n16 )==( ILA___bv_5_6_n70 ); 
  assign  ILA___n186 =( ILA___n185 ) ? ( ILA___n175 ):( ILA___x6 ); 
  assign  ILA___n187 =( ILA___n16 )==( ILA___bv_5_7_n68 ); 
  assign  ILA___n188 =( ILA___n187 ) ? ( ILA___n175 ):( ILA___x7 ); 
  assign  ILA___n189 =( ILA___n16 )==( ILA___bv_5_8_n66 ); 
  assign  ILA___n190 =( ILA___n189 ) ? ( ILA___n175 ):( ILA___x8 ); 
  assign  ILA___n191 =( ILA___n16 )==( ILA___bv_5_9_n64 ); 
  assign  ILA___n192 =( ILA___n191 ) ? ( ILA___n175 ):( ILA___x9 ); 
  assign  ILA___n193 =( ILA___n16 )==( ILA___bv_5_10_n62 ); 
  assign  ILA___n194 =( ILA___n193 ) ? ( ILA___n175 ):( ILA___x10 ); 
  assign  ILA___n195 =( ILA___n16 )==( ILA___bv_5_11_n60 ); 
  assign  ILA___n196 =( ILA___n195 ) ? ( ILA___n175 ):( ILA___x11 ); 
  assign  ILA___n197 =( ILA___n16 )==( ILA___bv_5_12_n58 ); 
  assign  ILA___n198 =( ILA___n197 ) ? ( ILA___n175 ):( ILA___x12 ); 
  assign  ILA___n199 =( ILA___n16 )==( ILA___bv_5_13_n56 ); 
  assign  ILA___n200 =( ILA___n199 ) ? ( ILA___n175 ):( ILA___x13 ); 
  assign  ILA___n201 =( ILA___n16 )==( ILA___bv_5_14_n54 ); 
  assign  ILA___n202 =( ILA___n201 ) ? ( ILA___n175 ):( ILA___x14 ); 
  assign  ILA___n203 =( ILA___n16 )==( ILA___bv_5_15_n52 ); 
  assign  ILA___n204 =( ILA___n203 ) ? ( ILA___n175 ):( ILA___x15 ); 
  assign  ILA___n205 =( ILA___n16 )==( ILA___bv_5_16_n50 ); 
  assign  ILA___n206 =( ILA___n205 ) ? ( ILA___n175 ):( ILA___x16 ); 
  assign  ILA___n207 =( ILA___n16 )==( ILA___bv_5_17_n48 ); 
  assign  ILA___n208 =( ILA___n207 ) ? ( ILA___n175 ):( ILA___x17 ); 
  assign  ILA___n209 =( ILA___n16 )==( ILA___bv_5_18_n46 ); 
  assign  ILA___n210 =( ILA___n209 ) ? ( ILA___n175 ):( ILA___x18 ); 
  assign  ILA___n211 =( ILA___n16 )==( ILA___bv_5_19_n44 ); 
  assign  ILA___n212 =( ILA___n211 ) ? ( ILA___n175 ):( ILA___x19 ); 
  assign  ILA___n213 =( ILA___n16 )==( ILA___bv_5_20_n42 ); 
  assign  ILA___n214 =( ILA___n213 ) ? ( ILA___n175 ):( ILA___x20 ); 
  assign  ILA___n215 =( ILA___n16 )==( ILA___bv_5_21_n40 ); 
  assign  ILA___n216 =( ILA___n215 ) ? ( ILA___n175 ):( ILA___x21 ); 
  assign  ILA___n217 =( ILA___n16 )==( ILA___bv_5_22_n38 ); 
  assign  ILA___n218 =( ILA___n217 ) ? ( ILA___n175 ):( ILA___x22 ); 
  assign  ILA___n219 =( ILA___n16 )==( ILA___bv_5_23_n36 ); 
  assign  ILA___n220 =( ILA___n219 ) ? ( ILA___n175 ):( ILA___x23 ); 
  assign  ILA___n221 =( ILA___n16 )==( ILA___bv_5_24_n34 ); 
  assign  ILA___n222 =( ILA___n221 ) ? ( ILA___n175 ):( ILA___x24 ); 
  assign  ILA___n223 =( ILA___n16 )==( ILA___bv_5_25_n32 ); 
  assign  ILA___n224 =( ILA___n223 ) ? ( ILA___n175 ):( ILA___x25 ); 
  assign  ILA___n225 =( ILA___n16 )==( ILA___bv_5_26_n30 ); 
  assign  ILA___n226 =( ILA___n225 ) ? ( ILA___n175 ):( ILA___x26 ); 
  assign  ILA___n227 =( ILA___n16 )==( ILA___bv_5_27_n28 ); 
  assign  ILA___n228 =( ILA___n227 ) ? ( ILA___n175 ):( ILA___x27 ); 
  assign  ILA___n229 =( ILA___n16 )==( ILA___bv_5_28_n26 ); 
  assign  ILA___n230 =( ILA___n229 ) ? ( ILA___n175 ):( ILA___x28 ); 
  assign  ILA___n231 =( ILA___n16 )==( ILA___bv_5_29_n24 ); 
  assign  ILA___n232 =( ILA___n231 ) ? ( ILA___n175 ):( ILA___x29 ); 
  assign  ILA___n233 =( ILA___n16 )==( ILA___bv_5_30_n22 ); 
  assign  ILA___n234 =( ILA___n233 ) ? ( ILA___n175 ):( ILA___x30 ); 
  assign  ILA___n235 =( ILA___n16 )==( ILA___bv_5_31_n20 ); 
  assign  ILA___n236 =( ILA___n235 ) ? ( ILA___n175 ):( ILA___x31 ); 
  always @( posedge  ILA___clk )
         begin 
             if ( ILA___rst )
                 begin  
                     ILA___pc  <= ILA___pc_randinit ; 
                     ILA___load_en  <= ILA___load_en_randinit ; 
                     ILA___load_addr  <= ILA___load_addr_randinit ; 
                     ILA___load_size  <= ILA___load_size_randinit ; 
                     ILA___load_data  <= ILA___load_data_randinit ; 
                     ILA___store_en  <= ILA___store_en_randinit ; 
                     ILA___store_addr  <= ILA___store_addr_randinit ; 
                     ILA___store_size  <= ILA___store_size_randinit ; 
                     ILA___store_data  <= ILA___store_data_randinit ; 
                     ILA___x0  <= ILA___x0_randinit ; 
                     ILA___x1  <= ILA___x1_randinit ; 
                     ILA___x2  <= ILA___x2_randinit ; 
                     ILA___x3  <= ILA___x3_randinit ; 
                     ILA___x4  <= ILA___x4_randinit ; 
                     ILA___x5  <= ILA___x5_randinit ; 
                     ILA___x6  <= ILA___x6_randinit ; 
                     ILA___x7  <= ILA___x7_randinit ; 
                     ILA___x8  <= ILA___x8_randinit ; 
                     ILA___x9  <= ILA___x9_randinit ; 
                     ILA___x10  <= ILA___x10_randinit ; 
                     ILA___x11  <= ILA___x11_randinit ; 
                     ILA___x12  <= ILA___x12_randinit ; 
                     ILA___x13  <= ILA___x13_randinit ; 
                     ILA___x14  <= ILA___x14_randinit ; 
                     ILA___x15  <= ILA___x15_randinit ; 
                     ILA___x16  <= ILA___x16_randinit ; 
                     ILA___x17  <= ILA___x17_randinit ; 
                     ILA___x18  <= ILA___x18_randinit ; 
                     ILA___x19  <= ILA___x19_randinit ; 
                     ILA___x20  <= ILA___x20_randinit ; 
                     ILA___x21  <= ILA___x21_randinit ; 
                     ILA___x22  <= ILA___x22_randinit ; 
                     ILA___x23  <= ILA___x23_randinit ; 
                     ILA___x24  <= ILA___x24_randinit ; 
                     ILA___x25  <= ILA___x25_randinit ; 
                     ILA___x26  <= ILA___x26_randinit ; 
                     ILA___x27  <= ILA___x27_randinit ; 
                     ILA___x28  <= ILA___x28_randinit ; 
                     ILA___x29  <= ILA___x29_randinit ; 
                     ILA___x30  <= ILA___x30_randinit ; 
                     ILA___x31  <= ILA___x31_randinit ; 
                     ILA_____COUNTER_start__n11  <=0;
                 end 
              else 
                 if ( ILA_____START__ && ILA_____ILA_riscv_valid__ )
                     begin 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA_____COUNTER_start__n11  <=1;
                             end 
                          else 
                             if (( ILA_____COUNTER_start__n11 >=1)&&( ILA_____COUNTER_start__n11 <255))
                                 begin  
                                     ILA_____COUNTER_start__n11  <= ILA_____COUNTER_start__n11 +1;
                                 end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___pc  <= ILA___n13 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___load_en  <= ILA___bv_1_0_n14 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___load_addr  <= ILA___load_addr ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___load_size  <= ILA___load_size ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___load_data  <= ILA___load_data ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___store_en  <= ILA___bv_1_0_n14 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___store_addr  <= ILA___store_addr ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___store_size  <= ILA___store_size ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___store_data  <= ILA___store_data ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x0  <= ILA___bv_32_0_n15 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x1  <= ILA___n176 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x2  <= ILA___n178 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x3  <= ILA___n180 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x4  <= ILA___n182 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x5  <= ILA___n184 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x6  <= ILA___n186 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x7  <= ILA___n188 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x8  <= ILA___n190 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x9  <= ILA___n192 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x10  <= ILA___n194 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x11  <= ILA___n196 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x12  <= ILA___n198 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x13  <= ILA___n200 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x14  <= ILA___n202 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x15  <= ILA___n204 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x16  <= ILA___n206 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x17  <= ILA___n208 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x18  <= ILA___n210 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x19  <= ILA___n212 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x20  <= ILA___n214 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x21  <= ILA___n216 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x22  <= ILA___n218 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x23  <= ILA___n220 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x24  <= ILA___n222 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x25  <= ILA___n224 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x26  <= ILA___n226 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x27  <= ILA___n228 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x28  <= ILA___n230 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x29  <= ILA___n232 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x30  <= ILA___n234 ;
                             end 
                         if ( ILA_____ILA_riscv_decode_of_ADD__ )
                             begin  
                                 ILA___x31  <= ILA___n236 ;
                             end 
                     end 
         end
 
    assign ILA_____START__ = __START__;
    assign ILA___clk = clk;
    assign ILA___inst = __ILA_I_inst;
    assign ILA___rst = rst;
    assign __ILA_riscv_decode_of_ADD__ = ILA_____ILA_riscv_decode_of_ADD__;
    assign __ILA_riscv_valid__ = ILA_____ILA_riscv_valid__;
    assign __ILA_SO_pc = ILA___pc;
    assign __ILA_SO_load_en = ILA___load_en;
    assign __ILA_SO_load_addr = ILA___load_addr;
    assign __ILA_SO_load_size = ILA___load_size;
    assign __ILA_SO_load_data = ILA___load_data;
    assign __ILA_SO_store_en = ILA___store_en;
    assign __ILA_SO_store_addr = ILA___store_addr;
    assign __ILA_SO_store_size = ILA___store_size;
    assign __ILA_SO_store_data = ILA___store_data;
    assign __ILA_SO_x0 = ILA___x0;
    assign __ILA_SO_x1 = ILA___x1;
    assign __ILA_SO_x2 = ILA___x2;
    assign __ILA_SO_x3 = ILA___x3;
    assign __ILA_SO_x4 = ILA___x4;
    assign __ILA_SO_x5 = ILA___x5;
    assign __ILA_SO_x6 = ILA___x6;
    assign __ILA_SO_x7 = ILA___x7;
    assign __ILA_SO_x8 = ILA___x8;
    assign __ILA_SO_x9 = ILA___x9;
    assign __ILA_SO_x10 = ILA___x10;
    assign __ILA_SO_x11 = ILA___x11;
    assign __ILA_SO_x12 = ILA___x12;
    assign __ILA_SO_x13 = ILA___x13;
    assign __ILA_SO_x14 = ILA___x14;
    assign __ILA_SO_x15 = ILA___x15;
    assign __ILA_SO_x16 = ILA___x16;
    assign __ILA_SO_x17 = ILA___x17;
    assign __ILA_SO_x18 = ILA___x18;
    assign __ILA_SO_x19 = ILA___x19;
    assign __ILA_SO_x20 = ILA___x20;
    assign __ILA_SO_x21 = ILA___x21;
    assign __ILA_SO_x22 = ILA___x22;
    assign __ILA_SO_x23 = ILA___x23;
    assign __ILA_SO_x24 = ILA___x24;
    assign __ILA_SO_x25 = ILA___x25;
    assign __ILA_SO_x26 = ILA___x26;
    assign __ILA_SO_x27 = ILA___x27;
    assign __ILA_SO_x28 = ILA___x28;
    assign __ILA_SO_x29 = ILA___x29;
    assign __ILA_SO_x30 = ILA___x30;
    assign __ILA_SO_x31 = ILA___x31;
    
assign __EDCOND__ = (end_of_pipeline)&&(__STARTED__) ;
assign __IEND__ = ((((end_of_pipeline)&&(__STARTED__))&&(__RESETED__))&&(!(__ENDED__)))&&(1'b1) ;
assign __VLG_II_m_external_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_nmi_req_set_not_clear = 1'b0 ;
assign __VLG_II_s_external_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_software_interrupt_req_set_not_clear = 1'b0 ;
assign __VLG_II_timer_interrupt_req_set_not_clear = 1'b0 ;
assign __auxvar10__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar10__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ ;
assign __auxvar11__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar11__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ ;
assign __auxvar12__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar12__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ ;
assign __auxvar13__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar13__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ ;
assign __auxvar14__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar14__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ ;
assign __auxvar15__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar15__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ ;
assign __auxvar16__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar16__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ ;
assign __auxvar17__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar17__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ ;
assign __auxvar18__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar18__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ ;
assign __auxvar19__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar19__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ ;
assign __auxvar1__recorder_sn_cond = ((monitor_s2)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar1__recorder_sn_value = RTL__DOT__near_mem$imem_pc ;
assign __auxvar20__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar20__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ ;
assign __auxvar21__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar21__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ ;
assign __auxvar22__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar22__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ ;
assign __auxvar23__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar23__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ ;
assign __auxvar24__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar24__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ ;
assign __auxvar25__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar25__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ ;
assign __auxvar26__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar26__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ ;
assign __auxvar27__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar27__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ ;
assign __auxvar28__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar28__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ ;
assign __auxvar29__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar29__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ ;
assign __auxvar2__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar2__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ ;
assign __auxvar30__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar30__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ ;
assign __auxvar31__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar31__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ ;
assign __auxvar32__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar32__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ ;
assign __auxvar33__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar33__recorder_sn_value = RTL__DOT__near_mem$dmem_req_addr ;
assign __auxvar34__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar34__recorder_sn_value = RTL__DOT__near_mem$EN_dmem_req ;
assign __auxvar35__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar35__recorder_sn_value = RTL__DOT__near_mem$dmem_req_f3 ;
assign __auxvar36__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar36__recorder_sn_value = RTL__DOT__near_mem$dmem_req_op ;
assign __auxvar37__recorder_sn_cond = ((monitor_s2)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar37__recorder_sn_value = RTL__DOT__near_mem$dmem_word64[31:0] ;
assign __auxvar38__recorder_sn_cond = ((monitor_s1)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar38__recorder_sn_value = RTL__DOT__near_mem$dmem_req_store_value[31:0] ;
assign __auxvar3__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar3__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ ;
assign __auxvar4__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar4__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ ;
assign __auxvar5__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar5__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ ;
assign __auxvar6__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar6__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ ;
assign __auxvar7__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar7__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ ;
assign __auxvar8__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar8__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ ;
assign __auxvar9__recorder_sn_cond = ((monitor_s3)&&((__START__)||(__STARTED__)))&&(!(__ENDED__)) ;
assign __auxvar9__recorder_sn_value = RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ ;
assign __auxvar0__delay_d_0 = monitor_s4 ;
assign end_of_pipeline = (monitor_s4)&&(~(__auxvar0__delay)) ;
assign monitor_s1 = ((RTL__DOT__stage1_rg_full)&(~(monitor_s1_already)))&(__START__) ;
assign s2_enter = ((RTL__DOT__s1_to_s2$D_IN)&(RTL__DOT__s1_to_s2$EN))&(monitor_s1) ;
assign s2_exit = (RTL__DOT__s2_to_s3$D_IN)&(RTL__DOT__s2_to_s3$EN) ;
assign s3_enter = ((RTL__DOT__s2_to_s3$D_IN)&(RTL__DOT__s2_to_s3$EN))&(monitor_s2) ;
assign s3_exit = (RTL__DOT__s3_deq$EN)&(RTL__DOT__s3_deq$D_IN) ;
assign s4_enter = (monitor_s3)&&(RTL__DOT__rg_retiring$EN) ;
assign monitor_s1_already_enter_cond = (monitor_s1)&&(s2_enter) ;
assign monitor_s2_enter_cond = s2_enter ;
assign monitor_s2_exit_cond = s2_exit ;
assign monitor_s3_enter_cond = s3_enter ;
assign monitor_s3_exit_cond = s3_exit ;
assign monitor_s4_enter_cond = s4_enter ;
assign mem_req_addr = __auxvar33__recorder ;
assign mem_req_en = __auxvar34__recorder ;
assign mem_req_funct3 = __auxvar35__recorder ;
assign mem_req_op = __auxvar36__recorder ;
assign mem_req_rd_data = __auxvar37__recorder ;
assign mem_req_wd_data = __auxvar38__recorder ;
assign input_map_assume___p0__ = (!(__START__))||((__ILA_I_inst)==(RTL__DOT__near_mem$imem_instr)) ;
assign invariant_assume__p1__ = !(((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p2__ = !(((RTL__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p3__ = !(((RTL__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p4__ = !(((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p5__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p6__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p7__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p8__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p9__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p10__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p11__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p12__ = !(((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg)==(0))) ;
assign invariant_assume__p13__ = !(((RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p14__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p15__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p16__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p17__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg)==(0))) ;
assign invariant_assume__p18__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p19__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg)==(0))) ;
assign invariant_assume__p20__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg)==(0))) ;
assign invariant_assume__p21__ = !(((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg)==(0))&&((RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg)==(0))) ;
assign invariant_assume__p22__ = !(((RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage1_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p23__ = !(((RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage1_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p24__ = !(((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage2_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p25__ = !(((RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage2_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p26__ = !(((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(0))&&((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(0))) ;
assign invariant_assume__p27__ = !(((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(0))&&((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(0))) ;
assign invariant_assume__p28__ = ((((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage3_rg_full)==(1'b1))))&&((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__f_reset_reqs__DOT__full_reg)==(1'b0)))))&&(((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage2_rg_full)==(1'b1)))) ;
assign invariant_assume__p29__ = ((!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b1))))&&((RTL__DOT__stage2_f_reset_reqs__DOT__full_reg)==(1'b1)) ;
assign invariant_assume__p30__ = (((!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1)))||(!((RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(1'b0))))&&((((!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1)))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(1'b0)))) ;
assign invariant_assume__p31__ = (((((((((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b1))))||(!((RTL__DOT__rg_run_on_reset)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!(RTL__DOT__stage2_rg_stage2[101:101])))||((RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr[4:4])==(1'b1)))||(!((RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa[4:4])==(1'b1))))&&(!((RTL__DOT__csr_regfile__DOT__rg_nmi)==(1'b1))))&&(((!((RTL__DOT__rg_state[0:0])==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b0)))))&&(((((((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b1))||(!(RTL__DOT__rg_trap_instr[22:22])))||(!(RTL__DOT__rg_trap_instr[20:20])))||(!(RTL__DOT__rg_trap_instr[26:26])))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__csr_regfile__DOT__rg_state)==(1'b0)))))&&(((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__rg_run_on_reset)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b0)))) ;
assign invariant_assume__p32__ = (((((!((RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg)==(1'b0)))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__full_reg)==(1'b0))))&&(((((!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0)))||(!((RTL__DOT__rg_state[0:0])==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(RTL__DOT__rg_run_on_reset)))&&(((((((!((RTL__DOT__stage2_rg_full)==(1'b1)))||(!((RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg)==(1'b0))))||(!((RTL__DOT__rg_state[0:0])==(1'b1))))||(!((RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg)==(1'b1))))||(!((RTL__DOT__stage3_f_reset_rsps__DOT__full_reg)==(1'b1))))||(RTL__DOT__stage2_rg_stage2[168:168]))||(!(RTL__DOT__rg_cur_priv[1:1]))) ;
assign issue_decode__p33__ = (!(__START__))||(__ILA_riscv_decode_of_ADD__) ;
assign issue_valid__p34__ = (!(__START__))||(__ILA_riscv_valid__) ;
assign noreset__p35__ = (!(__RESETED__))||(!(dummy_reset)) ;
assign post_value_holder__p36__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar10__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar10__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)) ;
assign post_value_holder__p37__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar11__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar11__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)) ;
assign post_value_holder__p38__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar12__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar12__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)) ;
assign post_value_holder__p39__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar13__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar13__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)) ;
assign post_value_holder__p40__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar14__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar14__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)) ;
assign post_value_holder__p41__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar15__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar15__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)) ;
assign post_value_holder__p42__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar16__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar16__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)) ;
assign post_value_holder__p43__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar17__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar17__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)) ;
assign post_value_holder__p44__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar18__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar18__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)) ;
assign post_value_holder__p45__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar19__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar19__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)) ;
assign post_value_holder__p46__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar1__recorder_sn_condmet)))&&(monitor_s2)))||((__auxvar1__recorder)==(RTL__DOT__near_mem$imem_pc)) ;
assign post_value_holder__p47__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar20__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar20__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)) ;
assign post_value_holder__p48__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar21__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar21__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)) ;
assign post_value_holder__p49__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar22__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar22__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)) ;
assign post_value_holder__p50__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar23__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar23__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)) ;
assign post_value_holder__p51__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar24__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar24__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)) ;
assign post_value_holder__p52__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar25__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar25__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)) ;
assign post_value_holder__p53__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar26__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar26__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)) ;
assign post_value_holder__p54__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar27__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar27__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)) ;
assign post_value_holder__p55__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar28__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar28__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)) ;
assign post_value_holder__p56__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar29__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar29__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)) ;
assign post_value_holder__p57__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar2__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar2__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)) ;
assign post_value_holder__p58__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar30__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar30__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)) ;
assign post_value_holder__p59__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar31__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar31__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)) ;
assign post_value_holder__p60__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar32__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar32__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)) ;
assign post_value_holder__p61__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar33__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar33__recorder)==(RTL__DOT__near_mem$dmem_req_addr)) ;
assign post_value_holder__p62__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar34__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar34__recorder)==(RTL__DOT__near_mem$EN_dmem_req)) ;
assign post_value_holder__p63__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar35__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar35__recorder)==(RTL__DOT__near_mem$dmem_req_f3)) ;
assign post_value_holder__p64__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar36__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar36__recorder)==(RTL__DOT__near_mem$dmem_req_op)) ;
assign post_value_holder__p65__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar37__recorder_sn_condmet)))&&(monitor_s2)))||((__auxvar37__recorder)==(RTL__DOT__near_mem$dmem_word64[31:0])) ;
assign post_value_holder__p66__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar38__recorder_sn_condmet)))&&(monitor_s1)))||((__auxvar38__recorder)==(RTL__DOT__near_mem$dmem_req_store_value[31:0])) ;
assign post_value_holder__p67__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar3__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar3__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)) ;
assign post_value_holder__p68__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar4__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar4__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)) ;
assign post_value_holder__p69__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar5__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar5__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)) ;
assign post_value_holder__p70__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar6__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar6__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)) ;
assign post_value_holder__p71__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar7__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar7__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)) ;
assign post_value_holder__p72__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar8__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar8__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)) ;
assign post_value_holder__p73__ = (!((((__START__)||(__STARTED__))&&(!(__auxvar9__recorder_sn_condmet)))&&(monitor_s3)))||((__auxvar9__recorder)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)) ;
assign rfassumptions__p74__ = (__ILA_SO_pc[1:0])==(2'b00) ;
assign rfassumptions__p75__ = (RTL__DOT__near_mem$imem_pc[1:0])==(2'b00) ;
assign rfassumptions__p76__ = (!(monitor_s2))||((RTL__DOT__near_mem$dmem_exc)==(0)) ;
assign variable_map_assume___p77__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_load_en)))||((__ILA_SO_load_addr)==(mem_req_addr))) ;
assign variable_map_assume___p78__ = (!(__START__))||((!((__START__)&&(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0)))))||((__ILA_SO_load_data)==(mem_req_rd_data))) ;
assign variable_map_assume___p79__ = (!(__START__))||((!(__IEND__))||((__ILA_SO_load_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0))))) ;
assign variable_map_assume___p80__ = (!(__START__))||(((((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))||(((mem_req_funct3)==(0))||((mem_req_funct3)==(4))))&&((!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2)))))||(((mem_req_funct3)==(1))||((mem_req_funct3)==(5)))))&&((!(((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(4)))))||(((mem_req_funct3)==(2))||((mem_req_funct3)==(6)))))&&((!((((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(!(((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(1))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(4))))))&&(((__IEND__)&&(__ILA_SO_load_en))&&((__ILA_SO_load_size)==(8)))))||((mem_req_funct3)==(3)))) ;
assign variable_map_assume___p81__ = (!(__START__))||(((!(__START__))||((__ILA_SO_pc)==(RTL__DOT__near_mem$imem_pc)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_pc)==(__auxvar1__recorder)))) ;
assign variable_map_assume___p82__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_store_en)))||((__ILA_SO_store_addr)==(mem_req_addr))) ;
assign variable_map_assume___p83__ = (!(__START__))||((!((__IEND__)&&(__ILA_SO_store_en)))||((__ILA_SO_store_data)==(mem_req_wd_data))) ;
assign variable_map_assume___p84__ = (!(__START__))||((!(__IEND__))||((__ILA_SO_store_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b1))))) ;
assign variable_map_assume___p85__ = (!(__START__))||(((((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))||(((mem_req_funct3)==(0))||((mem_req_funct3)==(4))))&&((!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2)))))||(((mem_req_funct3)==(1))||((mem_req_funct3)==(5)))))&&((!(((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(4)))))||(((mem_req_funct3)==(2))||((mem_req_funct3)==(6)))))&&((!((((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(!(((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(!((!(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(1))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(2))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(4))))))&&(((__IEND__)&&(__ILA_SO_store_en))&&((__ILA_SO_store_size)==(8)))))||((mem_req_funct3)==(3)))) ;
assign variable_map_assume___p86__ = (!(__START__))||((__ILA_SO_x0)==(0)) ;
assign variable_map_assume___p87__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x1)==(__auxvar2__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x1)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)))) ;
assign variable_map_assume___p88__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x10)==(__auxvar3__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x10)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)))) ;
assign variable_map_assume___p89__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x11)==(__auxvar4__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x11)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)))) ;
assign variable_map_assume___p90__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x12)==(__auxvar5__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x12)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)))) ;
assign variable_map_assume___p91__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x13)==(__auxvar6__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x13)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)))) ;
assign variable_map_assume___p92__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x14)==(__auxvar7__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x14)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)))) ;
assign variable_map_assume___p93__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x15)==(__auxvar8__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x15)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)))) ;
assign variable_map_assume___p94__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x16)==(__auxvar9__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x16)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)))) ;
assign variable_map_assume___p95__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x17)==(__auxvar10__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x17)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)))) ;
assign variable_map_assume___p96__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x18)==(__auxvar11__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x18)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)))) ;
assign variable_map_assume___p97__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x19)==(__auxvar12__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x19)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)))) ;
assign variable_map_assume___p98__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x2)==(__auxvar13__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x2)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)))) ;
assign variable_map_assume___p99__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x20)==(__auxvar14__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x20)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)))) ;
assign variable_map_assume___p100__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x21)==(__auxvar15__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x21)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)))) ;
assign variable_map_assume___p101__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x22)==(__auxvar16__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x22)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)))) ;
assign variable_map_assume___p102__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x23)==(__auxvar17__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x23)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)))) ;
assign variable_map_assume___p103__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x24)==(__auxvar18__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x24)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)))) ;
assign variable_map_assume___p104__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x25)==(__auxvar19__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x25)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)))) ;
assign variable_map_assume___p105__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x26)==(__auxvar20__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x26)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)))) ;
assign variable_map_assume___p106__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x27)==(__auxvar21__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x27)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)))) ;
assign variable_map_assume___p107__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x28)==(__auxvar22__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x28)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)))) ;
assign variable_map_assume___p108__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x29)==(__auxvar23__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x29)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)))) ;
assign variable_map_assume___p109__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x3)==(__auxvar24__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x3)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)))) ;
assign variable_map_assume___p110__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x30)==(__auxvar25__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x30)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)))) ;
assign variable_map_assume___p111__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x31)==(__auxvar26__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x31)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)))) ;
assign variable_map_assume___p112__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x4)==(__auxvar27__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x4)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)))) ;
assign variable_map_assume___p113__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x5)==(__auxvar28__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x5)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)))) ;
assign variable_map_assume___p114__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x6)==(__auxvar29__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x6)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)))) ;
assign variable_map_assume___p115__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x7)==(__auxvar30__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x7)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)))) ;
assign variable_map_assume___p116__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x8)==(__auxvar31__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x8)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)))) ;
assign variable_map_assume___p117__ = (!(__START__))||(((!(__START__))||((__ILA_SO_x9)==(__auxvar32__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x9)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)))) ;
assign variable_map_assert__p118__ = (!(__IEND__))||((!(__IEND__))||((__ILA_SO_load_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b0))))) ;
assign variable_map_assert__p119__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_pc)==(RTL__DOT__near_mem$imem_pc)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_pc)==(__auxvar1__recorder)))) ;
assign variable_map_assert__p120__ = (!(__IEND__))||((!(__IEND__))||((__ILA_SO_store_en)==(((mem_req_en)==(1'b1))&&((mem_req_op)==(1'b1))))) ;
assign variable_map_assert__p121__ = (!(__IEND__))||((__ILA_SO_x0)==(0)) ;
assign variable_map_assert__p122__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x1)==(__auxvar2__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x1)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_)))) ;
assign variable_map_assert__p123__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x10)==(__auxvar3__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x10)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_)))) ;
assign variable_map_assert__p124__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x11)==(__auxvar4__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x11)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_)))) ;
assign variable_map_assert__p125__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x12)==(__auxvar5__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x12)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_)))) ;
assign variable_map_assert__p126__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x13)==(__auxvar6__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x13)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_)))) ;
assign variable_map_assert__p127__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x14)==(__auxvar7__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x14)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_)))) ;
assign variable_map_assert__p128__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x15)==(__auxvar8__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x15)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_)))) ;
assign variable_map_assert__p129__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x16)==(__auxvar9__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x16)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_)))) ;
assign variable_map_assert__p130__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x17)==(__auxvar10__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x17)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_)))) ;
assign variable_map_assert__p131__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x18)==(__auxvar11__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x18)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_)))) ;
assign variable_map_assert__p132__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x19)==(__auxvar12__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x19)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_)))) ;
assign variable_map_assert__p133__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x2)==(__auxvar13__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x2)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_)))) ;
assign variable_map_assert__p134__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x20)==(__auxvar14__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x20)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_)))) ;
assign variable_map_assert__p135__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x21)==(__auxvar15__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x21)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_)))) ;
assign variable_map_assert__p136__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x22)==(__auxvar16__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x22)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_)))) ;
assign variable_map_assert__p137__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x23)==(__auxvar17__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x23)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_)))) ;
assign variable_map_assert__p138__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x24)==(__auxvar18__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x24)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_)))) ;
assign variable_map_assert__p139__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x25)==(__auxvar19__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x25)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_)))) ;
assign variable_map_assert__p140__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x26)==(__auxvar20__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x26)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_)))) ;
assign variable_map_assert__p141__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x27)==(__auxvar21__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x27)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_)))) ;
assign variable_map_assert__p142__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x28)==(__auxvar22__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x28)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_)))) ;
assign variable_map_assert__p143__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x29)==(__auxvar23__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x29)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_)))) ;
assign variable_map_assert__p144__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x3)==(__auxvar24__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x3)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_)))) ;
assign variable_map_assert__p145__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x30)==(__auxvar25__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x30)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_)))) ;
assign variable_map_assert__p146__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x31)==(__auxvar26__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x31)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_)))) ;
assign variable_map_assert__p147__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x4)==(__auxvar27__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x4)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_)))) ;
assign variable_map_assert__p148__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x5)==(__auxvar28__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x5)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_)))) ;
assign variable_map_assert__p149__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x6)==(__auxvar29__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x6)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_)))) ;
assign variable_map_assert__p150__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x7)==(__auxvar30__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x7)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_)))) ;
assign variable_map_assert__p151__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x8)==(__auxvar31__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x8)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_)))) ;
assign variable_map_assert__p152__ = (!(__IEND__))||(((!(__START__))||((__ILA_SO_x9)==(__auxvar32__recorder)))&&((!((!(__START__))&&(__IEND__)))||((__ILA_SO_x9)==(RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_)))) ;
assign post_value_holder_overly_constrained__p153__ = (!((__auxvar10__recorder_sn_condmet)&&(__auxvar10__recorder_sn_cond)))||((__auxvar10__recorder_sn_value)==(__auxvar10__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p154__ = (!((__auxvar11__recorder_sn_condmet)&&(__auxvar11__recorder_sn_cond)))||((__auxvar11__recorder_sn_value)==(__auxvar11__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p155__ = (!((__auxvar12__recorder_sn_condmet)&&(__auxvar12__recorder_sn_cond)))||((__auxvar12__recorder_sn_value)==(__auxvar12__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p156__ = (!((__auxvar13__recorder_sn_condmet)&&(__auxvar13__recorder_sn_cond)))||((__auxvar13__recorder_sn_value)==(__auxvar13__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p157__ = (!((__auxvar14__recorder_sn_condmet)&&(__auxvar14__recorder_sn_cond)))||((__auxvar14__recorder_sn_value)==(__auxvar14__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p158__ = (!((__auxvar15__recorder_sn_condmet)&&(__auxvar15__recorder_sn_cond)))||((__auxvar15__recorder_sn_value)==(__auxvar15__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p159__ = (!((__auxvar16__recorder_sn_condmet)&&(__auxvar16__recorder_sn_cond)))||((__auxvar16__recorder_sn_value)==(__auxvar16__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p160__ = (!((__auxvar17__recorder_sn_condmet)&&(__auxvar17__recorder_sn_cond)))||((__auxvar17__recorder_sn_value)==(__auxvar17__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p161__ = (!((__auxvar18__recorder_sn_condmet)&&(__auxvar18__recorder_sn_cond)))||((__auxvar18__recorder_sn_value)==(__auxvar18__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p162__ = (!((__auxvar19__recorder_sn_condmet)&&(__auxvar19__recorder_sn_cond)))||((__auxvar19__recorder_sn_value)==(__auxvar19__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p163__ = (!((__auxvar1__recorder_sn_condmet)&&(__auxvar1__recorder_sn_cond)))||((__auxvar1__recorder_sn_value)==(__auxvar1__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p164__ = (!((__auxvar20__recorder_sn_condmet)&&(__auxvar20__recorder_sn_cond)))||((__auxvar20__recorder_sn_value)==(__auxvar20__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p165__ = (!((__auxvar21__recorder_sn_condmet)&&(__auxvar21__recorder_sn_cond)))||((__auxvar21__recorder_sn_value)==(__auxvar21__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p166__ = (!((__auxvar22__recorder_sn_condmet)&&(__auxvar22__recorder_sn_cond)))||((__auxvar22__recorder_sn_value)==(__auxvar22__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p167__ = (!((__auxvar23__recorder_sn_condmet)&&(__auxvar23__recorder_sn_cond)))||((__auxvar23__recorder_sn_value)==(__auxvar23__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p168__ = (!((__auxvar24__recorder_sn_condmet)&&(__auxvar24__recorder_sn_cond)))||((__auxvar24__recorder_sn_value)==(__auxvar24__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p169__ = (!((__auxvar25__recorder_sn_condmet)&&(__auxvar25__recorder_sn_cond)))||((__auxvar25__recorder_sn_value)==(__auxvar25__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p170__ = (!((__auxvar26__recorder_sn_condmet)&&(__auxvar26__recorder_sn_cond)))||((__auxvar26__recorder_sn_value)==(__auxvar26__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p171__ = (!((__auxvar27__recorder_sn_condmet)&&(__auxvar27__recorder_sn_cond)))||((__auxvar27__recorder_sn_value)==(__auxvar27__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p172__ = (!((__auxvar28__recorder_sn_condmet)&&(__auxvar28__recorder_sn_cond)))||((__auxvar28__recorder_sn_value)==(__auxvar28__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p173__ = (!((__auxvar29__recorder_sn_condmet)&&(__auxvar29__recorder_sn_cond)))||((__auxvar29__recorder_sn_value)==(__auxvar29__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p174__ = (!((__auxvar2__recorder_sn_condmet)&&(__auxvar2__recorder_sn_cond)))||((__auxvar2__recorder_sn_value)==(__auxvar2__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p175__ = (!((__auxvar30__recorder_sn_condmet)&&(__auxvar30__recorder_sn_cond)))||((__auxvar30__recorder_sn_value)==(__auxvar30__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p176__ = (!((__auxvar31__recorder_sn_condmet)&&(__auxvar31__recorder_sn_cond)))||((__auxvar31__recorder_sn_value)==(__auxvar31__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p177__ = (!((__auxvar32__recorder_sn_condmet)&&(__auxvar32__recorder_sn_cond)))||((__auxvar32__recorder_sn_value)==(__auxvar32__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p178__ = (!((__auxvar33__recorder_sn_condmet)&&(__auxvar33__recorder_sn_cond)))||((__auxvar33__recorder_sn_value)==(__auxvar33__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p179__ = (!((__auxvar34__recorder_sn_condmet)&&(__auxvar34__recorder_sn_cond)))||((__auxvar34__recorder_sn_value)==(__auxvar34__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p180__ = (!((__auxvar35__recorder_sn_condmet)&&(__auxvar35__recorder_sn_cond)))||((__auxvar35__recorder_sn_value)==(__auxvar35__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p181__ = (!((__auxvar36__recorder_sn_condmet)&&(__auxvar36__recorder_sn_cond)))||((__auxvar36__recorder_sn_value)==(__auxvar36__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p182__ = (!((__auxvar37__recorder_sn_condmet)&&(__auxvar37__recorder_sn_cond)))||((__auxvar37__recorder_sn_value)==(__auxvar37__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p183__ = (!((__auxvar38__recorder_sn_condmet)&&(__auxvar38__recorder_sn_cond)))||((__auxvar38__recorder_sn_value)==(__auxvar38__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p184__ = (!((__auxvar3__recorder_sn_condmet)&&(__auxvar3__recorder_sn_cond)))||((__auxvar3__recorder_sn_value)==(__auxvar3__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p185__ = (!((__auxvar4__recorder_sn_condmet)&&(__auxvar4__recorder_sn_cond)))||((__auxvar4__recorder_sn_value)==(__auxvar4__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p186__ = (!((__auxvar5__recorder_sn_condmet)&&(__auxvar5__recorder_sn_cond)))||((__auxvar5__recorder_sn_value)==(__auxvar5__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p187__ = (!((__auxvar6__recorder_sn_condmet)&&(__auxvar6__recorder_sn_cond)))||((__auxvar6__recorder_sn_value)==(__auxvar6__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p188__ = (!((__auxvar7__recorder_sn_condmet)&&(__auxvar7__recorder_sn_cond)))||((__auxvar7__recorder_sn_value)==(__auxvar7__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p189__ = (!((__auxvar8__recorder_sn_condmet)&&(__auxvar8__recorder_sn_cond)))||((__auxvar8__recorder_sn_value)==(__auxvar8__recorder_sn_vhold)) ;
assign post_value_holder_overly_constrained__p190__ = (!((__auxvar9__recorder_sn_condmet)&&(__auxvar9__recorder_sn_cond)))||((__auxvar9__recorder_sn_value)==(__auxvar9__recorder_sn_vhold)) ;
assign post_value_holder_triggered__p191__ = (!(__IEND__))||((__auxvar10__recorder_sn_condmet)||(__auxvar10__recorder_sn_cond)) ;
assign post_value_holder_triggered__p192__ = (!(__IEND__))||((__auxvar11__recorder_sn_condmet)||(__auxvar11__recorder_sn_cond)) ;
assign post_value_holder_triggered__p193__ = (!(__IEND__))||((__auxvar12__recorder_sn_condmet)||(__auxvar12__recorder_sn_cond)) ;
assign post_value_holder_triggered__p194__ = (!(__IEND__))||((__auxvar13__recorder_sn_condmet)||(__auxvar13__recorder_sn_cond)) ;
assign post_value_holder_triggered__p195__ = (!(__IEND__))||((__auxvar14__recorder_sn_condmet)||(__auxvar14__recorder_sn_cond)) ;
assign post_value_holder_triggered__p196__ = (!(__IEND__))||((__auxvar15__recorder_sn_condmet)||(__auxvar15__recorder_sn_cond)) ;
assign post_value_holder_triggered__p197__ = (!(__IEND__))||((__auxvar16__recorder_sn_condmet)||(__auxvar16__recorder_sn_cond)) ;
assign post_value_holder_triggered__p198__ = (!(__IEND__))||((__auxvar17__recorder_sn_condmet)||(__auxvar17__recorder_sn_cond)) ;
assign post_value_holder_triggered__p199__ = (!(__IEND__))||((__auxvar18__recorder_sn_condmet)||(__auxvar18__recorder_sn_cond)) ;
assign post_value_holder_triggered__p200__ = (!(__IEND__))||((__auxvar19__recorder_sn_condmet)||(__auxvar19__recorder_sn_cond)) ;
assign post_value_holder_triggered__p201__ = (!(__IEND__))||((__auxvar1__recorder_sn_condmet)||(__auxvar1__recorder_sn_cond)) ;
assign post_value_holder_triggered__p202__ = (!(__IEND__))||((__auxvar20__recorder_sn_condmet)||(__auxvar20__recorder_sn_cond)) ;
assign post_value_holder_triggered__p203__ = (!(__IEND__))||((__auxvar21__recorder_sn_condmet)||(__auxvar21__recorder_sn_cond)) ;
assign post_value_holder_triggered__p204__ = (!(__IEND__))||((__auxvar22__recorder_sn_condmet)||(__auxvar22__recorder_sn_cond)) ;
assign post_value_holder_triggered__p205__ = (!(__IEND__))||((__auxvar23__recorder_sn_condmet)||(__auxvar23__recorder_sn_cond)) ;
assign post_value_holder_triggered__p206__ = (!(__IEND__))||((__auxvar24__recorder_sn_condmet)||(__auxvar24__recorder_sn_cond)) ;
assign post_value_holder_triggered__p207__ = (!(__IEND__))||((__auxvar25__recorder_sn_condmet)||(__auxvar25__recorder_sn_cond)) ;
assign post_value_holder_triggered__p208__ = (!(__IEND__))||((__auxvar26__recorder_sn_condmet)||(__auxvar26__recorder_sn_cond)) ;
assign post_value_holder_triggered__p209__ = (!(__IEND__))||((__auxvar27__recorder_sn_condmet)||(__auxvar27__recorder_sn_cond)) ;
assign post_value_holder_triggered__p210__ = (!(__IEND__))||((__auxvar28__recorder_sn_condmet)||(__auxvar28__recorder_sn_cond)) ;
assign post_value_holder_triggered__p211__ = (!(__IEND__))||((__auxvar29__recorder_sn_condmet)||(__auxvar29__recorder_sn_cond)) ;
assign post_value_holder_triggered__p212__ = (!(__IEND__))||((__auxvar2__recorder_sn_condmet)||(__auxvar2__recorder_sn_cond)) ;
assign post_value_holder_triggered__p213__ = (!(__IEND__))||((__auxvar30__recorder_sn_condmet)||(__auxvar30__recorder_sn_cond)) ;
assign post_value_holder_triggered__p214__ = (!(__IEND__))||((__auxvar31__recorder_sn_condmet)||(__auxvar31__recorder_sn_cond)) ;
assign post_value_holder_triggered__p215__ = (!(__IEND__))||((__auxvar32__recorder_sn_condmet)||(__auxvar32__recorder_sn_cond)) ;
assign post_value_holder_triggered__p216__ = (!(__IEND__))||((__auxvar33__recorder_sn_condmet)||(__auxvar33__recorder_sn_cond)) ;
assign post_value_holder_triggered__p217__ = (!(__IEND__))||((__auxvar34__recorder_sn_condmet)||(__auxvar34__recorder_sn_cond)) ;
assign post_value_holder_triggered__p218__ = (!(__IEND__))||((__auxvar35__recorder_sn_condmet)||(__auxvar35__recorder_sn_cond)) ;
assign post_value_holder_triggered__p219__ = (!(__IEND__))||((__auxvar36__recorder_sn_condmet)||(__auxvar36__recorder_sn_cond)) ;
assign post_value_holder_triggered__p220__ = (!(__IEND__))||((__auxvar37__recorder_sn_condmet)||(__auxvar37__recorder_sn_cond)) ;
assign post_value_holder_triggered__p221__ = (!(__IEND__))||((__auxvar38__recorder_sn_condmet)||(__auxvar38__recorder_sn_cond)) ;
assign post_value_holder_triggered__p222__ = (!(__IEND__))||((__auxvar3__recorder_sn_condmet)||(__auxvar3__recorder_sn_cond)) ;
assign post_value_holder_triggered__p223__ = (!(__IEND__))||((__auxvar4__recorder_sn_condmet)||(__auxvar4__recorder_sn_cond)) ;
assign post_value_holder_triggered__p224__ = (!(__IEND__))||((__auxvar5__recorder_sn_condmet)||(__auxvar5__recorder_sn_cond)) ;
assign post_value_holder_triggered__p225__ = (!(__IEND__))||((__auxvar6__recorder_sn_condmet)||(__auxvar6__recorder_sn_cond)) ;
assign post_value_holder_triggered__p226__ = (!(__IEND__))||((__auxvar7__recorder_sn_condmet)||(__auxvar7__recorder_sn_cond)) ;
assign post_value_holder_triggered__p227__ = (!(__IEND__))||((__auxvar8__recorder_sn_condmet)||(__auxvar8__recorder_sn_cond)) ;
assign post_value_holder_triggered__p228__ = (!(__IEND__))||((__auxvar9__recorder_sn_condmet)||(__auxvar9__recorder_sn_cond)) ;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem$dmem_req_op;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__rg_trap_instr;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire[63:0] RTL___RTL__DOT__near_mem$dmem_req_store_value;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire[63:0] RTL___RTL__DOT__near_mem$dmem_word64;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__s1_to_s2$D_IN;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire RTL___RTL__DOT__stage2_rg_full;
    wire RTL___RTL__DOT__csr_regfile__DOT__rg_state;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___RTL__DOT__stage1_rg_full;
    wire RTL___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire RTL___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__rg_run_on_reset;
    wire RTL___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___RTL__DOT__s2_to_s3$EN;
    wire[2:0] RTL___RTL__DOT__near_mem$dmem_req_f3;
    wire RTL___RTL__DOT__s1_to_s2$EN;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire RTL___RTL__DOT__s3_deq$EN;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire[3:0] RTL___RTL__DOT__rg_state;
    wire RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___RTL__DOT__rg_retiring$EN;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___RTL__DOT__s2_to_s3$D_IN;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire RTL___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__stage3_rg_full;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire[168:0] RTL___RTL__DOT__stage2_rg_stage2;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__csr_regfile__DOT__rg_nmi;
    wire[31:0] RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL___RTL__DOT__near_mem$EN_dmem_req;
    wire RTL___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire[1:0] RTL___RTL__DOT__rg_cur_priv;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire RTL___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__near_mem$dmem_req_addr;
    wire[31:0] RTL___RTL__DOT__near_mem$imem_instr;
    wire RTL___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire[31:0] RTL___RTL__DOT__near_mem$imem_pc;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem$dmem_exc;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___RTL__DOT__s3_deq$D_IN;
    wire RTL___CLK;
    wire RTL___RST_N;
    wire RTL___hart0_server_reset_request_put;
    wire RTL___EN_hart0_server_reset_request_put;
    wire RTL___EN_hart0_server_reset_response_get;
    wire RTL___imem_master_awready;
    wire RTL___imem_master_wready;
    wire RTL___imem_master_bvalid;
    wire[3:0] RTL___imem_master_bid;
    wire[1:0] RTL___imem_master_bresp;
    wire RTL___imem_master_arready;
    wire RTL___imem_master_rvalid;
    wire[3:0] RTL___imem_master_rid;
    wire[63:0] RTL___imem_master_rdata;
    wire[1:0] RTL___imem_master_rresp;
    wire RTL___imem_master_rlast;
    wire RTL___dmem_master_awready;
    wire RTL___dmem_master_wready;
    wire RTL___dmem_master_bvalid;
    wire[3:0] RTL___dmem_master_bid;
    wire[1:0] RTL___dmem_master_bresp;
    wire RTL___dmem_master_arready;
    wire RTL___dmem_master_rvalid;
    wire[3:0] RTL___dmem_master_rid;
    wire[63:0] RTL___dmem_master_rdata;
    wire[1:0] RTL___dmem_master_rresp;
    wire RTL___dmem_master_rlast;
    wire RTL___m_external_interrupt_req_set_not_clear;
    wire RTL___s_external_interrupt_req_set_not_clear;
    wire RTL___software_interrupt_req_set_not_clear;
    wire RTL___timer_interrupt_req_set_not_clear;
    wire RTL___nmi_req_set_not_clear;
    wire[3:0] RTL___set_verbosity_verbosity;
    wire[63:0] RTL___set_verbosity_logdelay;
    wire RTL___EN_set_verbosity;

    wire[63:0] RTL___dmem_master_araddr , RTL___dmem_master_awaddr , RTL___dmem_master_wdata , RTL___imem_master_araddr , RTL___imem_master_awaddr , RTL___imem_master_wdata ; 
    wire[7:0] RTL___dmem_master_arlen , RTL___dmem_master_awlen , RTL___dmem_master_wstrb , RTL___imem_master_arlen , RTL___imem_master_awlen , RTL___imem_master_wstrb ; 
    wire[3:0] RTL___dmem_master_arcache , RTL___dmem_master_arid , RTL___dmem_master_arqos , RTL___dmem_master_arregion , RTL___dmem_master_awcache , RTL___dmem_master_awid , RTL___dmem_master_awqos , RTL___dmem_master_awregion , RTL___imem_master_arcache , RTL___imem_master_arid , RTL___imem_master_arqos , RTL___imem_master_arregion , RTL___imem_master_awcache , RTL___imem_master_awid , RTL___imem_master_awqos , RTL___imem_master_awregion ; 
    wire[2:0] RTL___dmem_master_arprot , RTL___dmem_master_arsize , RTL___dmem_master_awprot , RTL___dmem_master_awsize , RTL___imem_master_arprot , RTL___imem_master_arsize , RTL___imem_master_awprot , RTL___imem_master_awsize ; 
    wire[1:0] RTL___dmem_master_arburst , RTL___dmem_master_awburst , RTL___imem_master_arburst , RTL___imem_master_awburst ; 
    wire RTL___RDY_hart0_server_reset_request_put , RTL___RDY_hart0_server_reset_response_get , RTL___RDY_set_verbosity , RTL___dmem_master_arlock , RTL___dmem_master_arvalid , RTL___dmem_master_awlock , RTL___dmem_master_awvalid , RTL___dmem_master_bready , RTL___dmem_master_rready , RTL___dmem_master_wlast , RTL___dmem_master_wvalid , RTL___hart0_server_reset_response_get , RTL___imem_master_arlock , RTL___imem_master_arvalid , RTL___imem_master_awlock , RTL___imem_master_awvalid , RTL___imem_master_bready , RTL___imem_master_rready , RTL___imem_master_wlast , RTL___imem_master_wvalid ; reg[63:0] RTL___cfg_logdelay ; 
    wire[63:0] RTL___cfg_logdelay$D_IN ; 
    wire RTL___cfg_logdelay$EN ; reg[3:0] RTL___cfg_verbosity ; 
    wire[3:0] RTL___cfg_verbosity$D_IN ; 
    wire RTL___cfg_verbosity$EN ; reg[31:0] RTL___rg_csr_pc ; 
    wire[31:0] RTL___rg_csr_pc$D_IN ; 
    wire RTL___rg_csr_pc$EN ; reg[31:0] RTL___rg_csr_val1 ; 
    wire[31:0] RTL___rg_csr_val1$D_IN ; 
    wire RTL___rg_csr_val1$EN ; reg[1:0] RTL___rg_cur_priv ; reg[1:0] RTL___rg_cur_priv$D_IN ; 
    wire RTL___rg_cur_priv$EN ; 
    reg RTL___rg_mstatus_MXR ; 
    wire RTL___rg_mstatus_MXR$D_IN , RTL___rg_mstatus_MXR$EN ; reg[31:0] RTL___rg_next_pc ; reg[31:0] RTL___rg_next_pc$D_IN ; 
    wire RTL___rg_next_pc$EN ; 
    reg RTL___rg_retiring ; 
    wire RTL___rg_retiring$D_IN , RTL___rg_retiring$EN ; 
    reg RTL___rg_run_on_reset ; 
    wire RTL___rg_run_on_reset$D_IN , RTL___rg_run_on_reset$EN ; 
    reg RTL___rg_sstatus_SUM ; 
    wire RTL___rg_sstatus_SUM$D_IN , RTL___rg_sstatus_SUM$EN ; reg[63:0] RTL___rg_start_CPI_cycles ; 
    wire[63:0] RTL___rg_start_CPI_cycles$D_IN ; 
    wire RTL___rg_start_CPI_cycles$EN ; reg[63:0] RTL___rg_start_CPI_instrs ; 
    wire[63:0] RTL___rg_start_CPI_instrs$D_IN ; 
    wire RTL___rg_start_CPI_instrs$EN ; reg[3:0] RTL___rg_state ; reg[3:0] RTL___rg_state$D_IN ; 
    wire RTL___rg_state$EN ; reg[67:0] RTL___rg_trap_info ; reg[67:0] RTL___rg_trap_info$D_IN ; 
    wire RTL___rg_trap_info$EN ; reg[31:0] RTL___rg_trap_instr ; 
    wire[31:0] RTL___rg_trap_instr$D_IN ; 
    wire RTL___rg_trap_instr$EN ; 
    reg RTL___rg_trap_interrupt ; 
    wire RTL___rg_trap_interrupt$D_IN , RTL___rg_trap_interrupt$EN ; 
    reg RTL___s1_to_s2 ; 
    wire RTL___s1_to_s2$D_IN , RTL___s1_to_s2$EN ; 
    reg RTL___s2_to_s3 ; 
    wire RTL___s2_to_s3$D_IN , RTL___s2_to_s3$EN ; 
    reg RTL___s3_deq ; 
    wire RTL___s3_deq$D_IN , RTL___s3_deq$EN ; 
    reg RTL___stage1_rg_full ; 
    reg RTL___stage1_rg_full$D_IN ; 
    wire RTL___stage1_rg_full$EN ; 
    reg RTL___stage2_rg_full ; 
    reg RTL___stage2_rg_full$D_IN ; 
    wire RTL___stage2_rg_full$EN ; 
    reg RTL___stage2_rg_resetting ; 
    wire RTL___stage2_rg_resetting$D_IN , RTL___stage2_rg_resetting$EN ; reg[168:0] RTL___stage2_rg_stage2 ; 
    wire[168:0] RTL___stage2_rg_stage2$D_IN ; 
    wire RTL___stage2_rg_stage2$EN ; 
    reg RTL___stage3_rg_full ; 
    reg RTL___stage3_rg_full$D_IN ; 
    wire RTL___stage3_rg_full$EN ; reg[103:0] RTL___stage3_rg_stage3 ; 
    wire[103:0] RTL___stage3_rg_stage3$D_IN ; 
    wire RTL___stage3_rg_stage3$EN ; reg[1:0] RTL___csr_regfile$csr_ret_actions_from_priv ; 
    wire[97:0] RTL___csr_regfile$csr_trap_actions ; 
    wire[65:0] RTL___csr_regfile$csr_ret_actions ; 
    wire[63:0] RTL___csr_regfile$read_csr_mcycle , RTL___csr_regfile$read_csr_minstret ; 
    wire[32:0] RTL___csr_regfile$read_csr ; 
    wire[31:0] RTL___csr_regfile$csr_trap_actions_pc , RTL___csr_regfile$csr_trap_actions_xtval , RTL___csr_regfile$mav_csr_write_word , RTL___csr_regfile$read_mstatus , RTL___csr_regfile$read_satp ; 
    wire[27:0] RTL___csr_regfile$read_misa ; 
    wire[11:0] RTL___csr_regfile$access_permitted_1_csr_addr , RTL___csr_regfile$access_permitted_2_csr_addr , RTL___csr_regfile$csr_counter_read_fault_csr_addr , RTL___csr_regfile$mav_csr_write_csr_addr , RTL___csr_regfile$mav_read_csr_csr_addr , RTL___csr_regfile$read_csr_csr_addr , RTL___csr_regfile$read_csr_port2_csr_addr ; 
    wire[4:0] RTL___csr_regfile$interrupt_pending ; 
    wire[3:0] RTL___csr_regfile$csr_trap_actions_exc_code ; 
    wire[1:0] RTL___csr_regfile$access_permitted_1_priv , RTL___csr_regfile$access_permitted_2_priv , RTL___csr_regfile$csr_counter_read_fault_priv , RTL___csr_regfile$csr_trap_actions_from_priv , RTL___csr_regfile$interrupt_pending_cur_priv ; 
    wire RTL___csr_regfile$EN_csr_minstret_incr , RTL___csr_regfile$EN_csr_ret_actions , RTL___csr_regfile$EN_csr_trap_actions , RTL___csr_regfile$EN_debug , RTL___csr_regfile$EN_mav_csr_write , RTL___csr_regfile$EN_mav_read_csr , RTL___csr_regfile$EN_server_reset_request_put , RTL___csr_regfile$EN_server_reset_response_get , RTL___csr_regfile$RDY_server_reset_request_put , RTL___csr_regfile$RDY_server_reset_response_get , RTL___csr_regfile$access_permitted_1 , RTL___csr_regfile$access_permitted_1_read_not_write , RTL___csr_regfile$access_permitted_2 , RTL___csr_regfile$access_permitted_2_read_not_write , RTL___csr_regfile$csr_trap_actions_interrupt , RTL___csr_regfile$csr_trap_actions_nmi , RTL___csr_regfile$m_external_interrupt_req_set_not_clear , RTL___csr_regfile$nmi_pending , RTL___csr_regfile$nmi_req_set_not_clear , RTL___csr_regfile$s_external_interrupt_req_set_not_clear , RTL___csr_regfile$software_interrupt_req_set_not_clear , RTL___csr_regfile$timer_interrupt_req_set_not_clear , RTL___csr_regfile$wfi_resume ; 
    wire RTL___f_reset_reqs$CLR , RTL___f_reset_reqs$DEQ , RTL___f_reset_reqs$D_IN , RTL___f_reset_reqs$D_OUT , RTL___f_reset_reqs$EMPTY_N , RTL___f_reset_reqs$ENQ , RTL___f_reset_reqs$FULL_N ; 
    wire RTL___f_reset_rsps$CLR , RTL___f_reset_rsps$DEQ , RTL___f_reset_rsps$D_IN , RTL___f_reset_rsps$D_OUT , RTL___f_reset_rsps$EMPTY_N , RTL___f_reset_rsps$ENQ , RTL___f_reset_rsps$FULL_N ; 
    wire[31:0] RTL___gpr_regfile$read_rs1 , RTL___gpr_regfile$read_rs2 , RTL___gpr_regfile$write_rd_rd_val ; 
    wire[4:0] RTL___gpr_regfile$read_rs1_port2_rs1 , RTL___gpr_regfile$read_rs1_rs1 , RTL___gpr_regfile$read_rs2_rs2 , RTL___gpr_regfile$write_rd_rd ; 
    wire RTL___gpr_regfile$EN_server_reset_request_put , RTL___gpr_regfile$EN_server_reset_response_get , RTL___gpr_regfile$EN_write_rd , RTL___gpr_regfile$RDY_server_reset_request_put , RTL___gpr_regfile$RDY_server_reset_response_get ; reg[31:0] RTL___near_mem$imem_req_addr ; 
    wire[63:0] RTL___near_mem$dmem_master_araddr , RTL___near_mem$dmem_master_awaddr , RTL___near_mem$dmem_master_rdata , RTL___near_mem$dmem_master_wdata , RTL___near_mem$dmem_req_store_value , RTL___near_mem$dmem_word64 , RTL___near_mem$imem_master_araddr , RTL___near_mem$imem_master_awaddr , RTL___near_mem$imem_master_rdata , RTL___near_mem$imem_master_wdata ; 
    wire[31:0] RTL___near_mem$dmem_req_addr , RTL___near_mem$dmem_req_satp , RTL___near_mem$imem_instr , RTL___near_mem$imem_pc , RTL___near_mem$imem_req_satp , RTL___near_mem$imem_tval ; 
    wire[7:0] RTL___near_mem$dmem_master_arlen , RTL___near_mem$dmem_master_awlen , RTL___near_mem$dmem_master_wstrb , RTL___near_mem$imem_master_arlen , RTL___near_mem$imem_master_awlen , RTL___near_mem$imem_master_wstrb , RTL___near_mem$server_fence_request_put ; 
    wire[3:0] RTL___near_mem$dmem_exc_code , RTL___near_mem$dmem_master_arcache , RTL___near_mem$dmem_master_arid , RTL___near_mem$dmem_master_arqos , RTL___near_mem$dmem_master_arregion , RTL___near_mem$dmem_master_awcache , RTL___near_mem$dmem_master_awid , RTL___near_mem$dmem_master_awqos , RTL___near_mem$dmem_master_awregion , RTL___near_mem$dmem_master_bid , RTL___near_mem$dmem_master_rid , RTL___near_mem$imem_exc_code , RTL___near_mem$imem_master_arcache , RTL___near_mem$imem_master_arid , RTL___near_mem$imem_master_arqos , RTL___near_mem$imem_master_arregion , RTL___near_mem$imem_master_awcache , RTL___near_mem$imem_master_awid , RTL___near_mem$imem_master_awqos , RTL___near_mem$imem_master_awregion , RTL___near_mem$imem_master_bid , RTL___near_mem$imem_master_rid ; 
    wire[2:0] RTL___near_mem$dmem_master_arprot , RTL___near_mem$dmem_master_arsize , RTL___near_mem$dmem_master_awprot , RTL___near_mem$dmem_master_awsize , RTL___near_mem$dmem_req_f3 , RTL___near_mem$imem_master_arprot , RTL___near_mem$imem_master_arsize , RTL___near_mem$imem_master_awprot , RTL___near_mem$imem_master_awsize , RTL___near_mem$imem_req_f3 ; 
    wire[1:0] RTL___near_mem$dmem_master_arburst , RTL___near_mem$dmem_master_awburst , RTL___near_mem$dmem_master_bresp , RTL___near_mem$dmem_master_rresp , RTL___near_mem$dmem_req_priv , RTL___near_mem$imem_master_arburst , RTL___near_mem$imem_master_awburst , RTL___near_mem$imem_master_bresp , RTL___near_mem$imem_master_rresp , RTL___near_mem$imem_req_priv ; 
    wire RTL___near_mem$EN_dmem_req , RTL___near_mem$EN_imem_req , RTL___near_mem$EN_server_fence_i_request_put , RTL___near_mem$EN_server_fence_i_response_get , RTL___near_mem$EN_server_fence_request_put , RTL___near_mem$EN_server_fence_response_get , RTL___near_mem$EN_server_reset_request_put , RTL___near_mem$EN_server_reset_response_get , RTL___near_mem$EN_sfence_vma , RTL___near_mem$RDY_server_fence_i_request_put , RTL___near_mem$RDY_server_fence_i_response_get , RTL___near_mem$RDY_server_fence_request_put , RTL___near_mem$RDY_server_fence_response_get , RTL___near_mem$RDY_server_reset_request_put , RTL___near_mem$RDY_server_reset_response_get , RTL___near_mem$dmem_exc , RTL___near_mem$dmem_master_arlock , RTL___near_mem$dmem_master_arready , RTL___near_mem$dmem_master_arvalid , RTL___near_mem$dmem_master_awlock , RTL___near_mem$dmem_master_awready , RTL___near_mem$dmem_master_awvalid , RTL___near_mem$dmem_master_bready , RTL___near_mem$dmem_master_bvalid , RTL___near_mem$dmem_master_rlast , RTL___near_mem$dmem_master_rready , RTL___near_mem$dmem_master_rvalid , RTL___near_mem$dmem_master_wlast , RTL___near_mem$dmem_master_wready , RTL___near_mem$dmem_master_wvalid , RTL___near_mem$dmem_req_mstatus_MXR , RTL___near_mem$dmem_req_op , RTL___near_mem$dmem_req_sstatus_SUM , RTL___near_mem$dmem_valid , RTL___near_mem$imem_exc , RTL___near_mem$imem_is_i32_not_i16 , RTL___near_mem$imem_master_arlock , RTL___near_mem$imem_master_arready , RTL___near_mem$imem_master_arvalid , RTL___near_mem$imem_master_awlock , RTL___near_mem$imem_master_awready , RTL___near_mem$imem_master_awvalid , RTL___near_mem$imem_master_bready , RTL___near_mem$imem_master_bvalid , RTL___near_mem$imem_master_rlast , RTL___near_mem$imem_master_rready , RTL___near_mem$imem_master_rvalid , RTL___near_mem$imem_master_wlast , RTL___near_mem$imem_master_wready , RTL___near_mem$imem_master_wvalid , RTL___near_mem$imem_req_mstatus_MXR , RTL___near_mem$imem_req_sstatus_SUM , RTL___near_mem$imem_valid ; 
    wire[63:0] RTL___soc_map$m_is_IO_addr_addr , RTL___soc_map$m_is_mem_addr_addr , RTL___soc_map$m_is_near_mem_IO_addr_addr , RTL___soc_map$m_pc_reset_value ; 
    wire RTL___stage1_f_reset_reqs$CLR , RTL___stage1_f_reset_reqs$DEQ , RTL___stage1_f_reset_reqs$EMPTY_N , RTL___stage1_f_reset_reqs$ENQ , RTL___stage1_f_reset_reqs$FULL_N ; 
    wire RTL___stage1_f_reset_rsps$CLR , RTL___stage1_f_reset_rsps$DEQ , RTL___stage1_f_reset_rsps$EMPTY_N , RTL___stage1_f_reset_rsps$ENQ , RTL___stage1_f_reset_rsps$FULL_N ; 
    wire RTL___stage2_f_reset_reqs$CLR , RTL___stage2_f_reset_reqs$DEQ , RTL___stage2_f_reset_reqs$EMPTY_N , RTL___stage2_f_reset_reqs$ENQ , RTL___stage2_f_reset_reqs$FULL_N ; 
    wire RTL___stage2_f_reset_rsps$CLR , RTL___stage2_f_reset_rsps$DEQ , RTL___stage2_f_reset_rsps$EMPTY_N , RTL___stage2_f_reset_rsps$ENQ , RTL___stage2_f_reset_rsps$FULL_N ; 
    wire RTL___stage3_f_reset_reqs$CLR , RTL___stage3_f_reset_reqs$DEQ , RTL___stage3_f_reset_reqs$EMPTY_N , RTL___stage3_f_reset_reqs$ENQ , RTL___stage3_f_reset_reqs$FULL_N ; 
    wire RTL___stage3_f_reset_rsps$CLR , RTL___stage3_f_reset_rsps$DEQ , RTL___stage3_f_reset_rsps$EMPTY_N , RTL___stage3_f_reset_rsps$ENQ , RTL___stage3_f_reset_rsps$FULL_N ; 
    wire RTL___CAN_FIRE_RL_rl_WFI_resume , RTL___CAN_FIRE_RL_rl_finish_FENCE , RTL___CAN_FIRE_RL_rl_finish_FENCE_I , RTL___CAN_FIRE_RL_rl_finish_SFENCE_VMA , RTL___CAN_FIRE_RL_rl_pipe , RTL___CAN_FIRE_RL_rl_reset_complete , RTL___CAN_FIRE_RL_rl_reset_from_WFI , RTL___CAN_FIRE_RL_rl_reset_start , RTL___CAN_FIRE_RL_rl_show_pipe , RTL___CAN_FIRE_RL_rl_stage1_CSRR_S_or_C , RTL___CAN_FIRE_RL_rl_stage1_CSRR_S_or_C_2 , RTL___CAN_FIRE_RL_rl_stage1_CSRR_W , RTL___CAN_FIRE_RL_rl_stage1_CSRR_W_2 , RTL___CAN_FIRE_RL_rl_stage1_FENCE , RTL___CAN_FIRE_RL_rl_stage1_FENCE_I , RTL___CAN_FIRE_RL_rl_stage1_SFENCE_VMA , RTL___CAN_FIRE_RL_rl_stage1_WFI , RTL___CAN_FIRE_RL_rl_stage1_interrupt , RTL___CAN_FIRE_RL_rl_stage1_restart_after_csrrx , RTL___CAN_FIRE_RL_rl_stage1_trap , RTL___CAN_FIRE_RL_rl_stage1_xRET , RTL___CAN_FIRE_RL_rl_stage2_nonpipe , RTL___CAN_FIRE_RL_rl_trap , RTL___CAN_FIRE_RL_rl_trap_fetch , RTL___CAN_FIRE_RL_stage1_rl_reset , RTL___CAN_FIRE_RL_stage2_rl_reset_begin , RTL___CAN_FIRE_RL_stage2_rl_reset_end , RTL___CAN_FIRE_RL_stage3_rl_reset , RTL___CAN_FIRE_dmem_master_m_arready , RTL___CAN_FIRE_dmem_master_m_awready , RTL___CAN_FIRE_dmem_master_m_bvalid , RTL___CAN_FIRE_dmem_master_m_rvalid , RTL___CAN_FIRE_dmem_master_m_wready , RTL___CAN_FIRE_hart0_server_reset_request_put , RTL___CAN_FIRE_hart0_server_reset_response_get , RTL___CAN_FIRE_imem_master_m_arready , RTL___CAN_FIRE_imem_master_m_awready , RTL___CAN_FIRE_imem_master_m_bvalid , RTL___CAN_FIRE_imem_master_m_rvalid , RTL___CAN_FIRE_imem_master_m_wready , RTL___CAN_FIRE_m_external_interrupt_req , RTL___CAN_FIRE_nmi_req , RTL___CAN_FIRE_s_external_interrupt_req , RTL___CAN_FIRE_set_verbosity , RTL___CAN_FIRE_software_interrupt_req , RTL___CAN_FIRE_timer_interrupt_req , RTL___WILL_FIRE_RL_rl_WFI_resume , RTL___WILL_FIRE_RL_rl_finish_FENCE , RTL___WILL_FIRE_RL_rl_finish_FENCE_I , RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA , RTL___WILL_FIRE_RL_rl_pipe , RTL___WILL_FIRE_RL_rl_reset_complete , RTL___WILL_FIRE_RL_rl_reset_from_WFI , RTL___WILL_FIRE_RL_rl_reset_start , RTL___WILL_FIRE_RL_rl_show_pipe , RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C , RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 , RTL___WILL_FIRE_RL_rl_stage1_CSRR_W , RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 , RTL___WILL_FIRE_RL_rl_stage1_FENCE , RTL___WILL_FIRE_RL_rl_stage1_FENCE_I , RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA , RTL___WILL_FIRE_RL_rl_stage1_WFI , RTL___WILL_FIRE_RL_rl_stage1_interrupt , RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx , RTL___WILL_FIRE_RL_rl_stage1_trap , RTL___WILL_FIRE_RL_rl_stage1_xRET , RTL___WILL_FIRE_RL_rl_stage2_nonpipe , RTL___WILL_FIRE_RL_rl_trap , RTL___WILL_FIRE_RL_rl_trap_fetch , RTL___WILL_FIRE_RL_stage1_rl_reset , RTL___WILL_FIRE_RL_stage2_rl_reset_begin , RTL___WILL_FIRE_RL_stage2_rl_reset_end , RTL___WILL_FIRE_RL_stage3_rl_reset , RTL___WILL_FIRE_dmem_master_m_arready , RTL___WILL_FIRE_dmem_master_m_awready , RTL___WILL_FIRE_dmem_master_m_bvalid , RTL___WILL_FIRE_dmem_master_m_rvalid , RTL___WILL_FIRE_dmem_master_m_wready , RTL___WILL_FIRE_hart0_server_reset_request_put , RTL___WILL_FIRE_hart0_server_reset_response_get , RTL___WILL_FIRE_imem_master_m_arready , RTL___WILL_FIRE_imem_master_m_awready , RTL___WILL_FIRE_imem_master_m_bvalid , RTL___WILL_FIRE_imem_master_m_rvalid , RTL___WILL_FIRE_imem_master_m_wready , RTL___WILL_FIRE_m_external_interrupt_req , RTL___WILL_FIRE_nmi_req , RTL___WILL_FIRE_s_external_interrupt_req , RTL___WILL_FIRE_set_verbosity , RTL___WILL_FIRE_software_interrupt_req , RTL___WILL_FIRE_timer_interrupt_req ; reg[31:0] RTL___MUX_csr_regfile$mav_csr_write_2__VAL_2 ; 
    wire[67:0] RTL___MUX_rg_trap_info$write_1__VAL_1 , RTL___MUX_rg_trap_info$write_1__VAL_2 , RTL___MUX_rg_trap_info$write_1__VAL_3 , RTL___MUX_rg_trap_info$write_1__VAL_4 ; 
    wire[3:0] RTL___MUX_rg_state$write_1__VAL_1 , RTL___MUX_rg_state$write_1__VAL_2 , RTL___MUX_rg_state$write_1__VAL_3 ; 
    wire RTL___MUX_csr_regfile$mav_csr_write_1__SEL_1 , RTL___MUX_gpr_regfile$write_rd_1__SEL_3 , RTL___MUX_near_mem$imem_req_1__SEL_1 , RTL___MUX_near_mem$imem_req_1__SEL_2 , RTL___MUX_near_mem$imem_req_1__SEL_5 , RTL___MUX_rg_next_pc$write_1__SEL_1 , RTL___MUX_rg_retiring$write_1__SEL_1 , RTL___MUX_rg_state$write_1__SEL_1 , RTL___MUX_rg_state$write_1__SEL_10 , RTL___MUX_rg_state$write_1__SEL_4 , RTL___MUX_rg_state$write_1__SEL_6 , RTL___MUX_rg_state$write_1__SEL_7 , RTL___MUX_rg_state$write_1__SEL_8 , RTL___MUX_rg_state$write_1__SEL_9 , RTL___MUX_rg_trap_info$write_1__SEL_1 , RTL___MUX_rg_trap_instr$write_1__SEL_1 , RTL___MUX_rg_trap_interrupt$write_1__SEL_1 , RTL___MUX_s1_to_s2$write_1__VAL_1 , RTL___MUX_stage1_rg_full$write_1__VAL_10 , RTL___MUX_stage2_rg_full$write_1__VAL_3 ; reg[31:0] RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570 , RTL____theResult_____1_fst__h6569 , RTL___rs1_val__h11920 , RTL___x_out_data_to_stage2_addr__h5223 , RTL___x_out_data_to_stage2_val1__h5224 , RTL___x_out_data_to_stage3_rd_val__h4668 ; reg[4:0] RTL___x_out_data_to_stage3_rd__h4667 ; reg[3:0] RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10 , RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12 , RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11 , RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13 , RTL___CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4 , RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3 , RTL___IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413 , RTL___alu_outputs_exc_code__h5862 ; reg[1:0] RTL___CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5 , RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ; 
    reg RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8 , RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9 , RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 , RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ; 
    wire[127:0] RTL___csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 ; 
    wire[63:0] RTL____theResult____h10743 , RTL___cpi__h10745 , RTL___cpifrac__h10746 , RTL___delta_CPI_cycles__h10741 , RTL___delta_CPI_instrs___1__h10778 , RTL___delta_CPI_instrs__h10742 , RTL___x__h10744 ; 
    wire[35:0] RTL___IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 ; 
    wire[31:0] RTL___IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 , RTL___IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 , RTL___SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 , RTL____theResult_____1_fst__h6562 , RTL____theResult_____1_fst__h6597 , RTL____theResult___snd__h7382 , RTL___alu_outputs___1_addr__h5365 , RTL___alu_outputs___1_addr__h5385 , RTL___alu_outputs___1_addr__h5410 , RTL___alu_outputs___1_addr__h5583 , RTL___alu_outputs___1_val1__h5386 , RTL___alu_outputs___1_val1__h5480 , RTL___alu_outputs___1_val1__h5516 , RTL___alu_outputs___1_val1__h5847 , RTL___alu_outputs___1_val2__h5367 , RTL___data_to_stage2_addr__h5215 , RTL___eaddr__h5553 , RTL___fall_through_pc__h5175 , RTL___output_stage2___1_bypass_rd_val__h4960 , RTL___rd_val___1__h6550 , RTL___rd_val___1__h6558 , RTL___rd_val___1__h6565 , RTL___rd_val___1__h6572 , RTL___rd_val___1__h6579 , RTL___rd_val___1__h6586 , RTL___rd_val__h5072 , RTL___rd_val__h5132 , RTL___rd_val__h5523 , RTL___rd_val__h5537 , RTL___rd_val__h7278 , RTL___rd_val__h7330 , RTL___rd_val__h7352 , RTL___rs1_val__h11213 , RTL___rs1_val_bypassed__h3337 , RTL___rs2_val__h5339 , RTL___trap_info_tval__h6925 , RTL___val__h5074 , RTL___val__h5134 , RTL___value__h6967 , RTL___x_out_bypass_rd_val__h4969 , RTL___x_out_data_to_stage2_val2__h5225 , RTL___x_out_next_pc__h5189 , RTL___y__h12191 ; 
    wire[20:0] RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 ; 
    wire[12:0] RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 ; 
    wire[11:0] RTL___near_memimem_instr_BITS_31_TO_20__q7 , RTL___near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 ; 
    wire[4:0] RTL___shamt__h5467 , RTL___x_out_data_to_stage2_rd__h5222 ; 
    wire[3:0] RTL___IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 , RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 , RTL___IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 , RTL___alu_outputs___1_exc_code__h5362 , RTL___alu_outputs___1_exc_code__h5843 , RTL___cur_verbosity__h1827 , RTL___x_exc_code__h15410 , RTL___x_out_trap_info_exc_code__h6928 ; 
    wire[1:0] RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 , RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 , RTL___IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 , RTL___IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 ; 
    wire RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 , RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 , RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 , RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649 , RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 , RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 , RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 , RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 , RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 , RTL___NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 , RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 , RTL___NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 , RTL___NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 , RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 , RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 , RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 , RTL____0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 , RTL___csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 , RTL___gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 , RTL___gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 , RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 , RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 , RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 , RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 , RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 , RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 , RTL___rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392 , RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 , RTL___rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 ; 
  assign  RTL___RDY_hart0_server_reset_request_put = RTL___f_reset_reqs$FULL_N ; 
  assign  RTL___CAN_FIRE_hart0_server_reset_request_put = RTL___f_reset_reqs$FULL_N ; 
  assign  RTL___WILL_FIRE_hart0_server_reset_request_put = RTL___EN_hart0_server_reset_request_put ; 
  assign  RTL___hart0_server_reset_response_get = RTL___f_reset_rsps$D_OUT ; 
  assign  RTL___RDY_hart0_server_reset_response_get = RTL___f_reset_rsps$EMPTY_N ; 
  assign  RTL___CAN_FIRE_hart0_server_reset_response_get = RTL___f_reset_rsps$EMPTY_N ; 
  assign  RTL___WILL_FIRE_hart0_server_reset_response_get = RTL___EN_hart0_server_reset_response_get ; 
  assign  RTL___imem_master_awvalid = RTL___near_mem$imem_master_awvalid ; 
  assign  RTL___imem_master_awid = RTL___near_mem$imem_master_awid ; 
  assign  RTL___imem_master_awaddr = RTL___near_mem$imem_master_awaddr ; 
  assign  RTL___imem_master_awlen = RTL___near_mem$imem_master_awlen ; 
  assign  RTL___imem_master_awsize = RTL___near_mem$imem_master_awsize ; 
  assign  RTL___imem_master_awburst = RTL___near_mem$imem_master_awburst ; 
  assign  RTL___imem_master_awlock = RTL___near_mem$imem_master_awlock ; 
  assign  RTL___imem_master_awcache = RTL___near_mem$imem_master_awcache ; 
  assign  RTL___imem_master_awprot = RTL___near_mem$imem_master_awprot ; 
  assign  RTL___imem_master_awqos = RTL___near_mem$imem_master_awqos ; 
  assign  RTL___imem_master_awregion = RTL___near_mem$imem_master_awregion ; 
  assign  RTL___CAN_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL___WILL_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL___imem_master_wvalid = RTL___near_mem$imem_master_wvalid ; 
  assign  RTL___imem_master_wdata = RTL___near_mem$imem_master_wdata ; 
  assign  RTL___imem_master_wstrb = RTL___near_mem$imem_master_wstrb ; 
  assign  RTL___imem_master_wlast = RTL___near_mem$imem_master_wlast ; 
  assign  RTL___CAN_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL___WILL_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL___CAN_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL___WILL_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL___imem_master_bready = RTL___near_mem$imem_master_bready ; 
  assign  RTL___imem_master_arvalid = RTL___near_mem$imem_master_arvalid ; 
  assign  RTL___imem_master_arid = RTL___near_mem$imem_master_arid ; 
  assign  RTL___imem_master_araddr = RTL___near_mem$imem_master_araddr ; 
  assign  RTL___imem_master_arlen = RTL___near_mem$imem_master_arlen ; 
  assign  RTL___imem_master_arsize = RTL___near_mem$imem_master_arsize ; 
  assign  RTL___imem_master_arburst = RTL___near_mem$imem_master_arburst ; 
  assign  RTL___imem_master_arlock = RTL___near_mem$imem_master_arlock ; 
  assign  RTL___imem_master_arcache = RTL___near_mem$imem_master_arcache ; 
  assign  RTL___imem_master_arprot = RTL___near_mem$imem_master_arprot ; 
  assign  RTL___imem_master_arqos = RTL___near_mem$imem_master_arqos ; 
  assign  RTL___imem_master_arregion = RTL___near_mem$imem_master_arregion ; 
  assign  RTL___CAN_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL___WILL_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL___CAN_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL___WILL_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL___imem_master_rready = RTL___near_mem$imem_master_rready ; 
  assign  RTL___dmem_master_awvalid = RTL___near_mem$dmem_master_awvalid ; 
  assign  RTL___dmem_master_awid = RTL___near_mem$dmem_master_awid ; 
  assign  RTL___dmem_master_awaddr = RTL___near_mem$dmem_master_awaddr ; 
  assign  RTL___dmem_master_awlen = RTL___near_mem$dmem_master_awlen ; 
  assign  RTL___dmem_master_awsize = RTL___near_mem$dmem_master_awsize ; 
  assign  RTL___dmem_master_awburst = RTL___near_mem$dmem_master_awburst ; 
  assign  RTL___dmem_master_awlock = RTL___near_mem$dmem_master_awlock ; 
  assign  RTL___dmem_master_awcache = RTL___near_mem$dmem_master_awcache ; 
  assign  RTL___dmem_master_awprot = RTL___near_mem$dmem_master_awprot ; 
  assign  RTL___dmem_master_awqos = RTL___near_mem$dmem_master_awqos ; 
  assign  RTL___dmem_master_awregion = RTL___near_mem$dmem_master_awregion ; 
  assign  RTL___CAN_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL___WILL_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL___dmem_master_wvalid = RTL___near_mem$dmem_master_wvalid ; 
  assign  RTL___dmem_master_wdata = RTL___near_mem$dmem_master_wdata ; 
  assign  RTL___dmem_master_wstrb = RTL___near_mem$dmem_master_wstrb ; 
  assign  RTL___dmem_master_wlast = RTL___near_mem$dmem_master_wlast ; 
  assign  RTL___CAN_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL___WILL_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL___CAN_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL___WILL_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL___dmem_master_bready = RTL___near_mem$dmem_master_bready ; 
  assign  RTL___dmem_master_arvalid = RTL___near_mem$dmem_master_arvalid ; 
  assign  RTL___dmem_master_arid = RTL___near_mem$dmem_master_arid ; 
  assign  RTL___dmem_master_araddr = RTL___near_mem$dmem_master_araddr ; 
  assign  RTL___dmem_master_arlen = RTL___near_mem$dmem_master_arlen ; 
  assign  RTL___dmem_master_arsize = RTL___near_mem$dmem_master_arsize ; 
  assign  RTL___dmem_master_arburst = RTL___near_mem$dmem_master_arburst ; 
  assign  RTL___dmem_master_arlock = RTL___near_mem$dmem_master_arlock ; 
  assign  RTL___dmem_master_arcache = RTL___near_mem$dmem_master_arcache ; 
  assign  RTL___dmem_master_arprot = RTL___near_mem$dmem_master_arprot ; 
  assign  RTL___dmem_master_arqos = RTL___near_mem$dmem_master_arqos ; 
  assign  RTL___dmem_master_arregion = RTL___near_mem$dmem_master_arregion ; 
  assign  RTL___CAN_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL___WILL_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL___CAN_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL___WILL_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL___dmem_master_rready = RTL___near_mem$dmem_master_rready ; 
  assign  RTL___CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___CAN_FIRE_nmi_req =1'd1; 
  assign  RTL___WILL_FIRE_nmi_req =1'd1; 
  assign  RTL___RDY_set_verbosity =1'd1; 
  assign  RTL___CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL___WILL_FIRE_set_verbosity = RTL___EN_set_verbosity ;  
    wire RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_nmi;
    wire RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_state;
    wire RTL___csr_regfile___CLK;
    wire RTL___csr_regfile___RST_N;
    wire RTL___csr_regfile___EN_server_reset_request_put;
    wire RTL___csr_regfile___EN_server_reset_response_get;
    wire[11:0] RTL___csr_regfile___read_csr_csr_addr;
    wire[11:0] RTL___csr_regfile___read_csr_port2_csr_addr;
    wire[11:0] RTL___csr_regfile___mav_read_csr_csr_addr;
    wire RTL___csr_regfile___EN_mav_read_csr;
    wire[11:0] RTL___csr_regfile___mav_csr_write_csr_addr;
    wire[31:0] RTL___csr_regfile___mav_csr_write_word;
    wire RTL___csr_regfile___EN_mav_csr_write;
    wire[1:0] RTL___csr_regfile___csr_trap_actions_from_priv;
    wire[31:0] RTL___csr_regfile___csr_trap_actions_pc;
    wire RTL___csr_regfile___csr_trap_actions_nmi;
    wire RTL___csr_regfile___csr_trap_actions_interrupt;
    wire[3:0] RTL___csr_regfile___csr_trap_actions_exc_code;
    wire[31:0] RTL___csr_regfile___csr_trap_actions_xtval;
    wire RTL___csr_regfile___EN_csr_trap_actions;
    wire[1:0] RTL___csr_regfile___csr_ret_actions_from_priv;
    wire RTL___csr_regfile___EN_csr_ret_actions;
    wire RTL___csr_regfile___EN_csr_minstret_incr;
    wire[1:0] RTL___csr_regfile___access_permitted_1_priv;
    wire[11:0] RTL___csr_regfile___access_permitted_1_csr_addr;
    wire RTL___csr_regfile___access_permitted_1_read_not_write;
    wire[1:0] RTL___csr_regfile___access_permitted_2_priv;
    wire[11:0] RTL___csr_regfile___access_permitted_2_csr_addr;
    wire RTL___csr_regfile___access_permitted_2_read_not_write;
    wire[1:0] RTL___csr_regfile___csr_counter_read_fault_priv;
    wire[11:0] RTL___csr_regfile___csr_counter_read_fault_csr_addr;
    wire RTL___csr_regfile___m_external_interrupt_req_set_not_clear;
    wire RTL___csr_regfile___s_external_interrupt_req_set_not_clear;
    wire RTL___csr_regfile___timer_interrupt_req_set_not_clear;
    wire RTL___csr_regfile___software_interrupt_req_set_not_clear;
    wire[1:0] RTL___csr_regfile___interrupt_pending_cur_priv;
    wire RTL___csr_regfile___nmi_req_set_not_clear;
    wire RTL___csr_regfile___EN_debug;

    wire[97:0] RTL___csr_regfile___csr_trap_actions ; 
    wire[65:0] RTL___csr_regfile___csr_ret_actions ; 
    wire[63:0] RTL___csr_regfile___read_csr_mcycle , RTL___csr_regfile___read_csr_minstret , RTL___csr_regfile___read_csr_mtime ; 
    wire[32:0] RTL___csr_regfile___mav_read_csr , RTL___csr_regfile___read_csr , RTL___csr_regfile___read_csr_port2 ; 
    wire[31:0] RTL___csr_regfile___csr_mip_read , RTL___csr_regfile___mav_csr_write , RTL___csr_regfile___read_mstatus , RTL___csr_regfile___read_satp , RTL___csr_regfile___read_ustatus ; 
    wire[27:0] RTL___csr_regfile___read_misa ; 
    wire[4:0] RTL___csr_regfile___interrupt_pending ; 
    wire RTL___csr_regfile___RDY_csr_ret_actions , RTL___csr_regfile___RDY_csr_trap_actions , RTL___csr_regfile___RDY_debug , RTL___csr_regfile___RDY_server_reset_request_put , RTL___csr_regfile___RDY_server_reset_response_get , RTL___csr_regfile___access_permitted_1 , RTL___csr_regfile___access_permitted_2 , RTL___csr_regfile___csr_counter_read_fault , RTL___csr_regfile___nmi_pending , RTL___csr_regfile___wfi_resume ; reg[3:0] RTL___csr_regfile___cfg_verbosity ; 
    wire[3:0] RTL___csr_regfile___cfg_verbosity$D_IN ; 
    wire RTL___csr_regfile___cfg_verbosity$EN ; reg[31:0] RTL___csr_regfile___csr_mstatus_rg_mstatus ; reg[31:0] RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN ; 
    wire RTL___csr_regfile___csr_mstatus_rg_mstatus$EN ; reg[31:0] RTL___csr_regfile___rg_dcsr ; 
    wire[31:0] RTL___csr_regfile___rg_dcsr$D_IN ; 
    wire RTL___csr_regfile___rg_dcsr$EN ; reg[31:0] RTL___csr_regfile___rg_dpc ; 
    wire[31:0] RTL___csr_regfile___rg_dpc$D_IN ; 
    wire RTL___csr_regfile___rg_dpc$EN ; reg[31:0] RTL___csr_regfile___rg_dscratch0 ; 
    wire[31:0] RTL___csr_regfile___rg_dscratch0$D_IN ; 
    wire RTL___csr_regfile___rg_dscratch0$EN ; reg[31:0] RTL___csr_regfile___rg_dscratch1 ; 
    wire[31:0] RTL___csr_regfile___rg_dscratch1$D_IN ; 
    wire RTL___csr_regfile___rg_dscratch1$EN ; reg[4:0] RTL___csr_regfile___rg_mcause ; reg[4:0] RTL___csr_regfile___rg_mcause$D_IN ; 
    wire RTL___csr_regfile___rg_mcause$EN ; reg[2:0] RTL___csr_regfile___rg_mcounteren ; 
    wire[2:0] RTL___csr_regfile___rg_mcounteren$D_IN ; 
    wire RTL___csr_regfile___rg_mcounteren$EN ; reg[63:0] RTL___csr_regfile___rg_mcycle ; 
    wire[63:0] RTL___csr_regfile___rg_mcycle$D_IN ; 
    wire RTL___csr_regfile___rg_mcycle$EN ; reg[31:0] RTL___csr_regfile___rg_mepc ; 
    wire[31:0] RTL___csr_regfile___rg_mepc$D_IN ; 
    wire RTL___csr_regfile___rg_mepc$EN ; reg[63:0] RTL___csr_regfile___rg_minstret ; 
    wire[63:0] RTL___csr_regfile___rg_minstret$D_IN ; 
    wire RTL___csr_regfile___rg_minstret$EN ; reg[31:0] RTL___csr_regfile___rg_mscratch ; 
    wire[31:0] RTL___csr_regfile___rg_mscratch$D_IN ; 
    wire RTL___csr_regfile___rg_mscratch$EN ; reg[31:0] RTL___csr_regfile___rg_mtval ; 
    wire[31:0] RTL___csr_regfile___rg_mtval$D_IN ; 
    wire RTL___csr_regfile___rg_mtval$EN ; reg[30:0] RTL___csr_regfile___rg_mtvec ; 
    wire[30:0] RTL___csr_regfile___rg_mtvec$D_IN ; 
    wire RTL___csr_regfile___rg_mtvec$EN ; 
    reg RTL___csr_regfile___rg_nmi ; 
    wire RTL___csr_regfile___rg_nmi$D_IN , RTL___csr_regfile___rg_nmi$EN ; reg[31:0] RTL___csr_regfile___rg_nmi_vector ; 
    wire[31:0] RTL___csr_regfile___rg_nmi_vector$D_IN ; 
    wire RTL___csr_regfile___rg_nmi_vector$EN ; 
    reg RTL___csr_regfile___rg_state ; 
    wire RTL___csr_regfile___rg_state$D_IN , RTL___csr_regfile___rg_state$EN ; reg[31:0] RTL___csr_regfile___rg_tdata1 ; 
    wire[31:0] RTL___csr_regfile___rg_tdata1$D_IN ; 
    wire RTL___csr_regfile___rg_tdata1$EN ; reg[31:0] RTL___csr_regfile___rg_tdata2 ; 
    wire[31:0] RTL___csr_regfile___rg_tdata2$D_IN ; 
    wire RTL___csr_regfile___rg_tdata2$EN ; reg[31:0] RTL___csr_regfile___rg_tdata3 ; 
    wire[31:0] RTL___csr_regfile___rg_tdata3$D_IN ; 
    wire RTL___csr_regfile___rg_tdata3$EN ; reg[31:0] RTL___csr_regfile___rg_tselect ; 
    wire[31:0] RTL___csr_regfile___rg_tselect$D_IN ; 
    wire RTL___csr_regfile___rg_tselect$EN ; 
    wire[31:0] RTL___csr_regfile___csr_mie$fav_write , RTL___csr_regfile___csr_mie$fav_write_wordxl , RTL___csr_regfile___csr_mie$fv_read ; 
    wire[27:0] RTL___csr_regfile___csr_mie$fav_write_misa ; 
    wire RTL___csr_regfile___csr_mie$EN_fav_write , RTL___csr_regfile___csr_mie$EN_reset ; 
    wire[31:0] RTL___csr_regfile___csr_mip$fav_write , RTL___csr_regfile___csr_mip$fav_write_wordxl , RTL___csr_regfile___csr_mip$fv_read ; 
    wire[27:0] RTL___csr_regfile___csr_mip$fav_write_misa ; 
    wire RTL___csr_regfile___csr_mip$EN_fav_write , RTL___csr_regfile___csr_mip$EN_reset , RTL___csr_regfile___csr_mip$m_external_interrupt_req_req , RTL___csr_regfile___csr_mip$s_external_interrupt_req_req , RTL___csr_regfile___csr_mip$software_interrupt_req_req , RTL___csr_regfile___csr_mip$timer_interrupt_req_req ; 
    wire RTL___csr_regfile___f_reset_rsps$CLR , RTL___csr_regfile___f_reset_rsps$DEQ , RTL___csr_regfile___f_reset_rsps$EMPTY_N , RTL___csr_regfile___f_reset_rsps$ENQ , RTL___csr_regfile___f_reset_rsps$FULL_N ; 
    wire[63:0] RTL___csr_regfile___soc_map$m_is_IO_addr_addr , RTL___csr_regfile___soc_map$m_is_mem_addr_addr , RTL___csr_regfile___soc_map$m_is_near_mem_IO_addr_addr , RTL___csr_regfile___soc_map$m_mtvec_reset_value , RTL___csr_regfile___soc_map$m_nmivec_reset_value ; 
    wire RTL___csr_regfile___CAN_FIRE_RL_rl_mcycle_incr , RTL___csr_regfile___CAN_FIRE_RL_rl_reset_start , RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_csrrx , RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_incr , RTL___csr_regfile___CAN_FIRE_csr_minstret_incr , RTL___csr_regfile___CAN_FIRE_csr_ret_actions , RTL___csr_regfile___CAN_FIRE_csr_trap_actions , RTL___csr_regfile___CAN_FIRE_debug , RTL___csr_regfile___CAN_FIRE_m_external_interrupt_req , RTL___csr_regfile___CAN_FIRE_mav_csr_write , RTL___csr_regfile___CAN_FIRE_mav_read_csr , RTL___csr_regfile___CAN_FIRE_nmi_req , RTL___csr_regfile___CAN_FIRE_s_external_interrupt_req , RTL___csr_regfile___CAN_FIRE_server_reset_request_put , RTL___csr_regfile___CAN_FIRE_server_reset_response_get , RTL___csr_regfile___CAN_FIRE_software_interrupt_req , RTL___csr_regfile___CAN_FIRE_timer_interrupt_req , RTL___csr_regfile___WILL_FIRE_RL_rl_mcycle_incr , RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start , RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_csrrx , RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_incr , RTL___csr_regfile___WILL_FIRE_csr_minstret_incr , RTL___csr_regfile___WILL_FIRE_csr_ret_actions , RTL___csr_regfile___WILL_FIRE_csr_trap_actions , RTL___csr_regfile___WILL_FIRE_debug , RTL___csr_regfile___WILL_FIRE_m_external_interrupt_req , RTL___csr_regfile___WILL_FIRE_mav_csr_write , RTL___csr_regfile___WILL_FIRE_mav_read_csr , RTL___csr_regfile___WILL_FIRE_nmi_req , RTL___csr_regfile___WILL_FIRE_s_external_interrupt_req , RTL___csr_regfile___WILL_FIRE_server_reset_request_put , RTL___csr_regfile___WILL_FIRE_server_reset_response_get , RTL___csr_regfile___WILL_FIRE_software_interrupt_req , RTL___csr_regfile___WILL_FIRE_timer_interrupt_req ; 
    wire[63:0] RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_1 , RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_2 , RTL___csr_regfile___MUX_rw_minstret$wset_1__VAL_1 ; 
    wire[31:0] RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ; 
    wire[30:0] RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_1 , RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_2 ; 
    wire[4:0] RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_2 , RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_3 ; 
    wire RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__SEL_2 , RTL___csr_regfile___MUX_rg_mcause$write_1__SEL_2 , RTL___csr_regfile___MUX_rg_mcounteren$write_1__SEL_1 , RTL___csr_regfile___MUX_rg_mepc$write_1__SEL_1 , RTL___csr_regfile___MUX_rg_mtval$write_1__SEL_1 , RTL___csr_regfile___MUX_rg_mtvec$write_1__SEL_1 , RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 , RTL___csr_regfile___MUX_rg_tdata1$write_1__SEL_1 , RTL___csr_regfile___MUX_rw_minstret$wset_1__SEL_1 ; reg[31:0] RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769 , RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574 , RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220 , RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397 ; 
    wire[63:0] RTL___csr_regfile___x__h5174 , RTL___csr_regfile___x__h5282 ; 
    wire[33:0] RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 ; 
    wire[31:0] RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 , RTL___csr_regfile____theResult___fst__h8211 , RTL___csr_regfile____theResult___fst__h8412 , RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 , RTL___csr_regfile___exc_pc___1__h7296 , RTL___csr_regfile___exc_pc__h7032 , RTL___csr_regfile___exc_pc__h7243 , RTL___csr_regfile___mask__h8232 , RTL___csr_regfile___mask__h8249 , RTL___csr_regfile___result__h4701 , RTL___csr_regfile___result__h5357 , RTL___csr_regfile___v__h4509 , RTL___csr_regfile___v__h4571 , RTL___csr_regfile___v__h4742 , RTL___csr_regfile___val__h8250 , RTL___csr_regfile___vector_offset__h7244 , RTL___csr_regfile___wordxl1__h4038 , RTL___csr_regfile___x__h5843 , RTL___csr_regfile___x__h8067 , RTL___csr_regfile___x__h8068 , RTL___csr_regfile___x__h8085 , RTL___csr_regfile___x__h8231 , RTL___csr_regfile___x__h8244 , RTL___csr_regfile___x__h8261 , RTL___csr_regfile___y__h8245 , RTL___csr_regfile___y__h8262 ; 
    wire[22:0] RTL___csr_regfile___fixed_up_val_23__h4079 , RTL___csr_regfile___fixed_up_val_23__h6471 , RTL___csr_regfile___fixed_up_val_23__h8130 ; 
    wire[5:0] RTL___csr_regfile___ie_from_x__h8195 , RTL___csr_regfile___pie_from_x__h8196 ; 
    wire[3:0] RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 , RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 , RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 , RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 , RTL___csr_regfile___exc_code__h7909 ; 
    wire[1:0] RTL___csr_regfile___mpp__h7337 , RTL___csr_regfile___to_y__h8411 ; 
    wire RTL___csr_regfile___NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 , RTL___csr_regfile___NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 , RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364 , RTL___csr_regfile___NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 , RTL___csr_regfile___NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746 , RTL___csr_regfile___b__h8248 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 , RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 , RTL___csr_regfile___csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 , RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 , RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 , RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 , RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 ; 
  assign  RTL___csr_regfile___RDY_server_reset_request_put = RTL___csr_regfile___f_reset_rsps$FULL_N ; 
  assign  RTL___csr_regfile___CAN_FIRE_server_reset_request_put = RTL___csr_regfile___f_reset_rsps$FULL_N ; 
  assign  RTL___csr_regfile___WILL_FIRE_server_reset_request_put = RTL___csr_regfile___EN_server_reset_request_put ; 
  assign  RTL___csr_regfile___RDY_server_reset_response_get = RTL___csr_regfile___rg_state && RTL___csr_regfile___f_reset_rsps$EMPTY_N ; 
  assign  RTL___csr_regfile___CAN_FIRE_server_reset_response_get = RTL___csr_regfile___rg_state && RTL___csr_regfile___f_reset_rsps$EMPTY_N ; 
  assign  RTL___csr_regfile___WILL_FIRE_server_reset_response_get = RTL___csr_regfile___EN_server_reset_response_get ; 
  assign  RTL___csr_regfile___read_csr ={ RTL___csr_regfile___read_csr_csr_addr >=12'hC03&& RTL___csr_regfile___read_csr_csr_addr <=12'hC1F|| RTL___csr_regfile___read_csr_csr_addr >=12'hC83&& RTL___csr_regfile___read_csr_csr_addr <=12'hC9F|| RTL___csr_regfile___read_csr_csr_addr >=12'hB03&& RTL___csr_regfile___read_csr_csr_addr <=12'hB1F|| RTL___csr_regfile___read_csr_csr_addr >=12'hB83&& RTL___csr_regfile___read_csr_csr_addr <=12'hB9F|| RTL___csr_regfile___read_csr_csr_addr >=12'h323&& RTL___csr_regfile___read_csr_csr_addr <=12'h33F|| RTL___csr_regfile___read_csr_csr_addr ==12'hC00|| RTL___csr_regfile___read_csr_csr_addr ==12'hC02|| RTL___csr_regfile___read_csr_csr_addr ==12'hC80|| RTL___csr_regfile___read_csr_csr_addr ==12'hC82|| RTL___csr_regfile___read_csr_csr_addr ==12'hF11|| RTL___csr_regfile___read_csr_csr_addr ==12'hF12|| RTL___csr_regfile___read_csr_csr_addr ==12'hF13|| RTL___csr_regfile___read_csr_csr_addr ==12'hF14|| RTL___csr_regfile___read_csr_csr_addr ==12'h300|| RTL___csr_regfile___read_csr_csr_addr ==12'h301|| RTL___csr_regfile___read_csr_csr_addr ==12'h304|| RTL___csr_regfile___read_csr_csr_addr ==12'h305|| RTL___csr_regfile___read_csr_csr_addr ==12'h306|| RTL___csr_regfile___read_csr_csr_addr ==12'h340|| RTL___csr_regfile___read_csr_csr_addr ==12'h341|| RTL___csr_regfile___read_csr_csr_addr ==12'h342|| RTL___csr_regfile___read_csr_csr_addr ==12'h343|| RTL___csr_regfile___read_csr_csr_addr ==12'h344|| RTL___csr_regfile___read_csr_csr_addr ==12'hB00|| RTL___csr_regfile___read_csr_csr_addr ==12'hB02|| RTL___csr_regfile___read_csr_csr_addr ==12'hB80|| RTL___csr_regfile___read_csr_csr_addr ==12'hB82|| RTL___csr_regfile___read_csr_csr_addr ==12'h7A0|| RTL___csr_regfile___read_csr_csr_addr ==12'h7A1|| RTL___csr_regfile___read_csr_csr_addr ==12'h7A2|| RTL___csr_regfile___read_csr_csr_addr ==12'h7A3,( RTL___csr_regfile___read_csr_csr_addr >=12'hC03&& RTL___csr_regfile___read_csr_csr_addr <=12'hC1F|| RTL___csr_regfile___read_csr_csr_addr >=12'hC83&& RTL___csr_regfile___read_csr_csr_addr <=12'hC9F|| RTL___csr_regfile___read_csr_csr_addr >=12'hB03&& RTL___csr_regfile___read_csr_csr_addr <=12'hB1F|| RTL___csr_regfile___read_csr_csr_addr >=12'hB83&& RTL___csr_regfile___read_csr_csr_addr <=12'hB9F|| RTL___csr_regfile___read_csr_csr_addr >=12'h323&& RTL___csr_regfile___read_csr_csr_addr <=12'h33F) ? 32'd0: RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220 }; 
  assign  RTL___csr_regfile___read_csr_port2 ={ RTL___csr_regfile___read_csr_port2_csr_addr >=12'hC03&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hC1F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hC83&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hC9F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hB03&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hB1F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hB83&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hB9F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'h323&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'h33F|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hC00|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hC02|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hC80|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hC82|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hF11|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hF12|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hF13|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hF14|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h300|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h301|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h304|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h305|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h306|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h340|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h341|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h342|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h343|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h344|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hB00|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hB02|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hB80|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'hB82|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h7A0|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h7A1|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h7A2|| RTL___csr_regfile___read_csr_port2_csr_addr ==12'h7A3,( RTL___csr_regfile___read_csr_port2_csr_addr >=12'hC03&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hC1F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hC83&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hC9F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hB03&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hB1F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'hB83&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'hB9F|| RTL___csr_regfile___read_csr_port2_csr_addr >=12'h323&& RTL___csr_regfile___read_csr_port2_csr_addr <=12'h33F) ? 32'd0: RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397 }; 
  assign  RTL___csr_regfile___mav_read_csr ={ RTL___csr_regfile___mav_read_csr_csr_addr >=12'hC03&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hC1F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hC83&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hC9F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hB03&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hB1F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hB83&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hB9F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'h323&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'h33F|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hC00|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hC02|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hC80|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hC82|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hF11|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hF12|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hF13|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hF14|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h300|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h301|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h304|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h305|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h306|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h340|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h341|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h342|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h343|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h344|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hB00|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hB02|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hB80|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'hB82|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h7A0|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h7A1|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h7A2|| RTL___csr_regfile___mav_read_csr_csr_addr ==12'h7A3,( RTL___csr_regfile___mav_read_csr_csr_addr >=12'hC03&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hC1F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hC83&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hC9F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hB03&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hB1F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'hB83&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'hB9F|| RTL___csr_regfile___mav_read_csr_csr_addr >=12'h323&& RTL___csr_regfile___mav_read_csr_csr_addr <=12'h33F) ? 32'd0: RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574 }; 
  assign  RTL___csr_regfile___CAN_FIRE_mav_read_csr =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_mav_read_csr = RTL___csr_regfile___EN_mav_read_csr ; 
  assign  RTL___csr_regfile___mav_csr_write = RTL___csr_regfile___NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746  ? 32'd0: RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769 ; 
  assign  RTL___csr_regfile___CAN_FIRE_mav_csr_write =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_mav_csr_write = RTL___csr_regfile___EN_mav_csr_write ; 
  assign  RTL___csr_regfile___read_misa =28'd68157696; 
  assign  RTL___csr_regfile___read_mstatus = RTL___csr_regfile___csr_mstatus_rg_mstatus ; 
  assign  RTL___csr_regfile___read_ustatus ={27'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus [4],3'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus [0]}; 
  assign  RTL___csr_regfile___read_satp =32'hAAAAAAAA; 
  assign  RTL___csr_regfile___csr_trap_actions ={ RTL___csr_regfile___x__h5843 , RTL___csr_regfile___x__h8067 , RTL___csr_regfile___x__h8068 ,2'b11}; 
  assign  RTL___csr_regfile___RDY_csr_trap_actions =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_csr_trap_actions =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_csr_trap_actions = RTL___csr_regfile___EN_csr_trap_actions ; 
  assign  RTL___csr_regfile___csr_ret_actions ={ RTL___csr_regfile___x__h8085 , RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 }; 
  assign  RTL___csr_regfile___RDY_csr_ret_actions =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_csr_ret_actions =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_csr_ret_actions = RTL___csr_regfile___EN_csr_ret_actions ; 
  assign  RTL___csr_regfile___read_csr_minstret = RTL___csr_regfile___rg_minstret ; 
  assign  RTL___csr_regfile___CAN_FIRE_csr_minstret_incr =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_csr_minstret_incr = RTL___csr_regfile___EN_csr_minstret_incr ; 
  assign  RTL___csr_regfile___read_csr_mcycle = RTL___csr_regfile___rg_mcycle ; 
  assign  RTL___csr_regfile___read_csr_mtime = RTL___csr_regfile___rg_mcycle ; 
  assign  RTL___csr_regfile___access_permitted_1 = RTL___csr_regfile___NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 &&( RTL___csr_regfile___access_permitted_1_read_not_write || RTL___csr_regfile___access_permitted_1_csr_addr [11:10]!=2'b11); 
  assign  RTL___csr_regfile___access_permitted_2 = RTL___csr_regfile___NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 &&( RTL___csr_regfile___access_permitted_2_read_not_write || RTL___csr_regfile___access_permitted_2_csr_addr [11:10]!=2'b11); 
  assign  RTL___csr_regfile___csr_counter_read_fault =( RTL___csr_regfile___csr_counter_read_fault_priv ==2'b01|| RTL___csr_regfile___csr_counter_read_fault_priv ==2'b0)&&( RTL___csr_regfile___csr_counter_read_fault_csr_addr ==12'hC00&&! RTL___csr_regfile___rg_mcounteren [0]|| RTL___csr_regfile___csr_counter_read_fault_csr_addr ==12'hC01&&! RTL___csr_regfile___rg_mcounteren [1]|| RTL___csr_regfile___csr_counter_read_fault_csr_addr ==12'hC02&&! RTL___csr_regfile___rg_mcounteren [2]|| RTL___csr_regfile___csr_counter_read_fault_csr_addr >=12'hC03&& RTL___csr_regfile___csr_counter_read_fault_csr_addr <=12'hC1F|| RTL___csr_regfile___csr_counter_read_fault_csr_addr >=12'hC83&& RTL___csr_regfile___csr_counter_read_fault_csr_addr <=12'hC9F); 
  assign  RTL___csr_regfile___csr_mip_read = RTL___csr_regfile___csr_mip$fv_read ; 
  assign  RTL___csr_regfile___CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___interrupt_pending ={ RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 , RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364  ? 4'd4: RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 }; 
  assign  RTL___csr_regfile___wfi_resume =( RTL___csr_regfile___csr_mip$fv_read & RTL___csr_regfile___csr_mie$fv_read )!=32'd0; 
  assign  RTL___csr_regfile___CAN_FIRE_nmi_req =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_nmi_req =1'd1; 
  assign  RTL___csr_regfile___nmi_pending = RTL___csr_regfile___rg_nmi ; 
  assign  RTL___csr_regfile___RDY_debug =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_debug =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_debug = RTL___csr_regfile___EN_debug ;  
    wire RTL___csr_regfile___csr_mie___CLK;
    wire RTL___csr_regfile___csr_mie___RST_N;
    wire RTL___csr_regfile___csr_mie___EN_reset;
    wire[27:0] RTL___csr_regfile___csr_mie___fav_write_misa;
    wire[31:0] RTL___csr_regfile___csr_mie___fav_write_wordxl;
    wire RTL___csr_regfile___csr_mie___EN_fav_write;

    wire[31:0] RTL___csr_regfile___csr_mie___fav_write , RTL___csr_regfile___csr_mie___fv_read ; reg[11:0] RTL___csr_regfile___csr_mie___rg_mie ; 
    wire[11:0] RTL___csr_regfile___csr_mie___rg_mie$D_IN ; 
    wire RTL___csr_regfile___csr_mie___rg_mie$EN ; 
    wire RTL___csr_regfile___csr_mie___CAN_FIRE_fav_write , RTL___csr_regfile___csr_mie___CAN_FIRE_reset , RTL___csr_regfile___csr_mie___WILL_FIRE_fav_write , RTL___csr_regfile___csr_mie___WILL_FIRE_reset ; 
    wire[11:0] RTL___csr_regfile___csr_mie___mie__h88 ; 
    wire RTL___csr_regfile___csr_mie___seie__h119 , RTL___csr_regfile___csr_mie___ssie__h113 , RTL___csr_regfile___csr_mie___stie__h116 , RTL___csr_regfile___csr_mie___ueie__h118 , RTL___csr_regfile___csr_mie___usie__h112 , RTL___csr_regfile___csr_mie___utie__h115 ; 
  assign  RTL___csr_regfile___csr_mie___CAN_FIRE_reset =1'd1; 
  assign  RTL___csr_regfile___csr_mie___WILL_FIRE_reset = RTL___csr_regfile___csr_mie___EN_reset ; 
  assign  RTL___csr_regfile___csr_mie___fv_read ={20'd0, RTL___csr_regfile___csr_mie___rg_mie }; 
  assign  RTL___csr_regfile___csr_mie___fav_write ={20'd0, RTL___csr_regfile___csr_mie___mie__h88 }; 
  assign  RTL___csr_regfile___csr_mie___CAN_FIRE_fav_write =1'd1; 
  assign  RTL___csr_regfile___csr_mie___WILL_FIRE_fav_write = RTL___csr_regfile___csr_mie___EN_fav_write ; 
  assign  RTL___csr_regfile___csr_mie___rg_mie$D_IN = RTL___csr_regfile___csr_mie___EN_fav_write  ?  RTL___csr_regfile___csr_mie___mie__h88 :12'd0; 
  assign  RTL___csr_regfile___csr_mie___rg_mie$EN = RTL___csr_regfile___csr_mie___EN_fav_write || RTL___csr_regfile___csr_mie___EN_reset ; 
  assign  RTL___csr_regfile___csr_mie___mie__h88 ={ RTL___csr_regfile___csr_mie___fav_write_wordxl [11],1'b0, RTL___csr_regfile___csr_mie___seie__h119 , RTL___csr_regfile___csr_mie___ueie__h118 , RTL___csr_regfile___csr_mie___fav_write_wordxl [7],1'b0, RTL___csr_regfile___csr_mie___stie__h116 , RTL___csr_regfile___csr_mie___utie__h115 , RTL___csr_regfile___csr_mie___fav_write_wordxl [3],1'b0, RTL___csr_regfile___csr_mie___ssie__h113 , RTL___csr_regfile___csr_mie___usie__h112 }; 
  assign  RTL___csr_regfile___csr_mie___seie__h119 = RTL___csr_regfile___csr_mie___fav_write_misa [18]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [9]; 
  assign  RTL___csr_regfile___csr_mie___ssie__h113 = RTL___csr_regfile___csr_mie___fav_write_misa [18]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [1]; 
  assign  RTL___csr_regfile___csr_mie___stie__h116 = RTL___csr_regfile___csr_mie___fav_write_misa [18]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [5]; 
  assign  RTL___csr_regfile___csr_mie___ueie__h118 = RTL___csr_regfile___csr_mie___fav_write_misa [13]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [8]; 
  assign  RTL___csr_regfile___csr_mie___usie__h112 = RTL___csr_regfile___csr_mie___fav_write_misa [13]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [0]; 
  assign  RTL___csr_regfile___csr_mie___utie__h115 = RTL___csr_regfile___csr_mie___fav_write_misa [13]&& RTL___csr_regfile___csr_mie___fav_write_wordxl [4]; 
  always @( posedge  RTL___csr_regfile___csr_mie___CLK )
         begin 
             if ( RTL___csr_regfile___csr_mie___RST_N ==1'b0)
                 begin  
                     RTL___csr_regfile___csr_mie___rg_mie  <=12'd0;
                 end 
              else 
                 begin 
                     if ( RTL___csr_regfile___csr_mie___rg_mie$EN ) 
                         RTL___csr_regfile___csr_mie___rg_mie  <= RTL___csr_regfile___csr_mie___rg_mie$D_IN ;
                 end 
         end
 
    assign RTL___csr_regfile___csr_mie___CLK = RTL___csr_regfile___CLK;
    assign RTL___csr_regfile___csr_mie___RST_N = RTL___csr_regfile___RST_N;
    assign RTL___csr_regfile___csr_mie___EN_reset = RTL___csr_regfile___csr_mie$EN_reset;
    assign RTL___csr_regfile___csr_mie$fv_read = RTL___csr_regfile___csr_mie___fv_read;
    assign RTL___csr_regfile___csr_mie___fav_write_misa = RTL___csr_regfile___csr_mie$fav_write_misa;
    assign RTL___csr_regfile___csr_mie___fav_write_wordxl = RTL___csr_regfile___csr_mie$fav_write_wordxl;
    assign RTL___csr_regfile___csr_mie___EN_fav_write = RTL___csr_regfile___csr_mie$EN_fav_write;
    assign RTL___csr_regfile___csr_mie$fav_write = RTL___csr_regfile___csr_mie___fav_write;
      
    wire RTL___csr_regfile___csr_mip___CLK;
    wire RTL___csr_regfile___csr_mip___RST_N;
    wire RTL___csr_regfile___csr_mip___EN_reset;
    wire[27:0] RTL___csr_regfile___csr_mip___fav_write_misa;
    wire[31:0] RTL___csr_regfile___csr_mip___fav_write_wordxl;
    wire RTL___csr_regfile___csr_mip___EN_fav_write;
    wire RTL___csr_regfile___csr_mip___m_external_interrupt_req_req;
    wire RTL___csr_regfile___csr_mip___s_external_interrupt_req_req;
    wire RTL___csr_regfile___csr_mip___software_interrupt_req_req;
    wire RTL___csr_regfile___csr_mip___timer_interrupt_req_req;

    wire[31:0] RTL___csr_regfile___csr_mip___fav_write , RTL___csr_regfile___csr_mip___fv_read ; 
    reg RTL___csr_regfile___csr_mip___rg_meip ; 
    wire RTL___csr_regfile___csr_mip___rg_meip$D_IN , RTL___csr_regfile___csr_mip___rg_meip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_msip ; 
    wire RTL___csr_regfile___csr_mip___rg_msip$D_IN , RTL___csr_regfile___csr_mip___rg_msip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_mtip ; 
    wire RTL___csr_regfile___csr_mip___rg_mtip$D_IN , RTL___csr_regfile___csr_mip___rg_mtip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_seip ; 
    wire RTL___csr_regfile___csr_mip___rg_seip$D_IN , RTL___csr_regfile___csr_mip___rg_seip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_ssip ; 
    wire RTL___csr_regfile___csr_mip___rg_ssip$D_IN , RTL___csr_regfile___csr_mip___rg_ssip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_stip ; 
    wire RTL___csr_regfile___csr_mip___rg_stip$D_IN , RTL___csr_regfile___csr_mip___rg_stip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_ueip ; 
    wire RTL___csr_regfile___csr_mip___rg_ueip$D_IN , RTL___csr_regfile___csr_mip___rg_ueip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_usip ; 
    wire RTL___csr_regfile___csr_mip___rg_usip$D_IN , RTL___csr_regfile___csr_mip___rg_usip$EN ; 
    reg RTL___csr_regfile___csr_mip___rg_utip ; 
    wire RTL___csr_regfile___csr_mip___rg_utip$D_IN , RTL___csr_regfile___csr_mip___rg_utip$EN ; 
    wire RTL___csr_regfile___csr_mip___CAN_FIRE_fav_write , RTL___csr_regfile___csr_mip___CAN_FIRE_m_external_interrupt_req , RTL___csr_regfile___csr_mip___CAN_FIRE_reset , RTL___csr_regfile___csr_mip___CAN_FIRE_s_external_interrupt_req , RTL___csr_regfile___csr_mip___CAN_FIRE_software_interrupt_req , RTL___csr_regfile___csr_mip___CAN_FIRE_timer_interrupt_req , RTL___csr_regfile___csr_mip___WILL_FIRE_fav_write , RTL___csr_regfile___csr_mip___WILL_FIRE_m_external_interrupt_req , RTL___csr_regfile___csr_mip___WILL_FIRE_reset , RTL___csr_regfile___csr_mip___WILL_FIRE_s_external_interrupt_req , RTL___csr_regfile___csr_mip___WILL_FIRE_software_interrupt_req , RTL___csr_regfile___csr_mip___WILL_FIRE_timer_interrupt_req ; 
    wire[11:0] RTL___csr_regfile___csr_mip___new_mip__h524 , RTL___csr_regfile___csr_mip___new_mip__h942 ; 
    wire RTL___csr_regfile___csr_mip___seip__h558 , RTL___csr_regfile___csr_mip___ssip__h562 , RTL___csr_regfile___csr_mip___stip__h560 , RTL___csr_regfile___csr_mip___ueip__h559 , RTL___csr_regfile___csr_mip___usip__h563 , RTL___csr_regfile___csr_mip___utip__h561 ; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_reset =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_reset = RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___fv_read ={20'd0, RTL___csr_regfile___csr_mip___new_mip__h524 }; 
  assign  RTL___csr_regfile___csr_mip___fav_write ={20'd0, RTL___csr_regfile___csr_mip___new_mip__h942 }; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_fav_write =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_fav_write = RTL___csr_regfile___csr_mip___EN_fav_write ; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_m_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_s_external_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_software_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___CAN_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___WILL_FIRE_timer_interrupt_req =1'd1; 
  assign  RTL___csr_regfile___csr_mip___rg_meip$D_IN = RTL___csr_regfile___csr_mip___m_external_interrupt_req_req ; 
  assign  RTL___csr_regfile___csr_mip___rg_meip$EN =1'b1; 
  assign  RTL___csr_regfile___csr_mip___rg_msip$D_IN = RTL___csr_regfile___csr_mip___software_interrupt_req_req ; 
  assign  RTL___csr_regfile___csr_mip___rg_msip$EN =1'b1; 
  assign  RTL___csr_regfile___csr_mip___rg_mtip$D_IN = RTL___csr_regfile___csr_mip___timer_interrupt_req_req ; 
  assign  RTL___csr_regfile___csr_mip___rg_mtip$EN =1'b1; 
  assign  RTL___csr_regfile___csr_mip___rg_seip$D_IN = RTL___csr_regfile___csr_mip___s_external_interrupt_req_req ; 
  assign  RTL___csr_regfile___csr_mip___rg_seip$EN =1'b1; 
  assign  RTL___csr_regfile___csr_mip___rg_ssip$D_IN =! RTL___csr_regfile___csr_mip___EN_reset && RTL___csr_regfile___csr_mip___ssip__h562 ; 
  assign  RTL___csr_regfile___csr_mip___rg_ssip$EN = RTL___csr_regfile___csr_mip___EN_fav_write || RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___rg_stip$D_IN =! RTL___csr_regfile___csr_mip___EN_reset && RTL___csr_regfile___csr_mip___stip__h560 ; 
  assign  RTL___csr_regfile___csr_mip___rg_stip$EN = RTL___csr_regfile___csr_mip___EN_fav_write || RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___rg_ueip$D_IN =! RTL___csr_regfile___csr_mip___EN_reset && RTL___csr_regfile___csr_mip___ueip__h559 ; 
  assign  RTL___csr_regfile___csr_mip___rg_ueip$EN = RTL___csr_regfile___csr_mip___EN_fav_write || RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___rg_usip$D_IN =! RTL___csr_regfile___csr_mip___EN_reset && RTL___csr_regfile___csr_mip___usip__h563 ; 
  assign  RTL___csr_regfile___csr_mip___rg_usip$EN = RTL___csr_regfile___csr_mip___EN_fav_write || RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___rg_utip$D_IN =! RTL___csr_regfile___csr_mip___EN_reset && RTL___csr_regfile___csr_mip___utip__h561 ; 
  assign  RTL___csr_regfile___csr_mip___rg_utip$EN = RTL___csr_regfile___csr_mip___EN_fav_write || RTL___csr_regfile___csr_mip___EN_reset ; 
  assign  RTL___csr_regfile___csr_mip___new_mip__h524 ={ RTL___csr_regfile___csr_mip___rg_meip ,1'b0, RTL___csr_regfile___csr_mip___rg_seip , RTL___csr_regfile___csr_mip___rg_ueip , RTL___csr_regfile___csr_mip___rg_mtip ,1'b0, RTL___csr_regfile___csr_mip___rg_stip , RTL___csr_regfile___csr_mip___rg_utip , RTL___csr_regfile___csr_mip___rg_msip ,1'b0, RTL___csr_regfile___csr_mip___rg_ssip , RTL___csr_regfile___csr_mip___rg_usip }; 
  assign  RTL___csr_regfile___csr_mip___new_mip__h942 ={ RTL___csr_regfile___csr_mip___rg_meip ,1'b0, RTL___csr_regfile___csr_mip___seip__h558 , RTL___csr_regfile___csr_mip___ueip__h559 , RTL___csr_regfile___csr_mip___rg_mtip ,1'b0, RTL___csr_regfile___csr_mip___stip__h560 , RTL___csr_regfile___csr_mip___utip__h561 , RTL___csr_regfile___csr_mip___rg_msip ,1'b0, RTL___csr_regfile___csr_mip___ssip__h562 , RTL___csr_regfile___csr_mip___usip__h563 }; 
  assign  RTL___csr_regfile___csr_mip___seip__h558 = RTL___csr_regfile___csr_mip___fav_write_misa [18]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [9]; 
  assign  RTL___csr_regfile___csr_mip___ssip__h562 = RTL___csr_regfile___csr_mip___fav_write_misa [18]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [1]; 
  assign  RTL___csr_regfile___csr_mip___stip__h560 = RTL___csr_regfile___csr_mip___fav_write_misa [18]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [5]; 
  assign  RTL___csr_regfile___csr_mip___ueip__h559 = RTL___csr_regfile___csr_mip___fav_write_misa [13]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [8]; 
  assign  RTL___csr_regfile___csr_mip___usip__h563 = RTL___csr_regfile___csr_mip___fav_write_misa [13]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [0]; 
  assign  RTL___csr_regfile___csr_mip___utip__h561 = RTL___csr_regfile___csr_mip___fav_write_misa [13]&& RTL___csr_regfile___csr_mip___fav_write_wordxl [4]; 
  always @( posedge  RTL___csr_regfile___csr_mip___CLK )
         begin 
             if ( RTL___csr_regfile___csr_mip___RST_N ==1'b0)
                 begin  
                     RTL___csr_regfile___csr_mip___rg_meip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_msip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_mtip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_seip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_ssip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_stip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_ueip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_usip  <=1'd0; 
                     RTL___csr_regfile___csr_mip___rg_utip  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL___csr_regfile___csr_mip___rg_meip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_meip  <= RTL___csr_regfile___csr_mip___rg_meip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_msip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_msip  <= RTL___csr_regfile___csr_mip___rg_msip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_mtip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_mtip  <= RTL___csr_regfile___csr_mip___rg_mtip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_seip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_seip  <= RTL___csr_regfile___csr_mip___rg_seip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_ssip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_ssip  <= RTL___csr_regfile___csr_mip___rg_ssip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_stip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_stip  <= RTL___csr_regfile___csr_mip___rg_stip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_ueip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_ueip  <= RTL___csr_regfile___csr_mip___rg_ueip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_usip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_usip  <= RTL___csr_regfile___csr_mip___rg_usip$D_IN ;
                     if ( RTL___csr_regfile___csr_mip___rg_utip$EN ) 
                         RTL___csr_regfile___csr_mip___rg_utip  <= RTL___csr_regfile___csr_mip___rg_utip$D_IN ;
                 end 
         end
 
    assign RTL___csr_regfile___csr_mip___CLK = RTL___csr_regfile___CLK;
    assign RTL___csr_regfile___csr_mip___RST_N = RTL___csr_regfile___RST_N;
    assign RTL___csr_regfile___csr_mip___EN_reset = RTL___csr_regfile___csr_mip$EN_reset;
    assign RTL___csr_regfile___csr_mip$fv_read = RTL___csr_regfile___csr_mip___fv_read;
    assign RTL___csr_regfile___csr_mip___fav_write_misa = RTL___csr_regfile___csr_mip$fav_write_misa;
    assign RTL___csr_regfile___csr_mip___fav_write_wordxl = RTL___csr_regfile___csr_mip$fav_write_wordxl;
    assign RTL___csr_regfile___csr_mip___EN_fav_write = RTL___csr_regfile___csr_mip$EN_fav_write;
    assign RTL___csr_regfile___csr_mip$fav_write = RTL___csr_regfile___csr_mip___fav_write;
    assign RTL___csr_regfile___csr_mip___m_external_interrupt_req_req = RTL___csr_regfile___csr_mip$m_external_interrupt_req_req;
    assign RTL___csr_regfile___csr_mip___s_external_interrupt_req_req = RTL___csr_regfile___csr_mip$s_external_interrupt_req_req;
    assign RTL___csr_regfile___csr_mip___software_interrupt_req_req = RTL___csr_regfile___csr_mip$software_interrupt_req_req;
    assign RTL___csr_regfile___csr_mip___timer_interrupt_req_req = RTL___csr_regfile___csr_mip$timer_interrupt_req_req;
      
    wire RTL___csr_regfile___f_reset_rsps___RST;
    wire RTL___csr_regfile___f_reset_rsps___CLK;
    wire RTL___csr_regfile___f_reset_rsps___ENQ;
    wire RTL___csr_regfile___f_reset_rsps___CLR;
    wire RTL___csr_regfile___f_reset_rsps___DEQ;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___csr_regfile___f_reset_rsps___FULL_N;
    wire RTL___csr_regfile___f_reset_rsps___EMPTY_N;
    wire RTL___stage1_f_reset_reqs___RST;
    wire RTL___stage1_f_reset_reqs___CLK;
    wire RTL___stage1_f_reset_reqs___ENQ;
    wire RTL___stage1_f_reset_reqs___CLR;
    wire RTL___stage1_f_reset_reqs___DEQ;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_reqs___FULL_N;
    wire RTL___stage1_f_reset_reqs___EMPTY_N;
    wire RTL___stage1_f_reset_rsps___RST;
    wire RTL___stage1_f_reset_rsps___CLK;
    wire RTL___stage1_f_reset_rsps___ENQ;
    wire RTL___stage1_f_reset_rsps___CLR;
    wire RTL___stage1_f_reset_rsps___DEQ;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage1_f_reset_rsps___FULL_N;
    wire RTL___stage1_f_reset_rsps___EMPTY_N;
    wire RTL___stage2_f_reset_reqs___RST;
    wire RTL___stage2_f_reset_reqs___CLK;
    wire RTL___stage2_f_reset_reqs___ENQ;
    wire RTL___stage2_f_reset_reqs___CLR;
    wire RTL___stage2_f_reset_reqs___DEQ;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_reqs___FULL_N;
    wire RTL___stage2_f_reset_reqs___EMPTY_N;
    wire RTL___stage2_f_reset_rsps___RST;
    wire RTL___stage2_f_reset_rsps___CLK;
    wire RTL___stage2_f_reset_rsps___ENQ;
    wire RTL___stage2_f_reset_rsps___CLR;
    wire RTL___stage2_f_reset_rsps___DEQ;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage2_f_reset_rsps___FULL_N;
    wire RTL___stage2_f_reset_rsps___EMPTY_N;
    wire RTL___stage3_f_reset_reqs___RST;
    wire RTL___stage3_f_reset_reqs___CLK;
    wire RTL___stage3_f_reset_reqs___ENQ;
    wire RTL___stage3_f_reset_reqs___CLR;
    wire RTL___stage3_f_reset_reqs___DEQ;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_reqs___FULL_N;
    wire RTL___stage3_f_reset_reqs___EMPTY_N;
    wire RTL___stage3_f_reset_rsps___RST;
    wire RTL___stage3_f_reset_rsps___CLK;
    wire RTL___stage3_f_reset_rsps___ENQ;
    wire RTL___stage3_f_reset_rsps___CLR;
    wire RTL___stage3_f_reset_rsps___DEQ;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___stage3_f_reset_rsps___FULL_N;
    wire RTL___stage3_f_reset_rsps___EMPTY_N;

    reg RTL___csr_regfile___f_reset_rsps___empty_reg ; 
    reg RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___FULL_N = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___EMPTY_N = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___csr_regfile___f_reset_rsps___CLK )
         begin 
             if ( RTL___csr_regfile___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___csr_regfile___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___csr_regfile___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___csr_regfile___f_reset_rsps___CLR )
                         begin  
                             RTL___csr_regfile___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___csr_regfile___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___csr_regfile___f_reset_rsps___ENQ &&! RTL___csr_regfile___f_reset_rsps___DEQ )
                             begin  
                                 RTL___csr_regfile___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___csr_regfile___f_reset_rsps___full_reg  <=! RTL___csr_regfile___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___csr_regfile___f_reset_rsps___ENQ && RTL___csr_regfile___f_reset_rsps___DEQ )
                                 begin  
                                     RTL___csr_regfile___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___csr_regfile___f_reset_rsps___empty_reg  <=! RTL___csr_regfile___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___csr_regfile___f_reset_rsps___CLK )
         begin : RTL___csr_regfile___f_reset_rsps___error_checks 
           reg RTL___csr_regfile___f_reset_rsps___deqerror , RTL___csr_regfile___f_reset_rsps___enqerror ; 
             RTL___csr_regfile___f_reset_rsps___deqerror  =0; 
             RTL___csr_regfile___f_reset_rsps___enqerror  =0;
             if ( RTL___csr_regfile___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___csr_regfile___f_reset_rsps___empty_reg && RTL___csr_regfile___f_reset_rsps___DEQ )
                         begin  
                             RTL___csr_regfile___f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___csr_regfile___f_reset_rsps___full_reg && RTL___csr_regfile___f_reset_rsps___ENQ &&(! RTL___csr_regfile___f_reset_rsps___DEQ || RTL___csr_regfile___f_reset_rsps___guarded ))
                         begin  
                             RTL___csr_regfile___f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___csr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___empty_reg ;
      
    wire RTL___csr_regfile___soc_map___CLK;
    wire RTL___csr_regfile___soc_map___RST_N;
    wire[63:0] RTL___csr_regfile___soc_map___m_is_mem_addr_addr;
    wire[63:0] RTL___csr_regfile___soc_map___m_is_IO_addr_addr;
    wire[63:0] RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr_addr;
    wire RTL___soc_map___CLK;
    wire RTL___soc_map___RST_N;
    wire[63:0] RTL___soc_map___m_is_mem_addr_addr;
    wire[63:0] RTL___soc_map___m_is_IO_addr_addr;
    wire[63:0] RTL___soc_map___m_is_near_mem_IO_addr_addr;

    wire[63:0] RTL___csr_regfile___soc_map___m_boot_rom_addr_base , RTL___csr_regfile___soc_map___m_boot_rom_addr_lim , RTL___csr_regfile___soc_map___m_boot_rom_addr_size , RTL___csr_regfile___soc_map___m_mem0_controller_addr_base , RTL___csr_regfile___soc_map___m_mem0_controller_addr_lim , RTL___csr_regfile___soc_map___m_mem0_controller_addr_size , RTL___csr_regfile___soc_map___m_mtvec_reset_value , RTL___csr_regfile___soc_map___m_near_mem_io_addr_base , RTL___csr_regfile___soc_map___m_near_mem_io_addr_lim , RTL___csr_regfile___soc_map___m_near_mem_io_addr_size , RTL___csr_regfile___soc_map___m_nmivec_reset_value , RTL___csr_regfile___soc_map___m_pc_reset_value , RTL___csr_regfile___soc_map___m_plic_addr_base , RTL___csr_regfile___soc_map___m_plic_addr_lim , RTL___csr_regfile___soc_map___m_plic_addr_size , RTL___csr_regfile___soc_map___m_tcm_addr_base , RTL___csr_regfile___soc_map___m_tcm_addr_lim , RTL___csr_regfile___soc_map___m_tcm_addr_size , RTL___csr_regfile___soc_map___m_uart0_addr_base , RTL___csr_regfile___soc_map___m_uart0_addr_lim , RTL___csr_regfile___soc_map___m_uart0_addr_size ; 
    wire RTL___csr_regfile___soc_map___m_is_IO_addr , RTL___csr_regfile___soc_map___m_is_mem_addr , RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr ; 
  assign  RTL___csr_regfile___soc_map___m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL___csr_regfile___soc_map___m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL___csr_regfile___soc_map___m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL___csr_regfile___soc_map___m_plic_addr_base =64'h000000000C000000; 
  assign  RTL___csr_regfile___soc_map___m_plic_addr_size =64'h0000000000400000; 
  assign  RTL___csr_regfile___soc_map___m_plic_addr_lim =64'd205520896; 
  assign  RTL___csr_regfile___soc_map___m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL___csr_regfile___soc_map___m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL___csr_regfile___soc_map___m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL___csr_regfile___soc_map___m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL___csr_regfile___soc_map___m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL___csr_regfile___soc_map___m_boot_rom_addr_lim =64'd8192; 
  assign  RTL___csr_regfile___soc_map___m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL___csr_regfile___soc_map___m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL___csr_regfile___soc_map___m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL___csr_regfile___soc_map___m_tcm_addr_base =64'h0; 
  assign  RTL___csr_regfile___soc_map___m_tcm_addr_size =64'd0; 
  assign  RTL___csr_regfile___soc_map___m_tcm_addr_lim =64'd0; 
  assign  RTL___csr_regfile___soc_map___m_is_mem_addr = RTL___csr_regfile___soc_map___m_is_mem_addr_addr >=64'h0000000000001000&& RTL___csr_regfile___soc_map___m_is_mem_addr_addr <64'd8192|| RTL___csr_regfile___soc_map___m_is_mem_addr_addr >=64'h0000000080000000&& RTL___csr_regfile___soc_map___m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL___csr_regfile___soc_map___m_is_IO_addr = RTL___csr_regfile___soc_map___m_is_IO_addr_addr >=64'h0000000002000000&& RTL___csr_regfile___soc_map___m_is_IO_addr_addr <64'd33603584|| RTL___csr_regfile___soc_map___m_is_IO_addr_addr >=64'h000000000C000000&& RTL___csr_regfile___soc_map___m_is_IO_addr_addr <64'd205520896|| RTL___csr_regfile___soc_map___m_is_IO_addr_addr >=64'h00000000C0000000&& RTL___csr_regfile___soc_map___m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr = RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL___csr_regfile___soc_map___m_pc_reset_value =64'h0000000000001000; 
  assign  RTL___csr_regfile___soc_map___m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL___csr_regfile___soc_map___m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL___csr_regfile___CAN_FIRE_RL_rl_reset_start =! RTL___csr_regfile___rg_state ; 
  assign  RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start = RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___csr_regfile___CAN_FIRE_RL_rl_mcycle_incr =1'd1; 
  assign  RTL___csr_regfile___WILL_FIRE_RL_rl_mcycle_incr =1'd1; 
  assign  RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_csrrx = RTL___csr_regfile___MUX_rw_minstret$wset_1__SEL_1 || RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_csrrx = RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_csrrx ; 
  assign  RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_incr =! RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_csrrx && RTL___csr_regfile___EN_csr_minstret_incr ; 
  assign  RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_incr = RTL___csr_regfile___CAN_FIRE_RL_rl_upd_minstret_incr ; 
  assign  RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__SEL_2 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h300; 
  assign  RTL___csr_regfile___MUX_rg_mcause$write_1__SEL_2 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h342; 
  assign  RTL___csr_regfile___MUX_rg_mcounteren$write_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h306; 
  assign  RTL___csr_regfile___MUX_rg_mepc$write_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h341; 
  assign  RTL___csr_regfile___MUX_rg_mtval$write_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h343; 
  assign  RTL___csr_regfile___MUX_rg_mtvec$write_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h305; 
  assign  RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 = RTL___csr_regfile___CAN_FIRE_RL_rl_reset_start &&! RTL___csr_regfile___EN_mav_csr_write ; 
  assign  RTL___csr_regfile___MUX_rg_tdata1$write_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h7A1; 
  assign  RTL___csr_regfile___MUX_rw_minstret$wset_1__SEL_1 = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 &&( RTL___csr_regfile___mav_csr_write_csr_addr ==12'hB02|| RTL___csr_regfile___mav_csr_write_csr_addr ==12'hB82); 
  assign  RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ={9'd0, RTL___csr_regfile___fixed_up_val_23__h8130 }; 
  assign  RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_2 ={ RTL___csr_regfile___mav_csr_write_word [31], RTL___csr_regfile___mav_csr_write_word [3:0]}; 
  assign  RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_3 ={! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt , RTL___csr_regfile___exc_code__h7909 }; 
  assign  RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_1 = RTL___csr_regfile___MUX_rw_minstret$wset_1__SEL_1  ?  RTL___csr_regfile___MUX_rw_minstret$wset_1__VAL_1 :64'd0; 
  assign  RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_2 = RTL___csr_regfile___rg_minstret +64'd1; 
  assign  RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_1 ={ RTL___csr_regfile___mav_csr_write_word [31:2], RTL___csr_regfile___mav_csr_write_word [0]}; 
  assign  RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_2 ={ RTL___csr_regfile___soc_map$m_mtvec_reset_value [31:2], RTL___csr_regfile___soc_map$m_mtvec_reset_value [0]}; 
  assign  RTL___csr_regfile___MUX_rw_minstret$wset_1__VAL_1 =( RTL___csr_regfile___mav_csr_write_csr_addr ==12'hB02) ?  RTL___csr_regfile___x__h5174 : RTL___csr_regfile___x__h5282 ; 
  assign  RTL___csr_regfile___cfg_verbosity$D_IN =4'h0; 
  assign  RTL___csr_regfile___cfg_verbosity$EN =1'b0; 
  always @(        RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start                      or   RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__SEL_2               or   RTL___csr_regfile___wordxl1__h4038              or   RTL___csr_regfile___EN_csr_ret_actions             or   RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__VAL_3            or   RTL___csr_regfile___EN_csr_trap_actions           or   RTL___csr_regfile___x__h8067  )
         case (1'b1) 
          RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start  : 
              RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN  =32'd0; 
          RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__SEL_2  : 
              RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN  = RTL___csr_regfile___wordxl1__h4038 ; 
          RTL___csr_regfile___EN_csr_ret_actions  : 
              RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN  = RTL___csr_regfile___MUX_csr_mstatus_rg_mstatus$write_1__VAL_3 ; 
          RTL___csr_regfile___EN_csr_trap_actions  : 
              RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN  = RTL___csr_regfile___x__h8067 ;
          default : 
              RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN  =32'hAAAAAAAA;endcase
  assign  RTL___csr_regfile___csr_mstatus_rg_mstatus$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h300|| RTL___csr_regfile___EN_csr_trap_actions || RTL___csr_regfile___EN_csr_ret_actions || RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_dcsr$D_IN =32'h0; 
  assign  RTL___csr_regfile___rg_dcsr$EN =1'b0; 
  assign  RTL___csr_regfile___rg_dpc$D_IN =32'h0; 
  assign  RTL___csr_regfile___rg_dpc$EN =1'b0; 
  assign  RTL___csr_regfile___rg_dscratch0$D_IN =32'h0; 
  assign  RTL___csr_regfile___rg_dscratch0$EN =1'b0; 
  assign  RTL___csr_regfile___rg_dscratch1$D_IN =32'h0; 
  assign  RTL___csr_regfile___rg_dscratch1$EN =1'b0; 
  always @(      RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start                  or   RTL___csr_regfile___MUX_rg_mcause$write_1__SEL_2             or   RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_2            or   RTL___csr_regfile___EN_csr_trap_actions           or   RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_3  )
         case (1'b1) 
          RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start  : 
              RTL___csr_regfile___rg_mcause$D_IN  =5'd0; 
          RTL___csr_regfile___MUX_rg_mcause$write_1__SEL_2  : 
              RTL___csr_regfile___rg_mcause$D_IN  = RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_2 ; 
          RTL___csr_regfile___EN_csr_trap_actions  : 
              RTL___csr_regfile___rg_mcause$D_IN  = RTL___csr_regfile___MUX_rg_mcause$write_1__VAL_3 ;
          default : 
              RTL___csr_regfile___rg_mcause$D_IN  =5'b01010;endcase
  assign  RTL___csr_regfile___rg_mcause$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h342|| RTL___csr_regfile___EN_csr_trap_actions || RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_mcounteren$D_IN = RTL___csr_regfile___MUX_rg_mcounteren$write_1__SEL_1  ?  RTL___csr_regfile___mav_csr_write_word [2:0]:3'd0; 
  assign  RTL___csr_regfile___rg_mcounteren$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h306|| RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_mcycle$D_IN = RTL___csr_regfile___rg_mcycle +64'd1; 
  assign  RTL___csr_regfile___rg_mcycle$EN =1'd1; 
  assign  RTL___csr_regfile___rg_mepc$D_IN = RTL___csr_regfile___MUX_rg_mepc$write_1__SEL_1  ?  RTL___csr_regfile___result__h4701 : RTL___csr_regfile___csr_trap_actions_pc ; 
  assign  RTL___csr_regfile___rg_mepc$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h341|| RTL___csr_regfile___EN_csr_trap_actions ; 
  assign  RTL___csr_regfile___rg_minstret$D_IN = RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_csrrx  ?  RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_1 : RTL___csr_regfile___MUX_rg_minstret$write_1__VAL_2 ; 
  assign  RTL___csr_regfile___rg_minstret$EN = RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_csrrx || RTL___csr_regfile___WILL_FIRE_RL_rl_upd_minstret_incr ; 
  assign  RTL___csr_regfile___rg_mscratch$D_IN = RTL___csr_regfile___mav_csr_write_word ; 
  assign  RTL___csr_regfile___rg_mscratch$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h340; 
  assign  RTL___csr_regfile___rg_mtval$D_IN = RTL___csr_regfile___MUX_rg_mtval$write_1__SEL_1  ?  RTL___csr_regfile___mav_csr_write_word : RTL___csr_regfile___csr_trap_actions_xtval ; 
  assign  RTL___csr_regfile___rg_mtval$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h343|| RTL___csr_regfile___EN_csr_trap_actions ; 
  assign  RTL___csr_regfile___rg_mtvec$D_IN = RTL___csr_regfile___MUX_rg_mtvec$write_1__SEL_1  ?  RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_1 : RTL___csr_regfile___MUX_rg_mtvec$write_1__VAL_2 ; 
  assign  RTL___csr_regfile___rg_mtvec$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h305|| RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_nmi$D_IN =! RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start && RTL___csr_regfile___nmi_req_set_not_clear ; 
  assign  RTL___csr_regfile___rg_nmi$EN =1'b1; 
  assign  RTL___csr_regfile___rg_nmi_vector$D_IN = RTL___csr_regfile___soc_map$m_nmivec_reset_value [31:0]; 
  assign  RTL___csr_regfile___rg_nmi_vector$EN = RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___csr_regfile___rg_state$D_IN =! RTL___csr_regfile___EN_server_reset_request_put ; 
  assign  RTL___csr_regfile___rg_state$EN = RTL___csr_regfile___EN_server_reset_request_put || RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_tdata1$D_IN = RTL___csr_regfile___MUX_rg_tdata1$write_1__SEL_1  ?  RTL___csr_regfile___result__h5357 :32'd0; 
  assign  RTL___csr_regfile___rg_tdata1$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h7A1|| RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___rg_tdata2$D_IN = RTL___csr_regfile___mav_csr_write_word ; 
  assign  RTL___csr_regfile___rg_tdata2$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h7A2; 
  assign  RTL___csr_regfile___rg_tdata3$D_IN = RTL___csr_regfile___mav_csr_write_word ; 
  assign  RTL___csr_regfile___rg_tdata3$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h7A3; 
  assign  RTL___csr_regfile___rg_tselect$D_IN =32'd0; 
  assign  RTL___csr_regfile___rg_tselect$EN = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h7A0|| RTL___csr_regfile___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile___csr_mie$fav_write_misa =28'd68157696; 
  assign  RTL___csr_regfile___csr_mie$fav_write_wordxl = RTL___csr_regfile___mav_csr_write_word ; 
  assign  RTL___csr_regfile___csr_mie$EN_reset = RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___csr_regfile___csr_mie$EN_fav_write = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h304; 
  assign  RTL___csr_regfile___csr_mip$fav_write_misa =28'd68157696; 
  assign  RTL___csr_regfile___csr_mip$fav_write_wordxl = RTL___csr_regfile___mav_csr_write_word ; 
  assign  RTL___csr_regfile___csr_mip$m_external_interrupt_req_req = RTL___csr_regfile___m_external_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile___csr_mip$s_external_interrupt_req_req = RTL___csr_regfile___s_external_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile___csr_mip$software_interrupt_req_req = RTL___csr_regfile___software_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile___csr_mip$timer_interrupt_req_req = RTL___csr_regfile___timer_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile___csr_mip$EN_reset = RTL___csr_regfile___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___csr_regfile___csr_mip$EN_fav_write = RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 && RTL___csr_regfile___mav_csr_write_csr_addr ==12'h344; 
  assign  RTL___csr_regfile___f_reset_rsps$ENQ = RTL___csr_regfile___EN_server_reset_request_put ; 
  assign  RTL___csr_regfile___f_reset_rsps$DEQ = RTL___csr_regfile___EN_server_reset_response_get ; 
  assign  RTL___csr_regfile___f_reset_rsps$CLR =1'b0; 
  assign  RTL___csr_regfile___soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL___csr_regfile___soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL___csr_regfile___soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 =(! RTL___csr_regfile___csr_mip$fv_read [11]||! RTL___csr_regfile___csr_mie$fv_read [11]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]) ? 4'd3:4'd11; 
  assign  RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339  ? 4'd9:( RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334  ? 4'd7: RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1370 ); 
  assign  RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349  ? 4'd5:( RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344  ? 4'd1: RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1372 ); 
  assign  RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1376 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359  ? 4'd0:( RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354  ? 4'd8: RTL___csr_regfile___IF_NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_N_ETC___d1374 ); 
  assign  RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 =( RTL___csr_regfile___csr_ret_actions_from_priv ==2'b11) ?  RTL___csr_regfile____theResult___fst__h8211 : RTL___csr_regfile____theResult___fst__h8412 ; 
  assign  RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1068 =( RTL___csr_regfile___csr_ret_actions_from_priv ==2'b11) ? { RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [12:11], RTL___csr_regfile____theResult___fst__h8211 }:{ RTL___csr_regfile___to_y__h8411 , RTL___csr_regfile____theResult___fst__h8412 }; 
  assign  RTL___csr_regfile___NOT_access_permitted_1_csr_addr_ULT_0xC03_069__ETC___d1155 =( RTL___csr_regfile___access_permitted_1_csr_addr >=12'hC03&& RTL___csr_regfile___access_permitted_1_csr_addr <=12'hC1F|| RTL___csr_regfile___access_permitted_1_csr_addr >=12'hB03&& RTL___csr_regfile___access_permitted_1_csr_addr <=12'hB1F|| RTL___csr_regfile___access_permitted_1_csr_addr >=12'hC83&& RTL___csr_regfile___access_permitted_1_csr_addr <=12'hC9F|| RTL___csr_regfile___access_permitted_1_csr_addr >=12'hB83&& RTL___csr_regfile___access_permitted_1_csr_addr <=12'hB9F|| RTL___csr_regfile___access_permitted_1_csr_addr >=12'h323&& RTL___csr_regfile___access_permitted_1_csr_addr <=12'h33F|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hC00|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hC02|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hC80|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hC81|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hC82|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hF11|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hF12|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hF13|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hF14|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h300|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h301|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h304|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h305|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h306|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h340|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h341|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h342|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h343|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h344|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hB00|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hB02|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hB80|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'hB82|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h7A0|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h7A1|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h7A2|| RTL___csr_regfile___access_permitted_1_csr_addr ==12'h7A3)&& RTL___csr_regfile___access_permitted_1_priv >= RTL___csr_regfile___access_permitted_1_csr_addr [9:8]&&( RTL___csr_regfile___access_permitted_1_csr_addr !=12'h180||! RTL___csr_regfile___csr_mstatus_rg_mstatus [20]); 
  assign  RTL___csr_regfile___NOT_access_permitted_2_csr_addr_ULT_0xC03_160__ETC___d1245 =( RTL___csr_regfile___access_permitted_2_csr_addr >=12'hC03&& RTL___csr_regfile___access_permitted_2_csr_addr <=12'hC1F|| RTL___csr_regfile___access_permitted_2_csr_addr >=12'hB03&& RTL___csr_regfile___access_permitted_2_csr_addr <=12'hB1F|| RTL___csr_regfile___access_permitted_2_csr_addr >=12'hC83&& RTL___csr_regfile___access_permitted_2_csr_addr <=12'hC9F|| RTL___csr_regfile___access_permitted_2_csr_addr >=12'hB83&& RTL___csr_regfile___access_permitted_2_csr_addr <=12'hB9F|| RTL___csr_regfile___access_permitted_2_csr_addr >=12'h323&& RTL___csr_regfile___access_permitted_2_csr_addr <=12'h33F|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hC00|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hC02|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hC80|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hC81|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hC82|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hF11|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hF12|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hF13|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hF14|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h300|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h301|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h304|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h305|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h306|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h340|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h341|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h342|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h343|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h344|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hB00|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hB02|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hB80|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'hB82|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h7A0|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h7A1|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h7A2|| RTL___csr_regfile___access_permitted_2_csr_addr ==12'h7A3)&& RTL___csr_regfile___access_permitted_2_priv >= RTL___csr_regfile___access_permitted_2_csr_addr [9:8]&&( RTL___csr_regfile___access_permitted_2_csr_addr !=12'h180||! RTL___csr_regfile___csr_mstatus_rg_mstatus [20]); 
  assign  RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 = RTL___csr_regfile___cfg_verbosity >4'd1; 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 =(! RTL___csr_regfile___csr_mip$fv_read [11]||! RTL___csr_regfile___csr_mie$fv_read [11]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3])&&(! RTL___csr_regfile___csr_mip$fv_read [3]||! RTL___csr_regfile___csr_mie$fv_read [3]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1334 &&(! RTL___csr_regfile___csr_mip$fv_read [7]||! RTL___csr_regfile___csr_mie$fv_read [7]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1339 &&(! RTL___csr_regfile___csr_mip$fv_read [9]||! RTL___csr_regfile___csr_mie$fv_read [9]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1344 &&(! RTL___csr_regfile___csr_mip$fv_read [1]||! RTL___csr_regfile___csr_mie$fv_read [1]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1349 &&(! RTL___csr_regfile___csr_mip$fv_read [5]||! RTL___csr_regfile___csr_mie$fv_read [5]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1354 &&(! RTL___csr_regfile___csr_mip$fv_read [8]||! RTL___csr_regfile___csr_mie$fv_read [8]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1364 = RTL___csr_regfile___NOT_csr_mip_fv_read__94_BIT_11_277_324_OR_NOT__ETC___d1359 &&(! RTL___csr_regfile___csr_mip$fv_read [0]||! RTL___csr_regfile___csr_mie$fv_read [0]|| RTL___csr_regfile___interrupt_pending_cur_priv ==2'b11&&! RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 =! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 !=4'd0&& RTL___csr_regfile___exc_code__h7909 !=4'd1&& RTL___csr_regfile___exc_code__h7909 !=4'd2&& RTL___csr_regfile___exc_code__h7909 !=4'd3&& RTL___csr_regfile___exc_code__h7909 !=4'd4&& RTL___csr_regfile___exc_code__h7909 !=4'd5&& RTL___csr_regfile___exc_code__h7909 !=4'd6&& RTL___csr_regfile___exc_code__h7909 !=4'd7&& RTL___csr_regfile___exc_code__h7909 !=4'd8&& RTL___csr_regfile___exc_code__h7909 !=4'd9&& RTL___csr_regfile___exc_code__h7909 !=4'd10&& RTL___csr_regfile___exc_code__h7909 !=4'd11; 
  assign  RTL___csr_regfile___NOT_mav_csr_write_csr_addr_ULT_0xB03_77_35_AND_ETC___d746 =! RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 && RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 && RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 && RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 || RTL___csr_regfile___mav_csr_write_csr_addr ==12'hF11|| RTL___csr_regfile___mav_csr_write_csr_addr ==12'hF12|| RTL___csr_regfile___mav_csr_write_csr_addr ==12'hF13|| RTL___csr_regfile___mav_csr_write_csr_addr ==12'hF14; 
  assign  RTL___csr_regfile____theResult___fst__h8211 ={ RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [31:13],2'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [10:0]}; 
  assign  RTL___csr_regfile____theResult___fst__h8412 ={ RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [31:9],1'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [7:0]}; 
  assign  RTL___csr_regfile___b__h8248 = RTL___csr_regfile___csr_mstatus_rg_mstatus [{3'd1, RTL___csr_regfile___csr_ret_actions_from_priv }]; 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 = RTL___csr_regfile___csr_mip$fv_read [11]&& RTL___csr_regfile___csr_mie$fv_read [11]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3])|| RTL___csr_regfile___csr_mip$fv_read [3]&& RTL___csr_regfile___csr_mie$fv_read [3]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1288 || RTL___csr_regfile___csr_mip$fv_read [7]&& RTL___csr_regfile___csr_mie$fv_read [7]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1293 || RTL___csr_regfile___csr_mip$fv_read [9]&& RTL___csr_regfile___csr_mie$fv_read [9]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1298 || RTL___csr_regfile___csr_mip$fv_read [1]&& RTL___csr_regfile___csr_mie$fv_read [1]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1303 || RTL___csr_regfile___csr_mip$fv_read [5]&& RTL___csr_regfile___csr_mie$fv_read [5]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1308 || RTL___csr_regfile___csr_mip$fv_read [8]&& RTL___csr_regfile___csr_mie$fv_read [8]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1313 || RTL___csr_regfile___csr_mip$fv_read [0]&& RTL___csr_regfile___csr_mie$fv_read [0]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1323 = RTL___csr_regfile___csr_mip_fv_read__94_BIT_11_277_AND_csr_mie_fv__ETC___d1318 || RTL___csr_regfile___csr_mip$fv_read [4]&& RTL___csr_regfile___csr_mie$fv_read [4]&&( RTL___csr_regfile___interrupt_pending_cur_priv !=2'b11|| RTL___csr_regfile___csr_mstatus_rg_mstatus [3]); 
  assign  RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 = RTL___csr_regfile___x__h8244 | RTL___csr_regfile___mask__h8232 ; 
  assign  RTL___csr_regfile___csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 =( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 !=4'd0&& RTL___csr_regfile___exc_code__h7909 !=4'd1&& RTL___csr_regfile___exc_code__h7909 !=4'd2&& RTL___csr_regfile___exc_code__h7909 !=4'd3&& RTL___csr_regfile___exc_code__h7909 !=4'd4&& RTL___csr_regfile___exc_code__h7909 !=4'd5&& RTL___csr_regfile___exc_code__h7909 !=4'd6&& RTL___csr_regfile___exc_code__h7909 !=4'd7&& RTL___csr_regfile___exc_code__h7909 !=4'd8&& RTL___csr_regfile___exc_code__h7909 !=4'd9&& RTL___csr_regfile___exc_code__h7909 !=4'd11&& RTL___csr_regfile___exc_code__h7909 !=4'd12&& RTL___csr_regfile___exc_code__h7909 !=4'd13&& RTL___csr_regfile___exc_code__h7909 !=4'd15; 
  assign  RTL___csr_regfile___exc_code__h7909 = RTL___csr_regfile___csr_trap_actions_nmi  ? 4'd0: RTL___csr_regfile___csr_trap_actions_exc_code ; 
  assign  RTL___csr_regfile___exc_pc___1__h7296 = RTL___csr_regfile___exc_pc__h7243 + RTL___csr_regfile___vector_offset__h7244 ; 
  assign  RTL___csr_regfile___exc_pc__h7032 ={ RTL___csr_regfile___rg_mtvec [30:1],2'd0}; 
  assign  RTL___csr_regfile___exc_pc__h7243 = RTL___csr_regfile___csr_trap_actions_nmi  ?  RTL___csr_regfile___rg_nmi_vector : RTL___csr_regfile___exc_pc__h7032 ; 
  assign  RTL___csr_regfile___fixed_up_val_23__h4079 ={ RTL___csr_regfile___mav_csr_write_word [22:17],4'd0,( RTL___csr_regfile___mav_csr_write_word [12:11]==2'b11) ?  RTL___csr_regfile___mav_csr_write_word [12:11]:2'b0, RTL___csr_regfile___mav_csr_write_word [10:9],1'd0, RTL___csr_regfile___mav_csr_write_word [7:6],2'd0, RTL___csr_regfile___mav_csr_write_word [3:2],2'd0}; 
  assign  RTL___csr_regfile___fixed_up_val_23__h6471 ={ RTL___csr_regfile___csr_mstatus_rg_mstatus [22:17],4'd0, RTL___csr_regfile___mpp__h7337 , RTL___csr_regfile___csr_mstatus_rg_mstatus [10:9],1'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus [3], RTL___csr_regfile___csr_mstatus_rg_mstatus [6],3'd0, RTL___csr_regfile___csr_mstatus_rg_mstatus [2],2'd0}; 
  assign  RTL___csr_regfile___fixed_up_val_23__h8130 ={ RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [22:17],4'd0,( RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [12:11]==2'b11) ?  RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [12:11]:2'b0, RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [10:9],1'd0, RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [7:6],2'd0, RTL___csr_regfile___IF_csr_ret_actions_from_priv_EQ_0b11_029_THEN__ETC___d1050 [3:2],2'd0}; 
  assign  RTL___csr_regfile___ie_from_x__h8195 ={4'd0, RTL___csr_regfile___csr_ret_actions_from_priv }; 
  assign  RTL___csr_regfile___mask__h8232 =32'd1<< RTL___csr_regfile___pie_from_x__h8196 ; 
  assign  RTL___csr_regfile___mask__h8249 =32'd1<< RTL___csr_regfile___ie_from_x__h8195 ; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 = RTL___csr_regfile___mav_csr_write_csr_addr <=12'h33F; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 = RTL___csr_regfile___mav_csr_write_csr_addr <=12'hB1F; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 = RTL___csr_regfile___mav_csr_write_csr_addr <=12'hB9F; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 =( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 )&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF11&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF12&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF13&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF14&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h300&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h301&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h304&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h305&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h306&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h340&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h341&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h342&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h343&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h344&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hB00&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hB02&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hB80&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hB82&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h7A0&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h7A1&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h7A2&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'h7A3; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 = RTL___csr_regfile___mav_csr_write_csr_addr <12'h323; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d590 =( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 )&&( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 ); 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d642 =( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 )&&( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323___d585 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0x33F___d586 )&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF11&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF12&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF13&& RTL___csr_regfile___mav_csr_write_csr_addr !=12'hF14; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 =( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB1F___d578 )&&( RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 ||! RTL___csr_regfile___mav_csr_write_csr_addr_ULE_0xB9F___d582 )&& RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0x323_85_OR_NOT_mav_ETC___d728 ; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03___d577 = RTL___csr_regfile___mav_csr_write_csr_addr <12'hB03; 
  assign  RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB83___d581 = RTL___csr_regfile___mav_csr_write_csr_addr <12'hB83; 
  assign  RTL___csr_regfile___mpp__h7337 =( RTL___csr_regfile___csr_trap_actions_from_priv ==2'b11) ?  RTL___csr_regfile___csr_trap_actions_from_priv :2'b0; 
  assign  RTL___csr_regfile___pie_from_x__h8196 ={4'd1, RTL___csr_regfile___csr_ret_actions_from_priv }; 
  assign  RTL___csr_regfile___result__h4701 ={ RTL___csr_regfile___mav_csr_write_word [31:2],2'd0}; 
  assign  RTL___csr_regfile___result__h5357 ={4'd0, RTL___csr_regfile___mav_csr_write_word [27:0]}; 
  assign  RTL___csr_regfile___to_y__h8411 ={1'b0, RTL___csr_regfile___csr_mstatus_rg_mstatus_76_AND_INV_1_SL_0_CONCA_ETC___d1043 [8]}; 
  assign  RTL___csr_regfile___v__h4509 ={ RTL___csr_regfile___mav_csr_write_word [31:2],1'b0, RTL___csr_regfile___mav_csr_write_word [0]}; 
  assign  RTL___csr_regfile___v__h4571 ={29'd0, RTL___csr_regfile___mav_csr_write_word [2:0]}; 
  assign  RTL___csr_regfile___v__h4742 ={ RTL___csr_regfile___mav_csr_write_word [31],27'd0, RTL___csr_regfile___mav_csr_write_word [3:0]}; 
  assign  RTL___csr_regfile___val__h8250 ={31'd0, RTL___csr_regfile___b__h8248 }<< RTL___csr_regfile___ie_from_x__h8195 ; 
  assign  RTL___csr_regfile___vector_offset__h7244 ={26'd0, RTL___csr_regfile___csr_trap_actions_exc_code ,2'd0}; 
  assign  RTL___csr_regfile___wordxl1__h4038 ={9'd0, RTL___csr_regfile___fixed_up_val_23__h4079 }; 
  assign  RTL___csr_regfile___x__h5174 ={ RTL___csr_regfile___rg_minstret [63:32], RTL___csr_regfile___mav_csr_write_word }; 
  assign  RTL___csr_regfile___x__h5282 ={ RTL___csr_regfile___mav_csr_write_word , RTL___csr_regfile___rg_minstret [31:0]}; 
  assign  RTL___csr_regfile___x__h5843 =( RTL___csr_regfile___csr_trap_actions_interrupt &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___rg_mtvec [0]) ?  RTL___csr_regfile___exc_pc___1__h7296 : RTL___csr_regfile___exc_pc__h7243 ; 
  assign  RTL___csr_regfile___x__h8067 ={9'd0, RTL___csr_regfile___fixed_up_val_23__h6471 }; 
  assign  RTL___csr_regfile___x__h8068 ={! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt ,27'd0, RTL___csr_regfile___exc_code__h7909 }; 
  assign  RTL___csr_regfile___x__h8085 ={ RTL___csr_regfile___rg_mepc [31:2],1'd0, RTL___csr_regfile___rg_mepc [0]}; 
  assign  RTL___csr_regfile___x__h8231 = RTL___csr_regfile___x__h8261 | RTL___csr_regfile___val__h8250 ; 
  assign  RTL___csr_regfile___x__h8244 = RTL___csr_regfile___x__h8231 & RTL___csr_regfile___y__h8245 ; 
  assign  RTL___csr_regfile___x__h8261 = RTL___csr_regfile___csr_mstatus_rg_mstatus & RTL___csr_regfile___y__h8262 ; 
  assign  RTL___csr_regfile___y__h8245 =~ RTL___csr_regfile___mask__h8232 ; 
  assign  RTL___csr_regfile___y__h8262 =~ RTL___csr_regfile___mask__h8249 ; 
  always @(                 RTL___csr_regfile___read_csr_csr_addr                                        or   RTL___csr_regfile___rg_tdata3                        or   RTL___csr_regfile___csr_mstatus_rg_mstatus                       or   RTL___csr_regfile___csr_mie$fv_read                      or   RTL___csr_regfile___rg_mtvec                     or   RTL___csr_regfile___rg_mcounteren                    or   RTL___csr_regfile___rg_mscratch                   or   RTL___csr_regfile___x__h8085                  or   RTL___csr_regfile___rg_mcause                 or   RTL___csr_regfile___rg_mtval                or   RTL___csr_regfile___csr_mip$fv_read               or   RTL___csr_regfile___rg_tselect              or   RTL___csr_regfile___rg_tdata1             or   RTL___csr_regfile___rg_tdata2            or   RTL___csr_regfile___rg_mcycle           or   RTL___csr_regfile___rg_minstret  )
         begin 
             case ( RTL___csr_regfile___read_csr_csr_addr )
              12 'h300: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  =32'd1074790656;
              12 'h304: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___csr_mie$fv_read ;
              12 'h305: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={ RTL___csr_regfile___rg_mtvec [30:1],1'b0, RTL___csr_regfile___rg_mtvec [0]};
              12 'h306: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={29'd0, RTL___csr_regfile___rg_mcounteren };
              12 'h340: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_mscratch ;
              12 'h341: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___x__h8085 ;
              12 'h342: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  ={ RTL___csr_regfile___rg_mcause [4],27'd0, RTL___csr_regfile___rg_mcause [3:0]};
              12 'h343: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_mtval ;
              12 'h344: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___csr_mip$fv_read ;
              12 'h7A0: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_tselect ;
              12 'h7A1: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_tdata1 ;
              12 'h7A2: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  =32'd0;
              default : 
                  RTL___csr_regfile___IF_read_csr_csr_addr_EQ_0xC00_9_THEN_rg_mcycle_ETC___d220  = RTL___csr_regfile___rg_tdata3 ;endcase
         end
  always @(                 RTL___csr_regfile___read_csr_port2_csr_addr                                        or   RTL___csr_regfile___rg_tdata3                        or   RTL___csr_regfile___csr_mstatus_rg_mstatus                       or   RTL___csr_regfile___csr_mie$fv_read                      or   RTL___csr_regfile___rg_mtvec                     or   RTL___csr_regfile___rg_mcounteren                    or   RTL___csr_regfile___rg_mscratch                   or   RTL___csr_regfile___x__h8085                  or   RTL___csr_regfile___rg_mcause                 or   RTL___csr_regfile___rg_mtval                or   RTL___csr_regfile___csr_mip$fv_read               or   RTL___csr_regfile___rg_tselect              or   RTL___csr_regfile___rg_tdata1             or   RTL___csr_regfile___rg_tdata2            or   RTL___csr_regfile___rg_mcycle           or   RTL___csr_regfile___rg_minstret  )
         begin 
             case ( RTL___csr_regfile___read_csr_port2_csr_addr )
              12 'h300: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  =32'd1074790656;
              12 'h304: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___csr_mie$fv_read ;
              12 'h305: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={ RTL___csr_regfile___rg_mtvec [30:1],1'b0, RTL___csr_regfile___rg_mtvec [0]};
              12 'h306: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={29'd0, RTL___csr_regfile___rg_mcounteren };
              12 'h340: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_mscratch ;
              12 'h341: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___x__h8085 ;
              12 'h342: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  ={ RTL___csr_regfile___rg_mcause [4],27'd0, RTL___csr_regfile___rg_mcause [3:0]};
              12 'h343: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_mtval ;
              12 'h344: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___csr_mip$fv_read ;
              12 'h7A0: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_tselect ;
              12 'h7A1: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_tdata1 ;
              12 'h7A2: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  =32'd0;
              default : 
                  RTL___csr_regfile___IF_read_csr_port2_csr_addr_EQ_0xC00_43_THEN_rg_ETC___d397  = RTL___csr_regfile___rg_tdata3 ;endcase
         end
  always @(                 RTL___csr_regfile___mav_read_csr_csr_addr                                        or   RTL___csr_regfile___rg_tdata3                        or   RTL___csr_regfile___csr_mstatus_rg_mstatus                       or   RTL___csr_regfile___csr_mie$fv_read                      or   RTL___csr_regfile___rg_mtvec                     or   RTL___csr_regfile___rg_mcounteren                    or   RTL___csr_regfile___rg_mscratch                   or   RTL___csr_regfile___x__h8085                  or   RTL___csr_regfile___rg_mcause                 or   RTL___csr_regfile___rg_mtval                or   RTL___csr_regfile___csr_mip$fv_read               or   RTL___csr_regfile___rg_tselect              or   RTL___csr_regfile___rg_tdata1             or   RTL___csr_regfile___rg_tdata2            or   RTL___csr_regfile___rg_mcycle           or   RTL___csr_regfile___rg_minstret  )
         begin 
             case ( RTL___csr_regfile___mav_read_csr_csr_addr )
              12 'h300: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___csr_mstatus_rg_mstatus ;
              12 'h301: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  =32'd1074790656;
              12 'h304: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___csr_mie$fv_read ;
              12 'h305: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={ RTL___csr_regfile___rg_mtvec [30:1],1'b0, RTL___csr_regfile___rg_mtvec [0]};
              12 'h306: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={29'd0, RTL___csr_regfile___rg_mcounteren };
              12 'h340: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_mscratch ;
              12 'h341: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___x__h8085 ;
              12 'h342: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  ={ RTL___csr_regfile___rg_mcause [4],27'd0, RTL___csr_regfile___rg_mcause [3:0]};
              12 'h343: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_mtval ;
              12 'h344: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___csr_mip$fv_read ;
              12 'h7A0: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_tselect ;
              12 'h7A1: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_tdata1 ;
              12 'h7A2: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_tdata2 ;
              12 'hB00,12'hC00: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_mcycle [31:0];
              12 'hB02,12'hC02: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_minstret [31:0];
              12 'hB80,12'hC80: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_mcycle [63:32];
              12 'hB82,12'hC82: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_minstret [63:32];
              12 'hF11,12'hF12,12'hF13,12'hF14: 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  =32'd0;
              default : 
                  RTL___csr_regfile___IF_mav_read_csr_csr_addr_EQ_0xC00_20_THEN_rg_m_ETC___d574  = RTL___csr_regfile___rg_tdata3 ;endcase
         end
  always @(           RTL___csr_regfile___mav_csr_write_csr_addr                            or   RTL___csr_regfile___mav_csr_write_word                  or   RTL___csr_regfile___wordxl1__h4038                 or   RTL___csr_regfile___csr_mie$fav_write                or   RTL___csr_regfile___v__h4509               or   RTL___csr_regfile___v__h4571              or   RTL___csr_regfile___result__h4701             or   RTL___csr_regfile___v__h4742            or   RTL___csr_regfile___csr_mip$fav_write           or   RTL___csr_regfile___result__h5357  )
         begin 
             case ( RTL___csr_regfile___mav_csr_write_csr_addr )
              12 'h300: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___wordxl1__h4038 ;
              12 'h301: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  =32'd1074790656;
              12 'h304: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___csr_mie$fav_write ;
              12 'h305: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___v__h4509 ;
              12 'h306: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___v__h4571 ;
              12 'h340,12'h343,12'hB00,12'hB02,12'hB80,12'hB82: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___mav_csr_write_word ;
              12 'h341: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___result__h4701 ;
              12 'h342: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___v__h4742 ;
              12 'h344: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___csr_mip$fav_write ;
              12 'h7A0: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  =32'd0;
              12 'h7A1: 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___result__h5357 ;
              default : 
                  RTL___csr_regfile___IF_mav_csr_write_csr_addr_EQ_0x300_91_THEN_0_C_ETC___d769  = RTL___csr_regfile___mav_csr_write_word ;endcase
         end
  always @( posedge  RTL___csr_regfile___CLK )
         begin 
             if ( RTL___csr_regfile___RST_N ==1'b0)
                 begin  
                     RTL___csr_regfile___cfg_verbosity  <=4'd0; 
                     RTL___csr_regfile___csr_mstatus_rg_mstatus  <=32'd0; 
                     RTL___csr_regfile___rg_mcycle  <=64'd0; 
                     RTL___csr_regfile___rg_minstret  <=64'd0; 
                     RTL___csr_regfile___rg_nmi  <=1'd0; 
                     RTL___csr_regfile___rg_state  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL___csr_regfile___cfg_verbosity$EN ) 
                         RTL___csr_regfile___cfg_verbosity  <= RTL___csr_regfile___cfg_verbosity$D_IN ;
                     if ( RTL___csr_regfile___csr_mstatus_rg_mstatus$EN ) 
                         RTL___csr_regfile___csr_mstatus_rg_mstatus  <= RTL___csr_regfile___csr_mstatus_rg_mstatus$D_IN ;
                     if ( RTL___csr_regfile___rg_mcycle$EN ) 
                         RTL___csr_regfile___rg_mcycle  <= RTL___csr_regfile___rg_mcycle$D_IN ;
                     if ( RTL___csr_regfile___rg_minstret$EN ) 
                         RTL___csr_regfile___rg_minstret  <= RTL___csr_regfile___rg_minstret$D_IN ;
                     if ( RTL___csr_regfile___rg_nmi$EN ) 
                         RTL___csr_regfile___rg_nmi  <= RTL___csr_regfile___rg_nmi$D_IN ;
                     if ( RTL___csr_regfile___rg_state$EN ) 
                         RTL___csr_regfile___rg_state  <= RTL___csr_regfile___rg_state$D_IN ;
                 end 
             if ( RTL___csr_regfile___rg_dcsr$EN ) 
                 RTL___csr_regfile___rg_dcsr  <= RTL___csr_regfile___rg_dcsr$D_IN ;
             if ( RTL___csr_regfile___rg_dpc$EN ) 
                 RTL___csr_regfile___rg_dpc  <= RTL___csr_regfile___rg_dpc$D_IN ;
             if ( RTL___csr_regfile___rg_dscratch0$EN ) 
                 RTL___csr_regfile___rg_dscratch0  <= RTL___csr_regfile___rg_dscratch0$D_IN ;
             if ( RTL___csr_regfile___rg_dscratch1$EN ) 
                 RTL___csr_regfile___rg_dscratch1  <= RTL___csr_regfile___rg_dscratch1$D_IN ;
             if ( RTL___csr_regfile___rg_mcause$EN ) 
                 RTL___csr_regfile___rg_mcause  <= RTL___csr_regfile___rg_mcause$D_IN ;
             if ( RTL___csr_regfile___rg_mcounteren$EN ) 
                 RTL___csr_regfile___rg_mcounteren  <= RTL___csr_regfile___rg_mcounteren$D_IN ;
             if ( RTL___csr_regfile___rg_mepc$EN ) 
                 RTL___csr_regfile___rg_mepc  <= RTL___csr_regfile___rg_mepc$D_IN ;
             if ( RTL___csr_regfile___rg_mscratch$EN ) 
                 RTL___csr_regfile___rg_mscratch  <= RTL___csr_regfile___rg_mscratch$D_IN ;
             if ( RTL___csr_regfile___rg_mtval$EN ) 
                 RTL___csr_regfile___rg_mtval  <= RTL___csr_regfile___rg_mtval$D_IN ;
             if ( RTL___csr_regfile___rg_mtvec$EN ) 
                 RTL___csr_regfile___rg_mtvec  <= RTL___csr_regfile___rg_mtvec$D_IN ;
             if ( RTL___csr_regfile___rg_nmi_vector$EN ) 
                 RTL___csr_regfile___rg_nmi_vector  <= RTL___csr_regfile___rg_nmi_vector$D_IN ;
             if ( RTL___csr_regfile___rg_tdata1$EN ) 
                 RTL___csr_regfile___rg_tdata1  <= RTL___csr_regfile___rg_tdata1$D_IN ;
             if ( RTL___csr_regfile___rg_tdata2$EN ) 
                 RTL___csr_regfile___rg_tdata2  <= RTL___csr_regfile___rg_tdata2$D_IN ;
             if ( RTL___csr_regfile___rg_tdata3$EN ) 
                 RTL___csr_regfile___rg_tdata3  <= RTL___csr_regfile___rg_tdata3$D_IN ;
             if ( RTL___csr_regfile___rg_tselect$EN ) 
                 RTL___csr_regfile___rg_tselect  <= RTL___csr_regfile___rg_tselect$D_IN ;
         end
  always @( negedge  RTL___csr_regfile___CLK )
         begin #0;
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_debug )$display("mstatus = 0x%0h", RTL___csr_regfile___csr_mstatus_rg_mstatus );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_debug )$display("mip     = 0x%0h", RTL___csr_regfile___csr_mip$fv_read );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_debug )$display("mie     = 0x%0h", RTL___csr_regfile___csr_mie$fv_read );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_Regfile.csr_trap_actions:", RTL___csr_regfile___rg_mcycle );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("    from priv %0d  pc 0x%0h  interrupt %0d  exc_code %0d  xtval 0x%0h", RTL___csr_regfile___csr_trap_actions_from_priv , RTL___csr_regfile___csr_trap_actions_pc , RTL___csr_regfile___csr_trap_actions_interrupt , RTL___csr_regfile___csr_trap_actions_exc_code , RTL___csr_regfile___csr_trap_actions_xtval );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("    priv %0d: ",2'b11);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ip: 0x%0h", RTL___csr_regfile___csr_mip$fv_read );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ie: 0x%0h", RTL___csr_regfile___csr_mie$fv_read );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" edeleg: 0x%0h",16'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ideleg: 0x%0h",12'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" cause:");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd0)$write("USER_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd1)$write("SUPERVISOR_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd2)$write("HYPERVISOR_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd3)$write("MACHINE_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd4)$write("USER_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd5)$write("SUPERVISOR_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd6)$write("HYPERVISOR_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd7)$write("MACHINE_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd8)$write("USER_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd9)$write("SUPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd10)$write("HYPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd11)$write("MACHINE_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]!=4'd0&& RTL___csr_regfile___rg_mcause [3:0]!=4'd1&& RTL___csr_regfile___rg_mcause [3:0]!=4'd2&& RTL___csr_regfile___rg_mcause [3:0]!=4'd3&& RTL___csr_regfile___rg_mcause [3:0]!=4'd4&& RTL___csr_regfile___rg_mcause [3:0]!=4'd5&& RTL___csr_regfile___rg_mcause [3:0]!=4'd6&& RTL___csr_regfile___rg_mcause [3:0]!=4'd7&& RTL___csr_regfile___rg_mcause [3:0]!=4'd8&& RTL___csr_regfile___rg_mcause [3:0]!=4'd9&& RTL___csr_regfile___rg_mcause [3:0]!=4'd10&& RTL___csr_regfile___rg_mcause [3:0]!=4'd11)$write("unknown interrupt Exc_Code %d", RTL___csr_regfile___rg_mcause [3:0]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd0)$write("INSTRUCTION_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd1)$write("INSTRUCTION_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd2)$write("ILLEGAL_INSTRUCTION");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd3)$write("BREAKPOINT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd4)$write("LOAD_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd5)$write("LOAD_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd6)$write("STORE_AMO_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd7)$write("STORE_AMO_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd8)$write("ECALL_FROM_U");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd9)$write("ECALL_FROM_S");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd11)$write("ECALL_FROM_M");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd12)$write("INSTRUCTION_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd13)$write("LOAD_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]==4'd15)$write("STORE_AMO_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___rg_mcause [4]&& RTL___csr_regfile___rg_mcause [3:0]!=4'd0&& RTL___csr_regfile___rg_mcause [3:0]!=4'd1&& RTL___csr_regfile___rg_mcause [3:0]!=4'd2&& RTL___csr_regfile___rg_mcause [3:0]!=4'd3&& RTL___csr_regfile___rg_mcause [3:0]!=4'd4&& RTL___csr_regfile___rg_mcause [3:0]!=4'd5&& RTL___csr_regfile___rg_mcause [3:0]!=4'd6&& RTL___csr_regfile___rg_mcause [3:0]!=4'd7&& RTL___csr_regfile___rg_mcause [3:0]!=4'd8&& RTL___csr_regfile___rg_mcause [3:0]!=4'd9&& RTL___csr_regfile___rg_mcause [3:0]!=4'd11&& RTL___csr_regfile___rg_mcause [3:0]!=4'd12&& RTL___csr_regfile___rg_mcause [3:0]!=4'd13&& RTL___csr_regfile___rg_mcause [3:0]!=4'd15)$write("unknown trap Exc_Code %d", RTL___csr_regfile___rg_mcause [3:0]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("        ");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" status: 0x%0h", RTL___csr_regfile___csr_mstatus_rg_mstatus );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tvec: 0x%0h",{ RTL___csr_regfile___rg_mtvec [30:1],1'b0, RTL___csr_regfile___rg_mtvec [0]});
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" epc: 0x%0h", RTL___csr_regfile___rg_mepc );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tval: 0x%0h", RTL___csr_regfile___rg_mtval );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("    Return: new pc 0x%0h  ", RTL___csr_regfile___x__h5843 );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new mstatus:");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("MStatus{","sd:%0d",1'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tsr:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [22]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tw:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [21]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" tvm:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [20]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mxr:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [19]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" sum:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [18]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mprv:%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [17]);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" xs:%0d",2'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" fs:%0d",2'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" mpp:%0d", RTL___csr_regfile___mpp__h7337 );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" spp:%0d",1'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" pies:%0d_%0d%0d", RTL___csr_regfile___csr_mstatus_rg_mstatus [3],1'd0,1'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" ies:%0d_%0d%0d",1'd0,1'd0,1'd0);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write("}");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new xcause:");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd0)$write("USER_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd1)$write("SUPERVISOR_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd2)$write("HYPERVISOR_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd3)$write("MACHINE_SW_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd4)$write("USER_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd5)$write("SUPERVISOR_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd6)$write("HYPERVISOR_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd7)$write("MACHINE_TIMER_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd8)$write("USER_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd9)$write("SUPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd10)$write("HYPERVISOR_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&! RTL___csr_regfile___csr_trap_actions_nmi && RTL___csr_regfile___csr_trap_actions_interrupt && RTL___csr_regfile___exc_code__h7909 ==4'd11)$write("MACHINE_EXTERNAL_INTERRUPT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___NOT_csr_trap_actions_nmi_97_AND_csr_trap_actio_ETC___d974 )$write("unknown interrupt Exc_Code %d", RTL___csr_regfile___exc_code__h7909 );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd0)$write("INSTRUCTION_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd1)$write("INSTRUCTION_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd2)$write("ILLEGAL_INSTRUCTION");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd3)$write("BREAKPOINT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd4)$write("LOAD_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd5)$write("LOAD_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd6)$write("STORE_AMO_ADDR_MISALIGNED");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd7)$write("STORE_AMO_ACCESS_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd8)$write("ECALL_FROM_U");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd9)$write("ECALL_FROM_S");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd11)$write("ECALL_FROM_M");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd12)$write("INSTRUCTION_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd13)$write("LOAD_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 &&( RTL___csr_regfile___csr_trap_actions_nmi ||! RTL___csr_regfile___csr_trap_actions_interrupt )&& RTL___csr_regfile___exc_code__h7909 ==4'd15)$write("STORE_AMO_PAGE_FAULT");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 && RTL___csr_regfile___csr_trap_actions_nmi_OR_NOT_csr_trap_actions_i_ETC___d1025 )$write("unknown trap Exc_Code %d", RTL___csr_regfile___exc_code__h7909 );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$write(" new priv %0d",2'b11);
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_csr_trap_actions && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("");
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___EN_mav_csr_write && RTL___csr_regfile___mav_csr_write_csr_addr_ULT_0xB03_77_OR_NOT_mav_ETC___d730 && RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: ERROR: CSR-write addr 0x%0h val 0x%0h not successful", RTL___csr_regfile___rg_mcycle , RTL___csr_regfile___mav_csr_write_csr_addr , RTL___csr_regfile___mav_csr_write_word );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: m_external_interrupt_req: %x", RTL___csr_regfile___rg_mcycle , RTL___csr_regfile___m_external_interrupt_req_set_not_clear );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: s_external_interrupt_req: %x", RTL___csr_regfile___rg_mcycle , RTL___csr_regfile___s_external_interrupt_req_set_not_clear );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: software_interrupt_req: %x", RTL___csr_regfile___rg_mcycle , RTL___csr_regfile___software_interrupt_req_set_not_clear );
             if ( RTL___csr_regfile___RST_N !=1'b0)
                 if ( RTL___csr_regfile___NOT_cfg_verbosity_read__31_ULE_1_32___d733 )$display("%0d: CSR_RegFile: timer_interrupt_req: %x", RTL___csr_regfile___rg_mcycle , RTL___csr_regfile___timer_interrupt_req_set_not_clear );
         end
  assign  RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_state = RTL___csr_regfile___rg_state ; 
  assign  RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_nmi = RTL___csr_regfile___rg_nmi ;
    assign RTL___RTL__DOT__csr_regfile__DOT__rg_nmi = RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_nmi;
    assign RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__csr_regfile__DOT__rg_state = RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__rg_state;
    assign RTL___csr_regfile___CLK = RTL___CLK;
    assign RTL___csr_regfile___RST_N = RTL___RST_N;
    assign RTL___csr_regfile___EN_server_reset_request_put = RTL___csr_regfile$EN_server_reset_request_put;
    assign RTL___csr_regfile$RDY_server_reset_request_put = RTL___csr_regfile___RDY_server_reset_request_put;
    assign RTL___csr_regfile___EN_server_reset_response_get = RTL___csr_regfile$EN_server_reset_response_get;
    assign RTL___csr_regfile$RDY_server_reset_response_get = RTL___csr_regfile___RDY_server_reset_response_get;
    assign RTL___csr_regfile___read_csr_csr_addr = RTL___csr_regfile$read_csr_csr_addr;
    assign RTL___csr_regfile$read_csr = RTL___csr_regfile___read_csr;
    assign RTL___csr_regfile___read_csr_port2_csr_addr = RTL___csr_regfile$read_csr_port2_csr_addr;
    assign RTL___csr_regfile___mav_read_csr_csr_addr = RTL___csr_regfile$mav_read_csr_csr_addr;
    assign RTL___csr_regfile___EN_mav_read_csr = RTL___csr_regfile$EN_mav_read_csr;
    assign RTL___csr_regfile___mav_csr_write_csr_addr = RTL___csr_regfile$mav_csr_write_csr_addr;
    assign RTL___csr_regfile___mav_csr_write_word = RTL___csr_regfile$mav_csr_write_word;
    assign RTL___csr_regfile___EN_mav_csr_write = RTL___csr_regfile$EN_mav_csr_write;
    assign RTL___csr_regfile$read_misa = RTL___csr_regfile___read_misa;
    assign RTL___csr_regfile$read_mstatus = RTL___csr_regfile___read_mstatus;
    assign RTL___csr_regfile$read_satp = RTL___csr_regfile___read_satp;
    assign RTL___csr_regfile___csr_trap_actions_from_priv = RTL___csr_regfile$csr_trap_actions_from_priv;
    assign RTL___csr_regfile___csr_trap_actions_pc = RTL___csr_regfile$csr_trap_actions_pc;
    assign RTL___csr_regfile___csr_trap_actions_nmi = RTL___csr_regfile$csr_trap_actions_nmi;
    assign RTL___csr_regfile___csr_trap_actions_interrupt = RTL___csr_regfile$csr_trap_actions_interrupt;
    assign RTL___csr_regfile___csr_trap_actions_exc_code = RTL___csr_regfile$csr_trap_actions_exc_code;
    assign RTL___csr_regfile___csr_trap_actions_xtval = RTL___csr_regfile$csr_trap_actions_xtval;
    assign RTL___csr_regfile___EN_csr_trap_actions = RTL___csr_regfile$EN_csr_trap_actions;
    assign RTL___csr_regfile$csr_trap_actions = RTL___csr_regfile___csr_trap_actions;
    assign RTL___csr_regfile___csr_ret_actions_from_priv = RTL___csr_regfile$csr_ret_actions_from_priv;
    assign RTL___csr_regfile___EN_csr_ret_actions = RTL___csr_regfile$EN_csr_ret_actions;
    assign RTL___csr_regfile$csr_ret_actions = RTL___csr_regfile___csr_ret_actions;
    assign RTL___csr_regfile$read_csr_minstret = RTL___csr_regfile___read_csr_minstret;
    assign RTL___csr_regfile___EN_csr_minstret_incr = RTL___csr_regfile$EN_csr_minstret_incr;
    assign RTL___csr_regfile$read_csr_mcycle = RTL___csr_regfile___read_csr_mcycle;
    assign RTL___csr_regfile___access_permitted_1_priv = RTL___csr_regfile$access_permitted_1_priv;
    assign RTL___csr_regfile___access_permitted_1_csr_addr = RTL___csr_regfile$access_permitted_1_csr_addr;
    assign RTL___csr_regfile___access_permitted_1_read_not_write = RTL___csr_regfile$access_permitted_1_read_not_write;
    assign RTL___csr_regfile$access_permitted_1 = RTL___csr_regfile___access_permitted_1;
    assign RTL___csr_regfile___access_permitted_2_priv = RTL___csr_regfile$access_permitted_2_priv;
    assign RTL___csr_regfile___access_permitted_2_csr_addr = RTL___csr_regfile$access_permitted_2_csr_addr;
    assign RTL___csr_regfile___access_permitted_2_read_not_write = RTL___csr_regfile$access_permitted_2_read_not_write;
    assign RTL___csr_regfile$access_permitted_2 = RTL___csr_regfile___access_permitted_2;
    assign RTL___csr_regfile___csr_counter_read_fault_priv = RTL___csr_regfile$csr_counter_read_fault_priv;
    assign RTL___csr_regfile___csr_counter_read_fault_csr_addr = RTL___csr_regfile$csr_counter_read_fault_csr_addr;
    assign RTL___csr_regfile___m_external_interrupt_req_set_not_clear = RTL___csr_regfile$m_external_interrupt_req_set_not_clear;
    assign RTL___csr_regfile___s_external_interrupt_req_set_not_clear = RTL___csr_regfile$s_external_interrupt_req_set_not_clear;
    assign RTL___csr_regfile___timer_interrupt_req_set_not_clear = RTL___csr_regfile$timer_interrupt_req_set_not_clear;
    assign RTL___csr_regfile___software_interrupt_req_set_not_clear = RTL___csr_regfile$software_interrupt_req_set_not_clear;
    assign RTL___csr_regfile___interrupt_pending_cur_priv = RTL___csr_regfile$interrupt_pending_cur_priv;
    assign RTL___csr_regfile$interrupt_pending = RTL___csr_regfile___interrupt_pending;
    assign RTL___csr_regfile$wfi_resume = RTL___csr_regfile___wfi_resume;
    assign RTL___csr_regfile___nmi_req_set_not_clear = RTL___csr_regfile$nmi_req_set_not_clear;
    assign RTL___csr_regfile$nmi_pending = RTL___csr_regfile___nmi_pending;
    assign RTL___csr_regfile___EN_debug = RTL___csr_regfile$EN_debug;
      
    wire RTL___f_reset_reqs___CLK;
    wire RTL___f_reset_reqs___RST;
    wire[RTL___f_reset_reqs___width-1:0] RTL___f_reset_reqs___D_IN;
    wire RTL___f_reset_reqs___ENQ;
    wire RTL___f_reset_reqs___DEQ;
    wire RTL___f_reset_reqs___CLR;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_reqs___FULL_N;
    wire RTL___f_reset_reqs___EMPTY_N;
    wire[RTL___f_reset_reqs___width-1:0] RTL___f_reset_reqs___D_OUT;
    wire RTL___f_reset_rsps___CLK;
    wire RTL___f_reset_rsps___RST;
    wire[RTL___f_reset_rsps___width-1:0] RTL___f_reset_rsps___D_IN;
    wire RTL___f_reset_rsps___ENQ;
    wire RTL___f_reset_rsps___DEQ;
    wire RTL___f_reset_rsps___CLR;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___f_reset_rsps___FULL_N;
    wire RTL___f_reset_rsps___EMPTY_N;
    wire[RTL___f_reset_rsps___width-1:0] RTL___f_reset_rsps___D_OUT;

    reg RTL___f_reset_reqs___full_reg ; 
    reg RTL___f_reset_reqs___empty_reg ; reg[ RTL___f_reset_reqs___width -1:0] RTL___f_reset_reqs___data0_reg ; reg[ RTL___f_reset_reqs___width -1:0] RTL___f_reset_reqs___data1_reg ; 
  assign  RTL___f_reset_reqs___FULL_N = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___EMPTY_N = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___D_OUT = RTL___f_reset_reqs___data0_reg ; 
    wire RTL___f_reset_reqs___d0di =( RTL___f_reset_reqs___ENQ &&! RTL___f_reset_reqs___empty_reg )||( RTL___f_reset_reqs___ENQ && RTL___f_reset_reqs___DEQ && RTL___f_reset_reqs___full_reg ); 
    wire RTL___f_reset_reqs___d0d1 = RTL___f_reset_reqs___DEQ &&! RTL___f_reset_reqs___full_reg ; 
    wire RTL___f_reset_reqs___d0h =((! RTL___f_reset_reqs___DEQ )&&(! RTL___f_reset_reqs___ENQ ))||(! RTL___f_reset_reqs___DEQ && RTL___f_reset_reqs___empty_reg )||(! RTL___f_reset_reqs___ENQ && RTL___f_reset_reqs___full_reg ); 
    wire RTL___f_reset_reqs___d1di = RTL___f_reset_reqs___ENQ & RTL___f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___f_reset_reqs___CLK )
         begin 
             if ( RTL___f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___f_reset_reqs___CLR )
                         begin  
                             RTL___f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___f_reset_reqs___ENQ &&! RTL___f_reset_reqs___DEQ )
                             begin  
                                 RTL___f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___f_reset_reqs___full_reg  <=! RTL___f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if ( RTL___f_reset_reqs___DEQ &&! RTL___f_reset_reqs___ENQ )
                                 begin  
                                     RTL___f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___f_reset_reqs___empty_reg  <=! RTL___f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___f_reset_reqs___CLK )
         begin 
             begin  
                 RTL___f_reset_reqs___data0_reg  <={ RTL___f_reset_reqs___width { RTL___f_reset_reqs___d0di }}& RTL___f_reset_reqs___D_IN |{ RTL___f_reset_reqs___width { RTL___f_reset_reqs___d0d1 }}& RTL___f_reset_reqs___data1_reg |{ RTL___f_reset_reqs___width { RTL___f_reset_reqs___d0h }}& RTL___f_reset_reqs___data0_reg ; 
                 RTL___f_reset_reqs___data1_reg  <= RTL___f_reset_reqs___d1di  ?  RTL___f_reset_reqs___D_IN : RTL___f_reset_reqs___data1_reg ;
             end 
         end
  always @( posedge  RTL___f_reset_reqs___CLK )
         begin : RTL___f_reset_reqs___error_checks 
           reg RTL___f_reset_reqs___deqerror , RTL___f_reset_reqs___enqerror ; 
             RTL___f_reset_reqs___deqerror  =0; 
             RTL___f_reset_reqs___enqerror  =0;
             if ( RTL___f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___f_reset_reqs___empty_reg && RTL___f_reset_reqs___DEQ )
                         begin  
                             RTL___f_reset_reqs___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___f_reset_reqs___full_reg && RTL___f_reset_reqs___ENQ &&(! RTL___f_reset_reqs___DEQ || RTL___f_reset_reqs___guarded ))
                         begin  
                             RTL___f_reset_reqs___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___f_reset_reqs___full_reg ; 
  assign  RTL___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___f_reset_reqs___empty_reg ;
    reg RTL___f_reset_rsps___full_reg ; 
    reg RTL___f_reset_rsps___empty_reg ; reg[ RTL___f_reset_rsps___width -1:0] RTL___f_reset_rsps___data0_reg ; reg[ RTL___f_reset_rsps___width -1:0] RTL___f_reset_rsps___data1_reg ; 
  assign  RTL___f_reset_rsps___FULL_N = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___EMPTY_N = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___D_OUT = RTL___f_reset_rsps___data0_reg ; 
    wire RTL___f_reset_rsps___d0di =( RTL___f_reset_rsps___ENQ &&! RTL___f_reset_rsps___empty_reg )||( RTL___f_reset_rsps___ENQ && RTL___f_reset_rsps___DEQ && RTL___f_reset_rsps___full_reg ); 
    wire RTL___f_reset_rsps___d0d1 = RTL___f_reset_rsps___DEQ &&! RTL___f_reset_rsps___full_reg ; 
    wire RTL___f_reset_rsps___d0h =((! RTL___f_reset_rsps___DEQ )&&(! RTL___f_reset_rsps___ENQ ))||(! RTL___f_reset_rsps___DEQ && RTL___f_reset_rsps___empty_reg )||(! RTL___f_reset_rsps___ENQ && RTL___f_reset_rsps___full_reg ); 
    wire RTL___f_reset_rsps___d1di = RTL___f_reset_rsps___ENQ & RTL___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___f_reset_rsps___CLK )
         begin 
             if ( RTL___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___f_reset_rsps___CLR )
                         begin  
                             RTL___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___f_reset_rsps___ENQ &&! RTL___f_reset_rsps___DEQ )
                             begin  
                                 RTL___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___f_reset_rsps___full_reg  <=! RTL___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if ( RTL___f_reset_rsps___DEQ &&! RTL___f_reset_rsps___ENQ )
                                 begin  
                                     RTL___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___f_reset_rsps___empty_reg  <=! RTL___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___f_reset_rsps___CLK )
         begin 
             begin  
                 RTL___f_reset_rsps___data0_reg  <={ RTL___f_reset_rsps___width { RTL___f_reset_rsps___d0di }}& RTL___f_reset_rsps___D_IN |{ RTL___f_reset_rsps___width { RTL___f_reset_rsps___d0d1 }}& RTL___f_reset_rsps___data1_reg |{ RTL___f_reset_rsps___width { RTL___f_reset_rsps___d0h }}& RTL___f_reset_rsps___data0_reg ; 
                 RTL___f_reset_rsps___data1_reg  <= RTL___f_reset_rsps___d1di  ?  RTL___f_reset_rsps___D_IN : RTL___f_reset_rsps___data1_reg ;
             end 
         end
  always @( posedge  RTL___f_reset_rsps___CLK )
         begin : RTL___f_reset_rsps___error_checks 
           reg RTL___f_reset_rsps___deqerror , RTL___f_reset_rsps___enqerror ; 
             RTL___f_reset_rsps___deqerror  =0; 
             RTL___f_reset_rsps___enqerror  =0;
             if ( RTL___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___f_reset_rsps___empty_reg && RTL___f_reset_rsps___DEQ )
                         begin  
                             RTL___f_reset_rsps___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___f_reset_rsps___full_reg && RTL___f_reset_rsps___ENQ &&(! RTL___f_reset_rsps___DEQ || RTL___f_reset_rsps___guarded ))
                         begin  
                             RTL___f_reset_rsps___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___f_reset_rsps___full_reg ; 
  assign  RTL___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___f_reset_rsps___empty_reg ;
    assign RTL___f_reset_reqs___CLK = RTL___CLK;
    assign RTL___f_reset_reqs___RST = RTL___RST_N;
    assign RTL___f_reset_reqs___D_IN = RTL___f_reset_reqs$D_IN;
    assign RTL___f_reset_reqs___ENQ = RTL___f_reset_reqs$ENQ;
    assign RTL___f_reset_reqs___DEQ = RTL___f_reset_reqs$DEQ;
    assign RTL___f_reset_reqs___CLR = RTL___f_reset_reqs$CLR;
    assign RTL___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___f_reset_reqs$FULL_N = RTL___f_reset_reqs___FULL_N;
    assign RTL___f_reset_reqs$EMPTY_N = RTL___f_reset_reqs___EMPTY_N;
    assign RTL___f_reset_reqs$D_OUT = RTL___f_reset_reqs___D_OUT;
    assign RTL___f_reset_rsps___CLK = RTL___CLK;
    assign RTL___f_reset_rsps___RST = RTL___RST_N;
    assign RTL___f_reset_rsps___D_IN = RTL___f_reset_rsps$D_IN;
    assign RTL___f_reset_rsps___ENQ = RTL___f_reset_rsps$ENQ;
    assign RTL___f_reset_rsps___DEQ = RTL___f_reset_rsps$DEQ;
    assign RTL___f_reset_rsps___CLR = RTL___f_reset_rsps$CLR;
    assign RTL___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___f_reset_rsps$FULL_N = RTL___f_reset_rsps___FULL_N;
    assign RTL___f_reset_rsps$EMPTY_N = RTL___f_reset_rsps___EMPTY_N;
    assign RTL___f_reset_rsps$D_OUT = RTL___f_reset_rsps___D_OUT;
      
    wire RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire RTL___gpr_regfile___CLK;
    wire RTL___gpr_regfile___RST_N;
    wire RTL___gpr_regfile___EN_server_reset_request_put;
    wire RTL___gpr_regfile___EN_server_reset_response_get;
    wire[4:0] RTL___gpr_regfile___read_rs1_rs1;
    wire[4:0] RTL___gpr_regfile___read_rs1_port2_rs1;
    wire[4:0] RTL___gpr_regfile___read_rs2_rs2;
    wire[4:0] RTL___gpr_regfile___write_rd_rd;
    wire[31:0] RTL___gpr_regfile___write_rd_rd_val;
    wire RTL___gpr_regfile___EN_write_rd;

    wire[31:0] RTL___gpr_regfile___read_rs1 , RTL___gpr_regfile___read_rs1_port2 , RTL___gpr_regfile___read_rs2 ; 
    wire RTL___gpr_regfile___RDY_server_reset_request_put , RTL___gpr_regfile___RDY_server_reset_response_get ; reg[1:0] RTL___gpr_regfile___rg_state ; reg[1:0] RTL___gpr_regfile___rg_state$D_IN ; 
    wire RTL___gpr_regfile___rg_state$EN ; 
    wire RTL___gpr_regfile___f_reset_rsps$CLR , RTL___gpr_regfile___f_reset_rsps$DEQ , RTL___gpr_regfile___f_reset_rsps$EMPTY_N , RTL___gpr_regfile___f_reset_rsps$ENQ , RTL___gpr_regfile___f_reset_rsps$FULL_N ; 
    wire[31:0] RTL___gpr_regfile___regfile$D_IN , RTL___gpr_regfile___regfile$D_OUT_1 , RTL___gpr_regfile___regfile$D_OUT_2 , RTL___gpr_regfile___regfile$D_OUT_3 ; 
    wire[4:0] RTL___gpr_regfile___regfile$ADDR_1 , RTL___gpr_regfile___regfile$ADDR_2 , RTL___gpr_regfile___regfile$ADDR_3 , RTL___gpr_regfile___regfile$ADDR_4 , RTL___gpr_regfile___regfile$ADDR_5 , RTL___gpr_regfile___regfile$ADDR_IN ; 
    wire RTL___gpr_regfile___regfile$WE ; 
    wire RTL___gpr_regfile___CAN_FIRE_RL_rl_reset_loop , RTL___gpr_regfile___CAN_FIRE_RL_rl_reset_start , RTL___gpr_regfile___CAN_FIRE_server_reset_request_put , RTL___gpr_regfile___CAN_FIRE_server_reset_response_get , RTL___gpr_regfile___CAN_FIRE_write_rd , RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_loop , RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_start , RTL___gpr_regfile___WILL_FIRE_server_reset_request_put , RTL___gpr_regfile___WILL_FIRE_server_reset_response_get , RTL___gpr_regfile___WILL_FIRE_write_rd ; 
  assign  RTL___gpr_regfile___RDY_server_reset_request_put = RTL___gpr_regfile___f_reset_rsps$FULL_N ; 
  assign  RTL___gpr_regfile___CAN_FIRE_server_reset_request_put = RTL___gpr_regfile___f_reset_rsps$FULL_N ; 
  assign  RTL___gpr_regfile___WILL_FIRE_server_reset_request_put = RTL___gpr_regfile___EN_server_reset_request_put ; 
  assign  RTL___gpr_regfile___RDY_server_reset_response_get = RTL___gpr_regfile___rg_state ==2'd2&& RTL___gpr_regfile___f_reset_rsps$EMPTY_N ; 
  assign  RTL___gpr_regfile___CAN_FIRE_server_reset_response_get = RTL___gpr_regfile___rg_state ==2'd2&& RTL___gpr_regfile___f_reset_rsps$EMPTY_N ; 
  assign  RTL___gpr_regfile___WILL_FIRE_server_reset_response_get = RTL___gpr_regfile___EN_server_reset_response_get ; 
  assign  RTL___gpr_regfile___read_rs1 =( RTL___gpr_regfile___read_rs1_rs1 ==5'd0) ? 32'd0: RTL___gpr_regfile___regfile$D_OUT_3 ; 
  assign  RTL___gpr_regfile___read_rs1_port2 =( RTL___gpr_regfile___read_rs1_port2_rs1 ==5'd0) ? 32'd0: RTL___gpr_regfile___regfile$D_OUT_2 ; 
  assign  RTL___gpr_regfile___read_rs2 =( RTL___gpr_regfile___read_rs2_rs2 ==5'd0) ? 32'd0: RTL___gpr_regfile___regfile$D_OUT_1 ; 
  assign  RTL___gpr_regfile___CAN_FIRE_write_rd =1'd1; 
  assign  RTL___gpr_regfile___WILL_FIRE_write_rd = RTL___gpr_regfile___EN_write_rd ;  
    wire RTL___gpr_regfile___f_reset_rsps___RST;
    wire RTL___gpr_regfile___f_reset_rsps___CLK;
    wire RTL___gpr_regfile___f_reset_rsps___ENQ;
    wire RTL___gpr_regfile___f_reset_rsps___CLR;
    wire RTL___gpr_regfile___f_reset_rsps___DEQ;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___gpr_regfile___f_reset_rsps___FULL_N;
    wire RTL___gpr_regfile___f_reset_rsps___EMPTY_N;

    reg RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
    reg RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___FULL_N = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___EMPTY_N = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___gpr_regfile___f_reset_rsps___CLK )
         begin 
             if ( RTL___gpr_regfile___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___gpr_regfile___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___gpr_regfile___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___gpr_regfile___f_reset_rsps___CLR )
                         begin  
                             RTL___gpr_regfile___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___gpr_regfile___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___gpr_regfile___f_reset_rsps___ENQ &&! RTL___gpr_regfile___f_reset_rsps___DEQ )
                             begin  
                                 RTL___gpr_regfile___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___gpr_regfile___f_reset_rsps___full_reg  <=! RTL___gpr_regfile___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___gpr_regfile___f_reset_rsps___ENQ && RTL___gpr_regfile___f_reset_rsps___DEQ )
                                 begin  
                                     RTL___gpr_regfile___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___gpr_regfile___f_reset_rsps___empty_reg  <=! RTL___gpr_regfile___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___gpr_regfile___f_reset_rsps___CLK )
         begin : RTL___gpr_regfile___f_reset_rsps___error_checks 
           reg RTL___gpr_regfile___f_reset_rsps___deqerror , RTL___gpr_regfile___f_reset_rsps___enqerror ; 
             RTL___gpr_regfile___f_reset_rsps___deqerror  =0; 
             RTL___gpr_regfile___f_reset_rsps___enqerror  =0;
             if ( RTL___gpr_regfile___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___gpr_regfile___f_reset_rsps___empty_reg && RTL___gpr_regfile___f_reset_rsps___DEQ )
                         begin  
                             RTL___gpr_regfile___f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___gpr_regfile___f_reset_rsps___full_reg && RTL___gpr_regfile___f_reset_rsps___ENQ &&(! RTL___gpr_regfile___f_reset_rsps___DEQ || RTL___gpr_regfile___f_reset_rsps___guarded ))
                         begin  
                             RTL___gpr_regfile___f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___full_reg ; 
  assign  RTL___gpr_regfile___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___empty_reg ;
    assign RTL___gpr_regfile___f_reset_rsps___RST = RTL___gpr_regfile___RST_N;
    assign RTL___gpr_regfile___f_reset_rsps___CLK = RTL___gpr_regfile___CLK;
    assign RTL___gpr_regfile___f_reset_rsps___ENQ = RTL___gpr_regfile___f_reset_rsps$ENQ;
    assign RTL___gpr_regfile___f_reset_rsps___CLR = RTL___gpr_regfile___f_reset_rsps$CLR;
    assign RTL___gpr_regfile___f_reset_rsps___DEQ = RTL___gpr_regfile___f_reset_rsps$DEQ;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___gpr_regfile___f_reset_rsps$FULL_N = RTL___gpr_regfile___f_reset_rsps___FULL_N;
    assign RTL___gpr_regfile___f_reset_rsps$EMPTY_N = RTL___gpr_regfile___f_reset_rsps___EMPTY_N;
      
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    wire[31:0] RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    wire RTL___gpr_regfile___regfile___CLK;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_IN;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_IN;
    wire RTL___gpr_regfile___regfile___WE;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_1;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_OUT_1;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_2;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_OUT_2;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_3;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_OUT_3;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_4;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_OUT_4;
    wire[RTL___gpr_regfile___regfile___addr_width-1:0] RTL___gpr_regfile___regfile___ADDR_5;
    wire[RTL___gpr_regfile___regfile___data_width-1:0] RTL___gpr_regfile___regfile___D_OUT_5;

    reg[ RTL___gpr_regfile___regfile___data_width -1:0] RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___lo : RTL___gpr_regfile___regfile___hi ]; 
  always @( posedge  RTL___gpr_regfile___regfile___CLK )
         begin 
             if ( RTL___gpr_regfile___regfile___WE ) 
                 RTL___gpr_regfile___regfile___arr  [ RTL___gpr_regfile___regfile___ADDR_IN ]<= RTL___gpr_regfile___regfile___D_IN ;
         end
  assign  RTL___gpr_regfile___regfile___D_OUT_1 = RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___ADDR_1 ]; 
  assign  RTL___gpr_regfile___regfile___D_OUT_2 = RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___ADDR_2 ]; 
  assign  RTL___gpr_regfile___regfile___D_OUT_3 = RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___ADDR_3 ]; 
  assign  RTL___gpr_regfile___regfile___D_OUT_4 = RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___ADDR_4 ]; 
  assign  RTL___gpr_regfile___regfile___D_OUT_5 = RTL___gpr_regfile___regfile___arr [ RTL___gpr_regfile___regfile___ADDR_5 ]; 
  always @( posedge  RTL___gpr_regfile___regfile___CLK )
         begin : RTL___gpr_regfile___regfile___runtime_check 
           reg RTL___gpr_regfile___regfile___enable_check ; 
             RTL___gpr_regfile___regfile___enable_check  =0;
             if ( RTL___gpr_regfile___regfile___enable_check )
                 begin 
                     if (( RTL___gpr_regfile___regfile___ADDR_1 < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_1 > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Address port 1 is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_1 );
                     if (( RTL___gpr_regfile___regfile___ADDR_2 < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_2 > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Address port 2 is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_2 );
                     if (( RTL___gpr_regfile___regfile___ADDR_3 < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_3 > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Address port 3 is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_3 );
                     if (( RTL___gpr_regfile___regfile___ADDR_4 < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_4 > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Address port 4 is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_4 );
                     if (( RTL___gpr_regfile___regfile___ADDR_5 < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_5 > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Address port 5 is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_5 );
                     if ( RTL___gpr_regfile___regfile___WE &&( RTL___gpr_regfile___regfile___ADDR_IN < RTL___gpr_regfile___regfile___lo )||( RTL___gpr_regfile___regfile___ADDR_IN > RTL___gpr_regfile___regfile___hi ))$display("Warning: RegFile: %m -- Write Address port is out of bounds: %h", RTL___gpr_regfile___regfile___ADDR_IN );
                 end 
         end
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL___gpr_regfile___regfile___arr [15]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL___gpr_regfile___regfile___arr [12]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL___gpr_regfile___regfile___arr [7]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL___gpr_regfile___regfile___arr [10]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL___gpr_regfile___regfile___arr [1]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL___gpr_regfile___regfile___arr [6]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL___gpr_regfile___regfile___arr [31]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL___gpr_regfile___regfile___arr [29]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL___gpr_regfile___regfile___arr [27]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL___gpr_regfile___regfile___arr [25]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL___gpr_regfile___regfile___arr [23]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL___gpr_regfile___regfile___arr [22]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL___gpr_regfile___regfile___arr [21]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL___gpr_regfile___regfile___arr [18]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL___gpr_regfile___regfile___arr [16]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL___gpr_regfile___regfile___arr [28]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL___gpr_regfile___regfile___arr [2]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL___gpr_regfile___regfile___arr [24]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL___gpr_regfile___regfile___arr [30]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL___gpr_regfile___regfile___arr [26]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL___gpr_regfile___regfile___arr [13]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL___gpr_regfile___regfile___arr [19]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL___gpr_regfile___regfile___arr [5]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL___gpr_regfile___regfile___arr [20]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL___gpr_regfile___regfile___arr [4]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL___gpr_regfile___regfile___arr [11]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL___gpr_regfile___regfile___arr [8]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL___gpr_regfile___regfile___arr [3]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL___gpr_regfile___regfile___arr [9]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL___gpr_regfile___regfile___arr [14]; 
  assign  RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL___gpr_regfile___regfile___arr [17];
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL___gpr_regfile___regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL___gpr_regfile___regfile___CLK = RTL___gpr_regfile___CLK;
    assign RTL___gpr_regfile___regfile___ADDR_IN = RTL___gpr_regfile___regfile$ADDR_IN;
    assign RTL___gpr_regfile___regfile___D_IN = RTL___gpr_regfile___regfile$D_IN;
    assign RTL___gpr_regfile___regfile___WE = RTL___gpr_regfile___regfile$WE;
    assign RTL___gpr_regfile___regfile___ADDR_1 = RTL___gpr_regfile___regfile$ADDR_1;
    assign RTL___gpr_regfile___regfile$D_OUT_1 = RTL___gpr_regfile___regfile___D_OUT_1;
    assign RTL___gpr_regfile___regfile___ADDR_2 = RTL___gpr_regfile___regfile$ADDR_2;
    assign RTL___gpr_regfile___regfile$D_OUT_2 = RTL___gpr_regfile___regfile___D_OUT_2;
    assign RTL___gpr_regfile___regfile___ADDR_3 = RTL___gpr_regfile___regfile$ADDR_3;
    assign RTL___gpr_regfile___regfile$D_OUT_3 = RTL___gpr_regfile___regfile___D_OUT_3;
    assign RTL___gpr_regfile___regfile___ADDR_4 = RTL___gpr_regfile___regfile$ADDR_4;
    assign RTL___gpr_regfile___regfile___ADDR_5 = RTL___gpr_regfile___regfile$ADDR_5;
     
  assign  RTL___gpr_regfile___CAN_FIRE_RL_rl_reset_start = RTL___gpr_regfile___rg_state ==2'd0; 
  assign  RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_start = RTL___gpr_regfile___rg_state ==2'd0; 
  assign  RTL___gpr_regfile___CAN_FIRE_RL_rl_reset_loop = RTL___gpr_regfile___rg_state ==2'd1; 
  assign  RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_loop = RTL___gpr_regfile___rg_state ==2'd1; 
  always @(    RTL___gpr_regfile___EN_server_reset_request_put              or   RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_loop           or   RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_start  )
         case (1'b1) 
          RTL___gpr_regfile___EN_server_reset_request_put  : 
              RTL___gpr_regfile___rg_state$D_IN  =2'd0; 
          RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_loop  : 
              RTL___gpr_regfile___rg_state$D_IN  =2'd2; 
          RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_start  : 
              RTL___gpr_regfile___rg_state$D_IN  =2'd1;
          default : 
              RTL___gpr_regfile___rg_state$D_IN  =2'b10;endcase
  assign  RTL___gpr_regfile___rg_state$EN = RTL___gpr_regfile___EN_server_reset_request_put || RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_start || RTL___gpr_regfile___WILL_FIRE_RL_rl_reset_loop ; 
  assign  RTL___gpr_regfile___f_reset_rsps$ENQ = RTL___gpr_regfile___EN_server_reset_request_put ; 
  assign  RTL___gpr_regfile___f_reset_rsps$DEQ = RTL___gpr_regfile___EN_server_reset_response_get ; 
  assign  RTL___gpr_regfile___f_reset_rsps$CLR =1'b0; 
  assign  RTL___gpr_regfile___regfile$ADDR_1 = RTL___gpr_regfile___read_rs2_rs2 ; 
  assign  RTL___gpr_regfile___regfile$ADDR_2 = RTL___gpr_regfile___read_rs1_port2_rs1 ; 
  assign  RTL___gpr_regfile___regfile$ADDR_3 = RTL___gpr_regfile___read_rs1_rs1 ; 
  assign  RTL___gpr_regfile___regfile$ADDR_4 =5'h0; 
  assign  RTL___gpr_regfile___regfile$ADDR_5 =5'h0; 
  assign  RTL___gpr_regfile___regfile$ADDR_IN = RTL___gpr_regfile___write_rd_rd ; 
  assign  RTL___gpr_regfile___regfile$D_IN = RTL___gpr_regfile___write_rd_rd_val ; 
  assign  RTL___gpr_regfile___regfile$WE = RTL___gpr_regfile___EN_write_rd && RTL___gpr_regfile___write_rd_rd !=5'd0; 
  always @( posedge  RTL___gpr_regfile___CLK )
         begin 
             if ( RTL___gpr_regfile___RST_N ==1'b0)
                 begin  
                     RTL___gpr_regfile___rg_state  <=2'd0;
                 end 
              else 
                 begin 
                     if ( RTL___gpr_regfile___rg_state$EN ) 
                         RTL___gpr_regfile___rg_state  <= RTL___gpr_regfile___rg_state$D_IN ;
                 end 
         end
 
    assign RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL___gpr_regfile___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL___gpr_regfile___CLK = RTL___CLK;
    assign RTL___gpr_regfile___RST_N = RTL___RST_N;
    assign RTL___gpr_regfile___EN_server_reset_request_put = RTL___gpr_regfile$EN_server_reset_request_put;
    assign RTL___gpr_regfile$RDY_server_reset_request_put = RTL___gpr_regfile___RDY_server_reset_request_put;
    assign RTL___gpr_regfile___EN_server_reset_response_get = RTL___gpr_regfile$EN_server_reset_response_get;
    assign RTL___gpr_regfile$RDY_server_reset_response_get = RTL___gpr_regfile___RDY_server_reset_response_get;
    assign RTL___gpr_regfile___read_rs1_rs1 = RTL___gpr_regfile$read_rs1_rs1;
    assign RTL___gpr_regfile$read_rs1 = RTL___gpr_regfile___read_rs1;
    assign RTL___gpr_regfile___read_rs1_port2_rs1 = RTL___gpr_regfile$read_rs1_port2_rs1;
    assign RTL___gpr_regfile___read_rs2_rs2 = RTL___gpr_regfile$read_rs2_rs2;
    assign RTL___gpr_regfile$read_rs2 = RTL___gpr_regfile___read_rs2;
    assign RTL___gpr_regfile___write_rd_rd = RTL___gpr_regfile$write_rd_rd;
    assign RTL___gpr_regfile___write_rd_rd_val = RTL___gpr_regfile$write_rd_rd_val;
    assign RTL___gpr_regfile___EN_write_rd = RTL___gpr_regfile$EN_write_rd;
      
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___CLK;
    wire RTL___near_mem___RST_N;
    wire RTL___near_mem___EN_server_reset_request_put;
    wire RTL___near_mem___EN_server_reset_response_get;
    wire[2:0] RTL___near_mem___imem_req_f3;
    wire[31:0] RTL___near_mem___imem_req_addr;
    wire[1:0] RTL___near_mem___imem_req_priv;
    wire RTL___near_mem___imem_req_sstatus_SUM;
    wire RTL___near_mem___imem_req_mstatus_MXR;
    wire[31:0] RTL___near_mem___imem_req_satp;
    wire RTL___near_mem___EN_imem_req;
    wire RTL___near_mem___imem_master_awready;
    wire RTL___near_mem___imem_master_wready;
    wire RTL___near_mem___imem_master_bvalid;
    wire[3:0] RTL___near_mem___imem_master_bid;
    wire[1:0] RTL___near_mem___imem_master_bresp;
    wire RTL___near_mem___imem_master_arready;
    wire RTL___near_mem___imem_master_rvalid;
    wire[3:0] RTL___near_mem___imem_master_rid;
    wire[63:0] RTL___near_mem___imem_master_rdata;
    wire[1:0] RTL___near_mem___imem_master_rresp;
    wire RTL___near_mem___imem_master_rlast;
    wire RTL___near_mem___dmem_req_op;
    wire[2:0] RTL___near_mem___dmem_req_f3;
    wire[31:0] RTL___near_mem___dmem_req_addr;
    wire[63:0] RTL___near_mem___dmem_req_store_value;
    wire[1:0] RTL___near_mem___dmem_req_priv;
    wire RTL___near_mem___dmem_req_sstatus_SUM;
    wire RTL___near_mem___dmem_req_mstatus_MXR;
    wire[31:0] RTL___near_mem___dmem_req_satp;
    wire RTL___near_mem___EN_dmem_req;
    wire RTL___near_mem___dmem_master_awready;
    wire RTL___near_mem___dmem_master_wready;
    wire RTL___near_mem___dmem_master_bvalid;
    wire[3:0] RTL___near_mem___dmem_master_bid;
    wire[1:0] RTL___near_mem___dmem_master_bresp;
    wire RTL___near_mem___dmem_master_arready;
    wire RTL___near_mem___dmem_master_rvalid;
    wire[3:0] RTL___near_mem___dmem_master_rid;
    wire[63:0] RTL___near_mem___dmem_master_rdata;
    wire[1:0] RTL___near_mem___dmem_master_rresp;
    wire RTL___near_mem___dmem_master_rlast;
    wire RTL___near_mem___EN_server_fence_i_request_put;
    wire RTL___near_mem___EN_server_fence_i_response_get;
    wire[7:0] RTL___near_mem___server_fence_request_put;
    wire RTL___near_mem___EN_server_fence_request_put;
    wire RTL___near_mem___EN_server_fence_response_get;
    wire RTL___near_mem___EN_sfence_vma;

    wire[63:0] RTL___near_mem___dmem_master_araddr , RTL___near_mem___dmem_master_awaddr , RTL___near_mem___dmem_master_wdata , RTL___near_mem___dmem_st_amo_val , RTL___near_mem___dmem_word64 , RTL___near_mem___imem_master_araddr , RTL___near_mem___imem_master_awaddr , RTL___near_mem___imem_master_wdata ; 
    wire[31:0] RTL___near_mem___imem_instr , RTL___near_mem___imem_pc , RTL___near_mem___imem_tval ; 
    wire[7:0] RTL___near_mem___dmem_master_arlen , RTL___near_mem___dmem_master_awlen , RTL___near_mem___dmem_master_wstrb , RTL___near_mem___imem_master_arlen , RTL___near_mem___imem_master_awlen , RTL___near_mem___imem_master_wstrb ; 
    wire[3:0] RTL___near_mem___dmem_exc_code , RTL___near_mem___dmem_master_arcache , RTL___near_mem___dmem_master_arid , RTL___near_mem___dmem_master_arqos , RTL___near_mem___dmem_master_arregion , RTL___near_mem___dmem_master_awcache , RTL___near_mem___dmem_master_awid , RTL___near_mem___dmem_master_awqos , RTL___near_mem___dmem_master_awregion , RTL___near_mem___imem_exc_code , RTL___near_mem___imem_master_arcache , RTL___near_mem___imem_master_arid , RTL___near_mem___imem_master_arqos , RTL___near_mem___imem_master_arregion , RTL___near_mem___imem_master_awcache , RTL___near_mem___imem_master_awid , RTL___near_mem___imem_master_awqos , RTL___near_mem___imem_master_awregion ; 
    wire[2:0] RTL___near_mem___dmem_master_arprot , RTL___near_mem___dmem_master_arsize , RTL___near_mem___dmem_master_awprot , RTL___near_mem___dmem_master_awsize , RTL___near_mem___imem_master_arprot , RTL___near_mem___imem_master_arsize , RTL___near_mem___imem_master_awprot , RTL___near_mem___imem_master_awsize ; 
    wire[1:0] RTL___near_mem___dmem_master_arburst , RTL___near_mem___dmem_master_awburst , RTL___near_mem___imem_master_arburst , RTL___near_mem___imem_master_awburst ; 
    wire RTL___near_mem___RDY_server_fence_i_request_put , RTL___near_mem___RDY_server_fence_i_response_get , RTL___near_mem___RDY_server_fence_request_put , RTL___near_mem___RDY_server_fence_response_get , RTL___near_mem___RDY_server_reset_request_put , RTL___near_mem___RDY_server_reset_response_get , RTL___near_mem___RDY_sfence_vma , RTL___near_mem___dmem_exc , RTL___near_mem___dmem_master_arlock , RTL___near_mem___dmem_master_arvalid , RTL___near_mem___dmem_master_awlock , RTL___near_mem___dmem_master_awvalid , RTL___near_mem___dmem_master_bready , RTL___near_mem___dmem_master_rready , RTL___near_mem___dmem_master_wlast , RTL___near_mem___dmem_master_wvalid , RTL___near_mem___dmem_valid , RTL___near_mem___imem_exc , RTL___near_mem___imem_is_i32_not_i16 , RTL___near_mem___imem_master_arlock , RTL___near_mem___imem_master_arvalid , RTL___near_mem___imem_master_awlock , RTL___near_mem___imem_master_awvalid , RTL___near_mem___imem_master_bready , RTL___near_mem___imem_master_rready , RTL___near_mem___imem_master_wlast , RTL___near_mem___imem_master_wvalid , RTL___near_mem___imem_valid ; reg[3:0] RTL___near_mem___cfg_verbosity ; 
    wire[3:0] RTL___near_mem___cfg_verbosity$D_IN ; 
    wire RTL___near_mem___cfg_verbosity$EN ; reg[1:0] RTL___near_mem___rg_state ; reg[1:0] RTL___near_mem___rg_state$D_IN ; 
    wire RTL___near_mem___rg_state$EN ; 
    wire[63:0] RTL___near_mem___dcache$mem_master_araddr , RTL___near_mem___dcache$mem_master_awaddr , RTL___near_mem___dcache$mem_master_rdata , RTL___near_mem___dcache$mem_master_wdata , RTL___near_mem___dcache$req_st_value , RTL___near_mem___dcache$word64 ; 
    wire[31:0] RTL___near_mem___dcache$req_addr , RTL___near_mem___dcache$req_satp ; 
    wire[7:0] RTL___near_mem___dcache$mem_master_arlen , RTL___near_mem___dcache$mem_master_awlen , RTL___near_mem___dcache$mem_master_wstrb ; 
    wire[3:0] RTL___near_mem___dcache$exc_code , RTL___near_mem___dcache$mem_master_arcache , RTL___near_mem___dcache$mem_master_arid , RTL___near_mem___dcache$mem_master_arqos , RTL___near_mem___dcache$mem_master_arregion , RTL___near_mem___dcache$mem_master_awcache , RTL___near_mem___dcache$mem_master_awid , RTL___near_mem___dcache$mem_master_awqos , RTL___near_mem___dcache$mem_master_awregion , RTL___near_mem___dcache$mem_master_bid , RTL___near_mem___dcache$mem_master_rid , RTL___near_mem___dcache$set_verbosity_verbosity ; 
    wire[2:0] RTL___near_mem___dcache$mem_master_arprot , RTL___near_mem___dcache$mem_master_arsize , RTL___near_mem___dcache$mem_master_awprot , RTL___near_mem___dcache$mem_master_awsize , RTL___near_mem___dcache$req_f3 ; 
    wire[1:0] RTL___near_mem___dcache$mem_master_arburst , RTL___near_mem___dcache$mem_master_awburst , RTL___near_mem___dcache$mem_master_bresp , RTL___near_mem___dcache$mem_master_rresp , RTL___near_mem___dcache$req_priv ; 
    wire RTL___near_mem___dcache$EN_req , RTL___near_mem___dcache$EN_server_flush_request_put , RTL___near_mem___dcache$EN_server_flush_response_get , RTL___near_mem___dcache$EN_server_reset_request_put , RTL___near_mem___dcache$EN_server_reset_response_get , RTL___near_mem___dcache$EN_set_verbosity , RTL___near_mem___dcache$EN_tlb_flush , RTL___near_mem___dcache$RDY_server_flush_request_put , RTL___near_mem___dcache$RDY_server_flush_response_get , RTL___near_mem___dcache$RDY_server_reset_request_put , RTL___near_mem___dcache$RDY_server_reset_response_get , RTL___near_mem___dcache$exc , RTL___near_mem___dcache$mem_master_arlock , RTL___near_mem___dcache$mem_master_arready , RTL___near_mem___dcache$mem_master_arvalid , RTL___near_mem___dcache$mem_master_awlock , RTL___near_mem___dcache$mem_master_awready , RTL___near_mem___dcache$mem_master_awvalid , RTL___near_mem___dcache$mem_master_bready , RTL___near_mem___dcache$mem_master_bvalid , RTL___near_mem___dcache$mem_master_rlast , RTL___near_mem___dcache$mem_master_rready , RTL___near_mem___dcache$mem_master_rvalid , RTL___near_mem___dcache$mem_master_wlast , RTL___near_mem___dcache$mem_master_wready , RTL___near_mem___dcache$mem_master_wvalid , RTL___near_mem___dcache$req_mstatus_MXR , RTL___near_mem___dcache$req_op , RTL___near_mem___dcache$req_sstatus_SUM , RTL___near_mem___dcache$valid ; 
    wire RTL___near_mem___f_reset_rsps$CLR , RTL___near_mem___f_reset_rsps$DEQ , RTL___near_mem___f_reset_rsps$EMPTY_N , RTL___near_mem___f_reset_rsps$ENQ , RTL___near_mem___f_reset_rsps$FULL_N ; 
    wire[63:0] RTL___near_mem___icache$mem_master_araddr , RTL___near_mem___icache$mem_master_awaddr , RTL___near_mem___icache$mem_master_rdata , RTL___near_mem___icache$mem_master_wdata , RTL___near_mem___icache$req_st_value , RTL___near_mem___icache$word64 ; 
    wire[31:0] RTL___near_mem___icache$addr , RTL___near_mem___icache$req_addr , RTL___near_mem___icache$req_satp ; 
    wire[7:0] RTL___near_mem___icache$mem_master_arlen , RTL___near_mem___icache$mem_master_awlen , RTL___near_mem___icache$mem_master_wstrb ; 
    wire[3:0] RTL___near_mem___icache$exc_code , RTL___near_mem___icache$mem_master_arcache , RTL___near_mem___icache$mem_master_arid , RTL___near_mem___icache$mem_master_arqos , RTL___near_mem___icache$mem_master_arregion , RTL___near_mem___icache$mem_master_awcache , RTL___near_mem___icache$mem_master_awid , RTL___near_mem___icache$mem_master_awqos , RTL___near_mem___icache$mem_master_awregion , RTL___near_mem___icache$mem_master_bid , RTL___near_mem___icache$mem_master_rid , RTL___near_mem___icache$set_verbosity_verbosity ; 
    wire[2:0] RTL___near_mem___icache$mem_master_arprot , RTL___near_mem___icache$mem_master_arsize , RTL___near_mem___icache$mem_master_awprot , RTL___near_mem___icache$mem_master_awsize , RTL___near_mem___icache$req_f3 ; 
    wire[1:0] RTL___near_mem___icache$mem_master_arburst , RTL___near_mem___icache$mem_master_awburst , RTL___near_mem___icache$mem_master_bresp , RTL___near_mem___icache$mem_master_rresp , RTL___near_mem___icache$req_priv ; 
    wire RTL___near_mem___icache$EN_req , RTL___near_mem___icache$EN_server_flush_request_put , RTL___near_mem___icache$EN_server_flush_response_get , RTL___near_mem___icache$EN_server_reset_request_put , RTL___near_mem___icache$EN_server_reset_response_get , RTL___near_mem___icache$EN_set_verbosity , RTL___near_mem___icache$EN_tlb_flush , RTL___near_mem___icache$RDY_server_flush_request_put , RTL___near_mem___icache$RDY_server_flush_response_get , RTL___near_mem___icache$RDY_server_reset_request_put , RTL___near_mem___icache$RDY_server_reset_response_get , RTL___near_mem___icache$exc , RTL___near_mem___icache$mem_master_arlock , RTL___near_mem___icache$mem_master_arready , RTL___near_mem___icache$mem_master_arvalid , RTL___near_mem___icache$mem_master_awlock , RTL___near_mem___icache$mem_master_awready , RTL___near_mem___icache$mem_master_awvalid , RTL___near_mem___icache$mem_master_bready , RTL___near_mem___icache$mem_master_bvalid , RTL___near_mem___icache$mem_master_rlast , RTL___near_mem___icache$mem_master_rready , RTL___near_mem___icache$mem_master_rvalid , RTL___near_mem___icache$mem_master_wlast , RTL___near_mem___icache$mem_master_wready , RTL___near_mem___icache$mem_master_wvalid , RTL___near_mem___icache$req_mstatus_MXR , RTL___near_mem___icache$req_op , RTL___near_mem___icache$req_sstatus_SUM , RTL___near_mem___icache$valid ; 
    wire[63:0] RTL___near_mem___soc_map$m_is_IO_addr_addr , RTL___near_mem___soc_map$m_is_mem_addr_addr , RTL___near_mem___soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL___near_mem___CAN_FIRE_RL_rl_reset , RTL___near_mem___CAN_FIRE_RL_rl_reset_complete , RTL___near_mem___CAN_FIRE_dmem_master_m_arready , RTL___near_mem___CAN_FIRE_dmem_master_m_awready , RTL___near_mem___CAN_FIRE_dmem_master_m_bvalid , RTL___near_mem___CAN_FIRE_dmem_master_m_rvalid , RTL___near_mem___CAN_FIRE_dmem_master_m_wready , RTL___near_mem___CAN_FIRE_dmem_req , RTL___near_mem___CAN_FIRE_imem_master_m_arready , RTL___near_mem___CAN_FIRE_imem_master_m_awready , RTL___near_mem___CAN_FIRE_imem_master_m_bvalid , RTL___near_mem___CAN_FIRE_imem_master_m_rvalid , RTL___near_mem___CAN_FIRE_imem_master_m_wready , RTL___near_mem___CAN_FIRE_imem_req , RTL___near_mem___CAN_FIRE_server_fence_i_request_put , RTL___near_mem___CAN_FIRE_server_fence_i_response_get , RTL___near_mem___CAN_FIRE_server_fence_request_put , RTL___near_mem___CAN_FIRE_server_fence_response_get , RTL___near_mem___CAN_FIRE_server_reset_request_put , RTL___near_mem___CAN_FIRE_server_reset_response_get , RTL___near_mem___CAN_FIRE_sfence_vma , RTL___near_mem___WILL_FIRE_RL_rl_reset , RTL___near_mem___WILL_FIRE_RL_rl_reset_complete , RTL___near_mem___WILL_FIRE_dmem_master_m_arready , RTL___near_mem___WILL_FIRE_dmem_master_m_awready , RTL___near_mem___WILL_FIRE_dmem_master_m_bvalid , RTL___near_mem___WILL_FIRE_dmem_master_m_rvalid , RTL___near_mem___WILL_FIRE_dmem_master_m_wready , RTL___near_mem___WILL_FIRE_dmem_req , RTL___near_mem___WILL_FIRE_imem_master_m_arready , RTL___near_mem___WILL_FIRE_imem_master_m_awready , RTL___near_mem___WILL_FIRE_imem_master_m_bvalid , RTL___near_mem___WILL_FIRE_imem_master_m_rvalid , RTL___near_mem___WILL_FIRE_imem_master_m_wready , RTL___near_mem___WILL_FIRE_imem_req , RTL___near_mem___WILL_FIRE_server_fence_i_request_put , RTL___near_mem___WILL_FIRE_server_fence_i_response_get , RTL___near_mem___WILL_FIRE_server_fence_request_put , RTL___near_mem___WILL_FIRE_server_fence_response_get , RTL___near_mem___WILL_FIRE_server_reset_request_put , RTL___near_mem___WILL_FIRE_server_reset_response_get , RTL___near_mem___WILL_FIRE_sfence_vma ; 
    wire RTL___near_mem___MUX_rg_state$write_1__SEL_2 , RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; reg[31:0] RTL___near_mem___v__h1643 ; reg[31:0] RTL___near_mem___v__h1794 ; reg[31:0] RTL___near_mem___v__h1637 ; reg[31:0] RTL___near_mem___v__h1788 ; 
    wire RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 ; 
  assign  RTL___near_mem___RDY_server_reset_request_put = RTL___near_mem___rg_state ==2'd2; 
  assign  RTL___near_mem___CAN_FIRE_server_reset_request_put = RTL___near_mem___rg_state ==2'd2; 
  assign  RTL___near_mem___WILL_FIRE_server_reset_request_put = RTL___near_mem___EN_server_reset_request_put ; 
  assign  RTL___near_mem___RDY_server_reset_response_get = RTL___near_mem___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___CAN_FIRE_server_reset_response_get = RTL___near_mem___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___WILL_FIRE_server_reset_response_get = RTL___near_mem___EN_server_reset_response_get ; 
  assign  RTL___near_mem___CAN_FIRE_imem_req =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_req = RTL___near_mem___EN_imem_req ; 
  assign  RTL___near_mem___imem_valid = RTL___near_mem___icache$valid ; 
  assign  RTL___near_mem___imem_is_i32_not_i16 =1'd1; 
  assign  RTL___near_mem___imem_pc = RTL___near_mem___icache$addr ; 
  assign  RTL___near_mem___imem_instr = RTL___near_mem___icache$word64 [31:0]; 
  assign  RTL___near_mem___imem_exc = RTL___near_mem___icache$exc ; 
  assign  RTL___near_mem___imem_exc_code = RTL___near_mem___icache$exc_code ; 
  assign  RTL___near_mem___imem_tval = RTL___near_mem___icache$addr ; 
  assign  RTL___near_mem___imem_master_awvalid = RTL___near_mem___icache$mem_master_awvalid ; 
  assign  RTL___near_mem___imem_master_awid = RTL___near_mem___icache$mem_master_awid ; 
  assign  RTL___near_mem___imem_master_awaddr = RTL___near_mem___icache$mem_master_awaddr ; 
  assign  RTL___near_mem___imem_master_awlen = RTL___near_mem___icache$mem_master_awlen ; 
  assign  RTL___near_mem___imem_master_awsize = RTL___near_mem___icache$mem_master_awsize ; 
  assign  RTL___near_mem___imem_master_awburst = RTL___near_mem___icache$mem_master_awburst ; 
  assign  RTL___near_mem___imem_master_awlock = RTL___near_mem___icache$mem_master_awlock ; 
  assign  RTL___near_mem___imem_master_awcache = RTL___near_mem___icache$mem_master_awcache ; 
  assign  RTL___near_mem___imem_master_awprot = RTL___near_mem___icache$mem_master_awprot ; 
  assign  RTL___near_mem___imem_master_awqos = RTL___near_mem___icache$mem_master_awqos ; 
  assign  RTL___near_mem___imem_master_awregion = RTL___near_mem___icache$mem_master_awregion ; 
  assign  RTL___near_mem___CAN_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_master_m_awready =1'd1; 
  assign  RTL___near_mem___imem_master_wvalid = RTL___near_mem___icache$mem_master_wvalid ; 
  assign  RTL___near_mem___imem_master_wdata = RTL___near_mem___icache$mem_master_wdata ; 
  assign  RTL___near_mem___imem_master_wstrb = RTL___near_mem___icache$mem_master_wstrb ; 
  assign  RTL___near_mem___imem_master_wlast = RTL___near_mem___icache$mem_master_wlast ; 
  assign  RTL___near_mem___CAN_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_master_m_wready =1'd1; 
  assign  RTL___near_mem___CAN_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___imem_master_bready = RTL___near_mem___icache$mem_master_bready ; 
  assign  RTL___near_mem___imem_master_arvalid = RTL___near_mem___icache$mem_master_arvalid ; 
  assign  RTL___near_mem___imem_master_arid = RTL___near_mem___icache$mem_master_arid ; 
  assign  RTL___near_mem___imem_master_araddr = RTL___near_mem___icache$mem_master_araddr ; 
  assign  RTL___near_mem___imem_master_arlen = RTL___near_mem___icache$mem_master_arlen ; 
  assign  RTL___near_mem___imem_master_arsize = RTL___near_mem___icache$mem_master_arsize ; 
  assign  RTL___near_mem___imem_master_arburst = RTL___near_mem___icache$mem_master_arburst ; 
  assign  RTL___near_mem___imem_master_arlock = RTL___near_mem___icache$mem_master_arlock ; 
  assign  RTL___near_mem___imem_master_arcache = RTL___near_mem___icache$mem_master_arcache ; 
  assign  RTL___near_mem___imem_master_arprot = RTL___near_mem___icache$mem_master_arprot ; 
  assign  RTL___near_mem___imem_master_arqos = RTL___near_mem___icache$mem_master_arqos ; 
  assign  RTL___near_mem___imem_master_arregion = RTL___near_mem___icache$mem_master_arregion ; 
  assign  RTL___near_mem___CAN_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_master_m_arready =1'd1; 
  assign  RTL___near_mem___CAN_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_imem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___imem_master_rready = RTL___near_mem___icache$mem_master_rready ; 
  assign  RTL___near_mem___CAN_FIRE_dmem_req =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_req = RTL___near_mem___EN_dmem_req ; 
  assign  RTL___near_mem___dmem_valid = RTL___near_mem___dcache$valid ; 
  assign  RTL___near_mem___dmem_word64 = RTL___near_mem___dcache$word64 ; 
  assign  RTL___near_mem___dmem_st_amo_val =64'hAAAAAAAAAAAAAAAA; 
  assign  RTL___near_mem___dmem_exc = RTL___near_mem___dcache$exc ; 
  assign  RTL___near_mem___dmem_exc_code = RTL___near_mem___dcache$exc_code ; 
  assign  RTL___near_mem___dmem_master_awvalid = RTL___near_mem___dcache$mem_master_awvalid ; 
  assign  RTL___near_mem___dmem_master_awid = RTL___near_mem___dcache$mem_master_awid ; 
  assign  RTL___near_mem___dmem_master_awaddr = RTL___near_mem___dcache$mem_master_awaddr ; 
  assign  RTL___near_mem___dmem_master_awlen = RTL___near_mem___dcache$mem_master_awlen ; 
  assign  RTL___near_mem___dmem_master_awsize = RTL___near_mem___dcache$mem_master_awsize ; 
  assign  RTL___near_mem___dmem_master_awburst = RTL___near_mem___dcache$mem_master_awburst ; 
  assign  RTL___near_mem___dmem_master_awlock = RTL___near_mem___dcache$mem_master_awlock ; 
  assign  RTL___near_mem___dmem_master_awcache = RTL___near_mem___dcache$mem_master_awcache ; 
  assign  RTL___near_mem___dmem_master_awprot = RTL___near_mem___dcache$mem_master_awprot ; 
  assign  RTL___near_mem___dmem_master_awqos = RTL___near_mem___dcache$mem_master_awqos ; 
  assign  RTL___near_mem___dmem_master_awregion = RTL___near_mem___dcache$mem_master_awregion ; 
  assign  RTL___near_mem___CAN_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_master_m_awready =1'd1; 
  assign  RTL___near_mem___dmem_master_wvalid = RTL___near_mem___dcache$mem_master_wvalid ; 
  assign  RTL___near_mem___dmem_master_wdata = RTL___near_mem___dcache$mem_master_wdata ; 
  assign  RTL___near_mem___dmem_master_wstrb = RTL___near_mem___dcache$mem_master_wstrb ; 
  assign  RTL___near_mem___dmem_master_wlast = RTL___near_mem___dcache$mem_master_wlast ; 
  assign  RTL___near_mem___CAN_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_master_m_wready =1'd1; 
  assign  RTL___near_mem___CAN_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___dmem_master_bready = RTL___near_mem___dcache$mem_master_bready ; 
  assign  RTL___near_mem___dmem_master_arvalid = RTL___near_mem___dcache$mem_master_arvalid ; 
  assign  RTL___near_mem___dmem_master_arid = RTL___near_mem___dcache$mem_master_arid ; 
  assign  RTL___near_mem___dmem_master_araddr = RTL___near_mem___dcache$mem_master_araddr ; 
  assign  RTL___near_mem___dmem_master_arlen = RTL___near_mem___dcache$mem_master_arlen ; 
  assign  RTL___near_mem___dmem_master_arsize = RTL___near_mem___dcache$mem_master_arsize ; 
  assign  RTL___near_mem___dmem_master_arburst = RTL___near_mem___dcache$mem_master_arburst ; 
  assign  RTL___near_mem___dmem_master_arlock = RTL___near_mem___dcache$mem_master_arlock ; 
  assign  RTL___near_mem___dmem_master_arcache = RTL___near_mem___dcache$mem_master_arcache ; 
  assign  RTL___near_mem___dmem_master_arprot = RTL___near_mem___dcache$mem_master_arprot ; 
  assign  RTL___near_mem___dmem_master_arqos = RTL___near_mem___dcache$mem_master_arqos ; 
  assign  RTL___near_mem___dmem_master_arregion = RTL___near_mem___dcache$mem_master_arregion ; 
  assign  RTL___near_mem___CAN_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_master_m_arready =1'd1; 
  assign  RTL___near_mem___CAN_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_dmem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___dmem_master_rready = RTL___near_mem___dcache$mem_master_rready ; 
  assign  RTL___near_mem___RDY_server_fence_i_request_put = RTL___near_mem___dcache$RDY_server_flush_request_put && RTL___near_mem___icache$RDY_server_flush_request_put ; 
  assign  RTL___near_mem___CAN_FIRE_server_fence_i_request_put = RTL___near_mem___dcache$RDY_server_flush_request_put && RTL___near_mem___icache$RDY_server_flush_request_put ; 
  assign  RTL___near_mem___WILL_FIRE_server_fence_i_request_put = RTL___near_mem___EN_server_fence_i_request_put ; 
  assign  RTL___near_mem___RDY_server_fence_i_response_get = RTL___near_mem___dcache$RDY_server_flush_response_get && RTL___near_mem___icache$RDY_server_flush_response_get ; 
  assign  RTL___near_mem___CAN_FIRE_server_fence_i_response_get = RTL___near_mem___dcache$RDY_server_flush_response_get && RTL___near_mem___icache$RDY_server_flush_response_get ; 
  assign  RTL___near_mem___WILL_FIRE_server_fence_i_response_get = RTL___near_mem___EN_server_fence_i_response_get ; 
  assign  RTL___near_mem___RDY_server_fence_request_put = RTL___near_mem___dcache$RDY_server_flush_request_put ; 
  assign  RTL___near_mem___CAN_FIRE_server_fence_request_put = RTL___near_mem___dcache$RDY_server_flush_request_put ; 
  assign  RTL___near_mem___WILL_FIRE_server_fence_request_put = RTL___near_mem___EN_server_fence_request_put ; 
  assign  RTL___near_mem___RDY_server_fence_response_get = RTL___near_mem___dcache$RDY_server_flush_response_get ; 
  assign  RTL___near_mem___CAN_FIRE_server_fence_response_get = RTL___near_mem___dcache$RDY_server_flush_response_get ; 
  assign  RTL___near_mem___WILL_FIRE_server_fence_response_get = RTL___near_mem___EN_server_fence_response_get ; 
  assign  RTL___near_mem___RDY_sfence_vma =1'd1; 
  assign  RTL___near_mem___CAN_FIRE_sfence_vma =1'd1; 
  assign  RTL___near_mem___WILL_FIRE_sfence_vma = RTL___near_mem___EN_sfence_vma ;  
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL___near_mem___dcache___CLK;
    wire RTL___near_mem___dcache___RST_N;
    wire[3:0] RTL___near_mem___dcache___set_verbosity_verbosity;
    wire RTL___near_mem___dcache___EN_set_verbosity;
    wire RTL___near_mem___dcache___EN_server_reset_request_put;
    wire RTL___near_mem___dcache___EN_server_reset_response_get;
    wire RTL___near_mem___dcache___req_op;
    wire[2:0] RTL___near_mem___dcache___req_f3;
    wire[31:0] RTL___near_mem___dcache___req_addr;
    wire[63:0] RTL___near_mem___dcache___req_st_value;
    wire[1:0] RTL___near_mem___dcache___req_priv;
    wire RTL___near_mem___dcache___req_sstatus_SUM;
    wire RTL___near_mem___dcache___req_mstatus_MXR;
    wire[31:0] RTL___near_mem___dcache___req_satp;
    wire RTL___near_mem___dcache___EN_req;
    wire RTL___near_mem___dcache___EN_server_flush_request_put;
    wire RTL___near_mem___dcache___EN_server_flush_response_get;
    wire RTL___near_mem___dcache___EN_tlb_flush;
    wire RTL___near_mem___dcache___mem_master_awready;
    wire RTL___near_mem___dcache___mem_master_wready;
    wire RTL___near_mem___dcache___mem_master_bvalid;
    wire[3:0] RTL___near_mem___dcache___mem_master_bid;
    wire[1:0] RTL___near_mem___dcache___mem_master_bresp;
    wire RTL___near_mem___dcache___mem_master_arready;
    wire RTL___near_mem___dcache___mem_master_rvalid;
    wire[3:0] RTL___near_mem___dcache___mem_master_rid;
    wire[63:0] RTL___near_mem___dcache___mem_master_rdata;
    wire[1:0] RTL___near_mem___dcache___mem_master_rresp;
    wire RTL___near_mem___dcache___mem_master_rlast;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire[31:0] RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire[31:0] RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    wire RTL___near_mem___icache___CLK;
    wire RTL___near_mem___icache___RST_N;
    wire[3:0] RTL___near_mem___icache___set_verbosity_verbosity;
    wire RTL___near_mem___icache___EN_set_verbosity;
    wire RTL___near_mem___icache___EN_server_reset_request_put;
    wire RTL___near_mem___icache___EN_server_reset_response_get;
    wire RTL___near_mem___icache___req_op;
    wire[2:0] RTL___near_mem___icache___req_f3;
    wire[31:0] RTL___near_mem___icache___req_addr;
    wire[63:0] RTL___near_mem___icache___req_st_value;
    wire[1:0] RTL___near_mem___icache___req_priv;
    wire RTL___near_mem___icache___req_sstatus_SUM;
    wire RTL___near_mem___icache___req_mstatus_MXR;
    wire[31:0] RTL___near_mem___icache___req_satp;
    wire RTL___near_mem___icache___EN_req;
    wire RTL___near_mem___icache___EN_server_flush_request_put;
    wire RTL___near_mem___icache___EN_server_flush_response_get;
    wire RTL___near_mem___icache___EN_tlb_flush;
    wire RTL___near_mem___icache___mem_master_awready;
    wire RTL___near_mem___icache___mem_master_wready;
    wire RTL___near_mem___icache___mem_master_bvalid;
    wire[3:0] RTL___near_mem___icache___mem_master_bid;
    wire[1:0] RTL___near_mem___icache___mem_master_bresp;
    wire RTL___near_mem___icache___mem_master_arready;
    wire RTL___near_mem___icache___mem_master_rvalid;
    wire[3:0] RTL___near_mem___icache___mem_master_rid;
    wire[63:0] RTL___near_mem___icache___mem_master_rdata;
    wire[1:0] RTL___near_mem___icache___mem_master_rresp;
    wire RTL___near_mem___icache___mem_master_rlast;

    reg[63:0] RTL___near_mem___dcache___word64 ; 
    wire[63:0] RTL___near_mem___dcache___mem_master_araddr , RTL___near_mem___dcache___mem_master_awaddr , RTL___near_mem___dcache___mem_master_wdata , RTL___near_mem___dcache___st_amo_val ; 
    wire[31:0] RTL___near_mem___dcache___addr ; 
    wire[7:0] RTL___near_mem___dcache___mem_master_arlen , RTL___near_mem___dcache___mem_master_awlen , RTL___near_mem___dcache___mem_master_wstrb ; 
    wire[3:0] RTL___near_mem___dcache___exc_code , RTL___near_mem___dcache___mem_master_arcache , RTL___near_mem___dcache___mem_master_arid , RTL___near_mem___dcache___mem_master_arqos , RTL___near_mem___dcache___mem_master_arregion , RTL___near_mem___dcache___mem_master_awcache , RTL___near_mem___dcache___mem_master_awid , RTL___near_mem___dcache___mem_master_awqos , RTL___near_mem___dcache___mem_master_awregion ; 
    wire[2:0] RTL___near_mem___dcache___mem_master_arprot , RTL___near_mem___dcache___mem_master_arsize , RTL___near_mem___dcache___mem_master_awprot , RTL___near_mem___dcache___mem_master_awsize ; 
    wire[1:0] RTL___near_mem___dcache___mem_master_arburst , RTL___near_mem___dcache___mem_master_awburst ; 
    wire RTL___near_mem___dcache___RDY_server_flush_request_put , RTL___near_mem___dcache___RDY_server_flush_response_get , RTL___near_mem___dcache___RDY_server_reset_request_put , RTL___near_mem___dcache___RDY_server_reset_response_get , RTL___near_mem___dcache___RDY_set_verbosity , RTL___near_mem___dcache___RDY_tlb_flush , RTL___near_mem___dcache___exc , RTL___near_mem___dcache___mem_master_arlock , RTL___near_mem___dcache___mem_master_arvalid , RTL___near_mem___dcache___mem_master_awlock , RTL___near_mem___dcache___mem_master_awvalid , RTL___near_mem___dcache___mem_master_bready , RTL___near_mem___dcache___mem_master_rready , RTL___near_mem___dcache___mem_master_wlast , RTL___near_mem___dcache___mem_master_wvalid , RTL___near_mem___dcache___valid ; 
    wire[3:0] RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port0__write_1 , RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port1__write_1 , RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port2__read , RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port3__read ; 
    wire RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN_port2__write , RTL___near_mem___dcache___dw_valid$whas ; reg[3:0] RTL___near_mem___dcache___cfg_verbosity ; 
    wire[3:0] RTL___near_mem___dcache___cfg_verbosity$D_IN ; 
    wire RTL___near_mem___dcache___cfg_verbosity$EN ; reg[3:0] RTL___near_mem___dcache___ctr_wr_rsps_pending_crg ; 
    wire[3:0] RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$D_IN ; 
    wire RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN ; reg[31:0] RTL___near_mem___dcache___rg_addr ; 
    wire[31:0] RTL___near_mem___dcache___rg_addr$D_IN ; 
    wire RTL___near_mem___dcache___rg_addr$EN ; reg[6:0] RTL___near_mem___dcache___rg_cset_in_cache ; 
    wire[6:0] RTL___near_mem___dcache___rg_cset_in_cache$D_IN ; 
    wire RTL___near_mem___dcache___rg_cset_in_cache$EN ; 
    reg RTL___near_mem___dcache___rg_error_during_refill ; 
    wire RTL___near_mem___dcache___rg_error_during_refill$D_IN , RTL___near_mem___dcache___rg_error_during_refill$EN ; reg[3:0] RTL___near_mem___dcache___rg_exc_code ; reg[3:0] RTL___near_mem___dcache___rg_exc_code$D_IN ; 
    wire RTL___near_mem___dcache___rg_exc_code$EN ; reg[2:0] RTL___near_mem___dcache___rg_f3 ; 
    wire[2:0] RTL___near_mem___dcache___rg_f3$D_IN ; 
    wire RTL___near_mem___dcache___rg_f3$EN ; reg[63:0] RTL___near_mem___dcache___rg_ld_val ; 
    wire[63:0] RTL___near_mem___dcache___rg_ld_val$D_IN ; 
    wire RTL___near_mem___dcache___rg_ld_val$EN ; reg[31:0] RTL___near_mem___dcache___rg_lower_word32 ; 
    wire[31:0] RTL___near_mem___dcache___rg_lower_word32$D_IN ; 
    wire RTL___near_mem___dcache___rg_lower_word32$EN ; 
    reg RTL___near_mem___dcache___rg_lower_word32_full ; 
    wire RTL___near_mem___dcache___rg_lower_word32_full$D_IN , RTL___near_mem___dcache___rg_lower_word32_full$EN ; 
    reg RTL___near_mem___dcache___rg_op ; 
    wire RTL___near_mem___dcache___rg_op$D_IN , RTL___near_mem___dcache___rg_op$EN ; reg[31:0] RTL___near_mem___dcache___rg_pa ; 
    wire[31:0] RTL___near_mem___dcache___rg_pa$D_IN ; 
    wire RTL___near_mem___dcache___rg_pa$EN ; reg[31:0] RTL___near_mem___dcache___rg_pte_pa ; 
    wire[31:0] RTL___near_mem___dcache___rg_pte_pa$D_IN ; 
    wire RTL___near_mem___dcache___rg_pte_pa$EN ; reg[63:0] RTL___near_mem___dcache___rg_st_amo_val ; 
    wire[63:0] RTL___near_mem___dcache___rg_st_amo_val$D_IN ; 
    wire RTL___near_mem___dcache___rg_st_amo_val$EN ; reg[3:0] RTL___near_mem___dcache___rg_state ; reg[3:0] RTL___near_mem___dcache___rg_state$D_IN ; 
    wire RTL___near_mem___dcache___rg_state$EN ; reg[8:0] RTL___near_mem___dcache___rg_word64_set_in_cache ; 
    wire[8:0] RTL___near_mem___dcache___rg_word64_set_in_cache$D_IN ; 
    wire RTL___near_mem___dcache___rg_word64_set_in_cache$EN ; 
    wire[98:0] RTL___near_mem___dcache___f_fabric_write_reqs$D_IN , RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT ; 
    wire RTL___near_mem___dcache___f_fabric_write_reqs$CLR , RTL___near_mem___dcache___f_fabric_write_reqs$DEQ , RTL___near_mem___dcache___f_fabric_write_reqs$EMPTY_N , RTL___near_mem___dcache___f_fabric_write_reqs$ENQ , RTL___near_mem___dcache___f_fabric_write_reqs$FULL_N ; 
    wire RTL___near_mem___dcache___f_reset_reqs$CLR , RTL___near_mem___dcache___f_reset_reqs$DEQ , RTL___near_mem___dcache___f_reset_reqs$D_IN , RTL___near_mem___dcache___f_reset_reqs$D_OUT , RTL___near_mem___dcache___f_reset_reqs$EMPTY_N , RTL___near_mem___dcache___f_reset_reqs$ENQ , RTL___near_mem___dcache___f_reset_reqs$FULL_N ; 
    wire RTL___near_mem___dcache___f_reset_rsps$CLR , RTL___near_mem___dcache___f_reset_rsps$DEQ , RTL___near_mem___dcache___f_reset_rsps$D_IN , RTL___near_mem___dcache___f_reset_rsps$D_OUT , RTL___near_mem___dcache___f_reset_rsps$EMPTY_N , RTL___near_mem___dcache___f_reset_rsps$ENQ , RTL___near_mem___dcache___f_reset_rsps$FULL_N ; 
    wire[96:0] RTL___near_mem___dcache___master_xactor_f_rd_addr$D_IN , RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr$CLR , RTL___near_mem___dcache___master_xactor_f_rd_addr$DEQ , RTL___near_mem___dcache___master_xactor_f_rd_addr$EMPTY_N , RTL___near_mem___dcache___master_xactor_f_rd_addr$ENQ , RTL___near_mem___dcache___master_xactor_f_rd_addr$FULL_N ; 
    wire[70:0] RTL___near_mem___dcache___master_xactor_f_rd_data$D_IN , RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_data$CLR , RTL___near_mem___dcache___master_xactor_f_rd_data$DEQ , RTL___near_mem___dcache___master_xactor_f_rd_data$EMPTY_N , RTL___near_mem___dcache___master_xactor_f_rd_data$ENQ , RTL___near_mem___dcache___master_xactor_f_rd_data$FULL_N ; 
    wire[96:0] RTL___near_mem___dcache___master_xactor_f_wr_addr$D_IN , RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr$CLR , RTL___near_mem___dcache___master_xactor_f_wr_addr$DEQ , RTL___near_mem___dcache___master_xactor_f_wr_addr$EMPTY_N , RTL___near_mem___dcache___master_xactor_f_wr_addr$ENQ , RTL___near_mem___dcache___master_xactor_f_wr_addr$FULL_N ; 
    wire[72:0] RTL___near_mem___dcache___master_xactor_f_wr_data$D_IN , RTL___near_mem___dcache___master_xactor_f_wr_data$D_OUT ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_data$CLR , RTL___near_mem___dcache___master_xactor_f_wr_data$DEQ , RTL___near_mem___dcache___master_xactor_f_wr_data$EMPTY_N , RTL___near_mem___dcache___master_xactor_f_wr_data$ENQ , RTL___near_mem___dcache___master_xactor_f_wr_data$FULL_N ; 
    wire[5:0] RTL___near_mem___dcache___master_xactor_f_wr_resp$D_IN , RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp$CLR , RTL___near_mem___dcache___master_xactor_f_wr_resp$DEQ , RTL___near_mem___dcache___master_xactor_f_wr_resp$EMPTY_N , RTL___near_mem___dcache___master_xactor_f_wr_resp$ENQ , RTL___near_mem___dcache___master_xactor_f_wr_resp$FULL_N ; 
    wire[22:0] RTL___near_mem___dcache___ram_state_and_ctag_cset$DIA , RTL___near_mem___dcache___ram_state_and_ctag_cset$DIB , RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB ; 
    wire[6:0] RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRA , RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRB ; 
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset$ENA , RTL___near_mem___dcache___ram_state_and_ctag_cset$ENB , RTL___near_mem___dcache___ram_state_and_ctag_cset$WEA , RTL___near_mem___dcache___ram_state_and_ctag_cset$WEB ; reg[63:0] RTL___near_mem___dcache___ram_word64_set$DIB ; reg[8:0] RTL___near_mem___dcache___ram_word64_set$ADDRB ; 
    wire[63:0] RTL___near_mem___dcache___ram_word64_set$DIA , RTL___near_mem___dcache___ram_word64_set$DOB ; 
    wire[8:0] RTL___near_mem___dcache___ram_word64_set$ADDRA ; 
    wire RTL___near_mem___dcache___ram_word64_set$ENA , RTL___near_mem___dcache___ram_word64_set$ENB , RTL___near_mem___dcache___ram_word64_set$WEA , RTL___near_mem___dcache___ram_word64_set$WEB ; 
    wire[63:0] RTL___near_mem___dcache___soc_map$m_is_IO_addr_addr , RTL___near_mem___dcache___soc_map$m_is_mem_addr_addr , RTL___near_mem___dcache___soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL___near_mem___dcache___soc_map$m_is_mem_addr ; 
    wire RTL___near_mem___dcache___CAN_FIRE_RL_rl_ST_AMO_response , RTL___near_mem___dcache___CAN_FIRE_RL_rl_cache_refill_rsps_loop , RTL___near_mem___dcache___CAN_FIRE_RL_rl_discard_write_rsp , RTL___near_mem___dcache___CAN_FIRE_RL_rl_drive_exception_rsp , RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req , RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_req , RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_rsp , RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_write_req , RTL___near_mem___dcache___CAN_FIRE_RL_rl_maintain_io_read_rsp , RTL___near_mem___dcache___CAN_FIRE_RL_rl_probe_and_immed_rsp , RTL___near_mem___dcache___CAN_FIRE_RL_rl_rereq , RTL___near_mem___dcache___CAN_FIRE_RL_rl_reset , RTL___near_mem___dcache___CAN_FIRE_RL_rl_start_cache_refill , RTL___near_mem___dcache___CAN_FIRE_RL_rl_start_reset , RTL___near_mem___dcache___CAN_FIRE_mem_master_m_arready , RTL___near_mem___dcache___CAN_FIRE_mem_master_m_awready , RTL___near_mem___dcache___CAN_FIRE_mem_master_m_bvalid , RTL___near_mem___dcache___CAN_FIRE_mem_master_m_rvalid , RTL___near_mem___dcache___CAN_FIRE_mem_master_m_wready , RTL___near_mem___dcache___CAN_FIRE_req , RTL___near_mem___dcache___CAN_FIRE_server_flush_request_put , RTL___near_mem___dcache___CAN_FIRE_server_flush_response_get , RTL___near_mem___dcache___CAN_FIRE_server_reset_request_put , RTL___near_mem___dcache___CAN_FIRE_server_reset_response_get , RTL___near_mem___dcache___CAN_FIRE_set_verbosity , RTL___near_mem___dcache___CAN_FIRE_tlb_flush , RTL___near_mem___dcache___WILL_FIRE_RL_rl_ST_AMO_response , RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop , RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp , RTL___near_mem___dcache___WILL_FIRE_RL_rl_drive_exception_rsp , RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req , RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req , RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp , RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req , RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp , RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp , RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq , RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset , RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill , RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset , RTL___near_mem___dcache___WILL_FIRE_mem_master_m_arready , RTL___near_mem___dcache___WILL_FIRE_mem_master_m_awready , RTL___near_mem___dcache___WILL_FIRE_mem_master_m_bvalid , RTL___near_mem___dcache___WILL_FIRE_mem_master_m_rvalid , RTL___near_mem___dcache___WILL_FIRE_mem_master_m_wready , RTL___near_mem___dcache___WILL_FIRE_req , RTL___near_mem___dcache___WILL_FIRE_server_flush_request_put , RTL___near_mem___dcache___WILL_FIRE_server_flush_response_get , RTL___near_mem___dcache___WILL_FIRE_server_reset_request_put , RTL___near_mem___dcache___WILL_FIRE_server_reset_response_get , RTL___near_mem___dcache___WILL_FIRE_set_verbosity , RTL___near_mem___dcache___WILL_FIRE_tlb_flush ; reg[63:0] RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2 ; 
    wire[98:0] RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_1 , RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
    wire[96:0] RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 , RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
    wire[22:0] RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ; 
    wire[8:0] RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_2 , RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_4 ; 
    wire[6:0] RTL___near_mem___dcache___MUX_rg_cset_in_cache$write_1__VAL_1 ; 
    wire[3:0] RTL___near_mem___dcache___MUX_rg_exc_code$write_1__VAL_1 , RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_1 , RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_4 , RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_7 , RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_9 ; 
    wire RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_1 , RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_2 , RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_3 , RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__SEL_1 , RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 , RTL___near_mem___dcache___MUX_ram_word64_set$a_put_1__SEL_1 , RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2 , RTL___near_mem___dcache___MUX_rg_error_during_refill$write_1__SEL_1 , RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_1 , RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_2 , RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_10 , RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_2 , RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_3 , RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_7 , RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_9 ; reg[31:0] RTL___near_mem___dcache___v__h2948 ; reg[31:0] RTL___near_mem___dcache___v__h3848 ; reg[31:0] RTL___near_mem___dcache___v__h3949 ; reg[31:0] RTL___near_mem___dcache___v__h4098 ; reg[31:0] RTL___near_mem___dcache___v__h12540 ; reg[31:0] RTL___near_mem___dcache___v__h14531 ; reg[31:0] RTL___near_mem___dcache___v__h15336 ; reg[31:0] RTL___near_mem___dcache___v__h15578 ; reg[31:0] RTL___near_mem___dcache___v__h17191 ; reg[31:0] RTL___near_mem___dcache___v__h17485 ; reg[31:0] RTL___near_mem___dcache___v__h18585 ; reg[31:0] RTL___near_mem___dcache___v__h18692 ; reg[31:0] RTL___near_mem___dcache___v__h18797 ; reg[31:0] RTL___near_mem___dcache___v__h18877 ; reg[31:0] RTL___near_mem___dcache___v__h19505 ; reg[31:0] RTL___near_mem___dcache___v__h19466 ; reg[31:0] RTL___near_mem___dcache___v__h3483 ; reg[31:0] RTL___near_mem___dcache___v__h19852 ; reg[31:0] RTL___near_mem___dcache___v__h2942 ; reg[31:0] RTL___near_mem___dcache___v__h3477 ; reg[31:0] RTL___near_mem___dcache___v__h3842 ; reg[31:0] RTL___near_mem___dcache___v__h3943 ; reg[31:0] RTL___near_mem___dcache___v__h4092 ; reg[31:0] RTL___near_mem___dcache___v__h12534 ; reg[31:0] RTL___near_mem___dcache___v__h14525 ; reg[31:0] RTL___near_mem___dcache___v__h15330 ; reg[31:0] RTL___near_mem___dcache___v__h15572 ; reg[31:0] RTL___near_mem___dcache___v__h17185 ; reg[31:0] RTL___near_mem___dcache___v__h17479 ; reg[31:0] RTL___near_mem___dcache___v__h18579 ; reg[31:0] RTL___near_mem___dcache___v__h18686 ; reg[31:0] RTL___near_mem___dcache___v__h18791 ; reg[31:0] RTL___near_mem___dcache___v__h18871 ; reg[31:0] RTL___near_mem___dcache___v__h19460 ; reg[31:0] RTL___near_mem___dcache___v__h19499 ; reg[31:0] RTL___near_mem___dcache___v__h19846 ; reg[63:0] RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 , RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 , RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 , RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 , RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 , RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 , RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 , RTL___near_mem___dcache___ld_val__h17594 , RTL___near_mem___dcache___mem_req_wr_data_wdata__h2699 ; reg[7:0] RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700 ; reg[2:0] RTL___near_mem___dcache___value__h17372 , RTL___near_mem___dcache___x__h2520 ; 
    wire[63:0] RTL___near_mem___dcache____theResult___snd_fst__h2707 , RTL___near_mem___dcache___cline_fabric_addr__h14584 , RTL___near_mem___dcache___fabric_addr__h17243 , RTL___near_mem___dcache___mem_req_wr_addr_awaddr__h2473 , RTL___near_mem___dcache___result__h11657 , RTL___near_mem___dcache___result__h11685 , RTL___near_mem___dcache___result__h11713 , RTL___near_mem___dcache___result__h11741 , RTL___near_mem___dcache___result__h11769 , RTL___near_mem___dcache___result__h11797 , RTL___near_mem___dcache___result__h11825 , RTL___near_mem___dcache___result__h11870 , RTL___near_mem___dcache___result__h11898 , RTL___near_mem___dcache___result__h11926 , RTL___near_mem___dcache___result__h11954 , RTL___near_mem___dcache___result__h11982 , RTL___near_mem___dcache___result__h12010 , RTL___near_mem___dcache___result__h12038 , RTL___near_mem___dcache___result__h12066 , RTL___near_mem___dcache___result__h12111 , RTL___near_mem___dcache___result__h12139 , RTL___near_mem___dcache___result__h12167 , RTL___near_mem___dcache___result__h12195 , RTL___near_mem___dcache___result__h12236 , RTL___near_mem___dcache___result__h12264 , RTL___near_mem___dcache___result__h12292 , RTL___near_mem___dcache___result__h12320 , RTL___near_mem___dcache___result__h12361 , RTL___near_mem___dcache___result__h12389 , RTL___near_mem___dcache___result__h12428 , RTL___near_mem___dcache___result__h12456 , RTL___near_mem___dcache___result__h17654 , RTL___near_mem___dcache___result__h17684 , RTL___near_mem___dcache___result__h17711 , RTL___near_mem___dcache___result__h17738 , RTL___near_mem___dcache___result__h17765 , RTL___near_mem___dcache___result__h17792 , RTL___near_mem___dcache___result__h17819 , RTL___near_mem___dcache___result__h17846 , RTL___near_mem___dcache___result__h17890 , RTL___near_mem___dcache___result__h17917 , RTL___near_mem___dcache___result__h17944 , RTL___near_mem___dcache___result__h17971 , RTL___near_mem___dcache___result__h17998 , RTL___near_mem___dcache___result__h18025 , RTL___near_mem___dcache___result__h18052 , RTL___near_mem___dcache___result__h18079 , RTL___near_mem___dcache___result__h18123 , RTL___near_mem___dcache___result__h18150 , RTL___near_mem___dcache___result__h18177 , RTL___near_mem___dcache___result__h18204 , RTL___near_mem___dcache___result__h18244 , RTL___near_mem___dcache___result__h18271 , RTL___near_mem___dcache___result__h18298 , RTL___near_mem___dcache___result__h18325 , RTL___near_mem___dcache___result__h18365 , RTL___near_mem___dcache___result__h18392 , RTL___near_mem___dcache___result__h18430 , RTL___near_mem___dcache___result__h18457 , RTL___near_mem___dcache___result__h5301 , RTL___near_mem___dcache___word64__h5094 , RTL___near_mem___dcache___y__h5337 ; 
    wire[31:0] RTL___near_mem___dcache___cline_addr__h14583 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 , RTL___near_mem___dcache___word64094_BITS_31_TO_0__q17 , RTL___near_mem___dcache___word64094_BITS_63_TO_32__q24 ; 
    wire[21:0] RTL___near_mem___dcache___pa_ctag__h4952 ; 
    wire[15:0] RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 , RTL___near_mem___dcache___word64094_BITS_15_TO_0__q16 , RTL___near_mem___dcache___word64094_BITS_31_TO_16__q20 , RTL___near_mem___dcache___word64094_BITS_47_TO_32__q23 , RTL___near_mem___dcache___word64094_BITS_63_TO_48__q27 ; 
    wire[7:0] RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 , RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 , RTL___near_mem___dcache___strobe64__h2637 , RTL___near_mem___dcache___strobe64__h2639 , RTL___near_mem___dcache___strobe64__h2641 , RTL___near_mem___dcache___word64094_BITS_15_TO_8__q18 , RTL___near_mem___dcache___word64094_BITS_23_TO_16__q19 , RTL___near_mem___dcache___word64094_BITS_31_TO_24__q21 , RTL___near_mem___dcache___word64094_BITS_39_TO_32__q22 , RTL___near_mem___dcache___word64094_BITS_47_TO_40__q25 , RTL___near_mem___dcache___word64094_BITS_55_TO_48__q26 , RTL___near_mem___dcache___word64094_BITS_63_TO_56__q28 , RTL___near_mem___dcache___word64094_BITS_7_TO_0__q15 ; 
    wire[5:0] RTL___near_mem___dcache___shift_bits__h2487 ; 
    wire[3:0] RTL___near_mem___dcache___access_exc_code__h2256 , RTL___near_mem___dcache___b__h14485 ; 
    wire RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 , RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 , RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 , RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 , RTL___near_mem___dcache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 , RTL___near_mem___dcache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 , RTL___near_mem___dcache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 , RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 , RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 , RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 ; 
  assign  RTL___near_mem___dcache___RDY_set_verbosity =1'd1; 
  assign  RTL___near_mem___dcache___CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_set_verbosity = RTL___near_mem___dcache___EN_set_verbosity ; 
  assign  RTL___near_mem___dcache___RDY_server_reset_request_put = RTL___near_mem___dcache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_server_reset_request_put = RTL___near_mem___dcache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_server_reset_request_put = RTL___near_mem___dcache___EN_server_reset_request_put ; 
  assign  RTL___near_mem___dcache___RDY_server_reset_response_get =! RTL___near_mem___dcache___f_reset_rsps$D_OUT && RTL___near_mem___dcache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_server_reset_response_get =! RTL___near_mem___dcache___f_reset_rsps$D_OUT && RTL___near_mem___dcache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_server_reset_response_get = RTL___near_mem___dcache___EN_server_reset_response_get ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_req =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_req = RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___valid = RTL___near_mem___dcache___dw_valid$whas ; 
  assign  RTL___near_mem___dcache___addr = RTL___near_mem___dcache___rg_addr ; 
  always @(       RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_1                    or   RTL___near_mem___dcache___ld_val__h17594              or   RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_2             or   RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2            or   RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_3           or   RTL___near_mem___dcache___rg_ld_val  )
         begin 
             case (1'b1) 
              RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_1  : 
                  RTL___near_mem___dcache___word64  = RTL___near_mem___dcache___ld_val__h17594 ; 
              RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_2  : 
                  RTL___near_mem___dcache___word64  = RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2 ; 
              RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_3  : 
                  RTL___near_mem___dcache___word64  = RTL___near_mem___dcache___rg_ld_val ;
              default : 
                  RTL___near_mem___dcache___word64  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL___near_mem___dcache___st_amo_val = RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_2  ? 64'd0: RTL___near_mem___dcache___rg_st_amo_val ; 
  assign  RTL___near_mem___dcache___exc = RTL___near_mem___dcache___rg_state ==4'd4; 
  assign  RTL___near_mem___dcache___exc_code = RTL___near_mem___dcache___rg_exc_code ; 
  assign  RTL___near_mem___dcache___RDY_server_flush_request_put = RTL___near_mem___dcache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_server_flush_request_put = RTL___near_mem___dcache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_server_flush_request_put = RTL___near_mem___dcache___EN_server_flush_request_put ; 
  assign  RTL___near_mem___dcache___RDY_server_flush_response_get = RTL___near_mem___dcache___f_reset_rsps$D_OUT && RTL___near_mem___dcache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_server_flush_response_get = RTL___near_mem___dcache___f_reset_rsps$D_OUT && RTL___near_mem___dcache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_server_flush_response_get = RTL___near_mem___dcache___EN_server_flush_response_get ; 
  assign  RTL___near_mem___dcache___RDY_tlb_flush =1'd1; 
  assign  RTL___near_mem___dcache___CAN_FIRE_tlb_flush =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_tlb_flush = RTL___near_mem___dcache___EN_tlb_flush ; 
  assign  RTL___near_mem___dcache___mem_master_awvalid = RTL___near_mem___dcache___master_xactor_f_wr_addr$EMPTY_N ; 
  assign  RTL___near_mem___dcache___mem_master_awid = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [96:93]; 
  assign  RTL___near_mem___dcache___mem_master_awaddr = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [92:29]; 
  assign  RTL___near_mem___dcache___mem_master_awlen = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [28:21]; 
  assign  RTL___near_mem___dcache___mem_master_awsize = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [20:18]; 
  assign  RTL___near_mem___dcache___mem_master_awburst = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [17:16]; 
  assign  RTL___near_mem___dcache___mem_master_awlock = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [15]; 
  assign  RTL___near_mem___dcache___mem_master_awcache = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [14:11]; 
  assign  RTL___near_mem___dcache___mem_master_awprot = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [10:8]; 
  assign  RTL___near_mem___dcache___mem_master_awqos = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [7:4]; 
  assign  RTL___near_mem___dcache___mem_master_awregion = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT [3:0]; 
  assign  RTL___near_mem___dcache___CAN_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL___near_mem___dcache___mem_master_wvalid = RTL___near_mem___dcache___master_xactor_f_wr_data$EMPTY_N ; 
  assign  RTL___near_mem___dcache___mem_master_wdata = RTL___near_mem___dcache___master_xactor_f_wr_data$D_OUT [72:9]; 
  assign  RTL___near_mem___dcache___mem_master_wstrb = RTL___near_mem___dcache___master_xactor_f_wr_data$D_OUT [8:1]; 
  assign  RTL___near_mem___dcache___mem_master_wlast = RTL___near_mem___dcache___master_xactor_f_wr_data$D_OUT [0]; 
  assign  RTL___near_mem___dcache___CAN_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL___near_mem___dcache___CAN_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___dcache___mem_master_bready = RTL___near_mem___dcache___master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL___near_mem___dcache___mem_master_arvalid = RTL___near_mem___dcache___master_xactor_f_rd_addr$EMPTY_N ; 
  assign  RTL___near_mem___dcache___mem_master_arid = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [96:93]; 
  assign  RTL___near_mem___dcache___mem_master_araddr = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [92:29]; 
  assign  RTL___near_mem___dcache___mem_master_arlen = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [28:21]; 
  assign  RTL___near_mem___dcache___mem_master_arsize = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [20:18]; 
  assign  RTL___near_mem___dcache___mem_master_arburst = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [17:16]; 
  assign  RTL___near_mem___dcache___mem_master_arlock = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [15]; 
  assign  RTL___near_mem___dcache___mem_master_arcache = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [14:11]; 
  assign  RTL___near_mem___dcache___mem_master_arprot = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [10:8]; 
  assign  RTL___near_mem___dcache___mem_master_arqos = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [7:4]; 
  assign  RTL___near_mem___dcache___mem_master_arregion = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT [3:0]; 
  assign  RTL___near_mem___dcache___CAN_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL___near_mem___dcache___CAN_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___dcache___mem_master_rready = RTL___near_mem___dcache___master_xactor_f_rd_data$FULL_N ;  
    wire RTL___near_mem___dcache___f_fabric_write_reqs___CLK;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RST;
    wire[RTL___near_mem___dcache___f_fabric_write_reqs___width-1:0] RTL___near_mem___dcache___f_fabric_write_reqs___D_IN;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___ENQ;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___DEQ;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___CLR;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___FULL_N;
    wire RTL___near_mem___dcache___f_fabric_write_reqs___EMPTY_N;
    wire[RTL___near_mem___dcache___f_fabric_write_reqs___width-1:0] RTL___near_mem___dcache___f_fabric_write_reqs___D_OUT;
    wire RTL___near_mem___dcache___f_reset_reqs___CLK;
    wire RTL___near_mem___dcache___f_reset_reqs___RST;
    wire[RTL___near_mem___dcache___f_reset_reqs___width-1:0] RTL___near_mem___dcache___f_reset_reqs___D_IN;
    wire RTL___near_mem___dcache___f_reset_reqs___ENQ;
    wire RTL___near_mem___dcache___f_reset_reqs___DEQ;
    wire RTL___near_mem___dcache___f_reset_reqs___CLR;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_reqs___FULL_N;
    wire RTL___near_mem___dcache___f_reset_reqs___EMPTY_N;
    wire[RTL___near_mem___dcache___f_reset_reqs___width-1:0] RTL___near_mem___dcache___f_reset_reqs___D_OUT;
    wire RTL___near_mem___dcache___f_reset_rsps___CLK;
    wire RTL___near_mem___dcache___f_reset_rsps___RST;
    wire[RTL___near_mem___dcache___f_reset_rsps___width-1:0] RTL___near_mem___dcache___f_reset_rsps___D_IN;
    wire RTL___near_mem___dcache___f_reset_rsps___ENQ;
    wire RTL___near_mem___dcache___f_reset_rsps___DEQ;
    wire RTL___near_mem___dcache___f_reset_rsps___CLR;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___f_reset_rsps___FULL_N;
    wire RTL___near_mem___dcache___f_reset_rsps___EMPTY_N;
    wire[RTL___near_mem___dcache___f_reset_rsps___width-1:0] RTL___near_mem___dcache___f_reset_rsps___D_OUT;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___CLK;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RST;
    wire[RTL___near_mem___dcache___master_xactor_f_rd_addr___width-1:0] RTL___near_mem___dcache___master_xactor_f_rd_addr___D_IN;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___CLR;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___FULL_N;
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___EMPTY_N;
    wire[RTL___near_mem___dcache___master_xactor_f_rd_addr___width-1:0] RTL___near_mem___dcache___master_xactor_f_rd_addr___D_OUT;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___CLK;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RST;
    wire[RTL___near_mem___dcache___master_xactor_f_rd_data___width-1:0] RTL___near_mem___dcache___master_xactor_f_rd_data___D_IN;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___CLR;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___FULL_N;
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___EMPTY_N;
    wire[RTL___near_mem___dcache___master_xactor_f_rd_data___width-1:0] RTL___near_mem___dcache___master_xactor_f_rd_data___D_OUT;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___CLK;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RST;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_addr___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_addr___D_IN;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___CLR;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___FULL_N;
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___EMPTY_N;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_addr___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_addr___D_OUT;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___CLK;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RST;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_data___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_data___D_IN;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___CLR;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___FULL_N;
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___EMPTY_N;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_data___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_data___D_OUT;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___CLK;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RST;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_resp___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_resp___D_IN;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___CLR;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___FULL_N;
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___EMPTY_N;
    wire[RTL___near_mem___dcache___master_xactor_f_wr_resp___width-1:0] RTL___near_mem___dcache___master_xactor_f_wr_resp___D_OUT;
    wire RTL___near_mem___icache___f_fabric_write_reqs___CLK;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RST;
    wire[RTL___near_mem___icache___f_fabric_write_reqs___width-1:0] RTL___near_mem___icache___f_fabric_write_reqs___D_IN;
    wire RTL___near_mem___icache___f_fabric_write_reqs___ENQ;
    wire RTL___near_mem___icache___f_fabric_write_reqs___DEQ;
    wire RTL___near_mem___icache___f_fabric_write_reqs___CLR;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_fabric_write_reqs___FULL_N;
    wire RTL___near_mem___icache___f_fabric_write_reqs___EMPTY_N;
    wire[RTL___near_mem___icache___f_fabric_write_reqs___width-1:0] RTL___near_mem___icache___f_fabric_write_reqs___D_OUT;
    wire RTL___near_mem___icache___f_reset_reqs___CLK;
    wire RTL___near_mem___icache___f_reset_reqs___RST;
    wire[RTL___near_mem___icache___f_reset_reqs___width-1:0] RTL___near_mem___icache___f_reset_reqs___D_IN;
    wire RTL___near_mem___icache___f_reset_reqs___ENQ;
    wire RTL___near_mem___icache___f_reset_reqs___DEQ;
    wire RTL___near_mem___icache___f_reset_reqs___CLR;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_reqs___FULL_N;
    wire RTL___near_mem___icache___f_reset_reqs___EMPTY_N;
    wire[RTL___near_mem___icache___f_reset_reqs___width-1:0] RTL___near_mem___icache___f_reset_reqs___D_OUT;
    wire RTL___near_mem___icache___f_reset_rsps___CLK;
    wire RTL___near_mem___icache___f_reset_rsps___RST;
    wire[RTL___near_mem___icache___f_reset_rsps___width-1:0] RTL___near_mem___icache___f_reset_rsps___D_IN;
    wire RTL___near_mem___icache___f_reset_rsps___ENQ;
    wire RTL___near_mem___icache___f_reset_rsps___DEQ;
    wire RTL___near_mem___icache___f_reset_rsps___CLR;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___f_reset_rsps___FULL_N;
    wire RTL___near_mem___icache___f_reset_rsps___EMPTY_N;
    wire[RTL___near_mem___icache___f_reset_rsps___width-1:0] RTL___near_mem___icache___f_reset_rsps___D_OUT;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___CLK;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RST;
    wire[RTL___near_mem___icache___master_xactor_f_rd_addr___width-1:0] RTL___near_mem___icache___master_xactor_f_rd_addr___D_IN;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___CLR;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___FULL_N;
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___EMPTY_N;
    wire[RTL___near_mem___icache___master_xactor_f_rd_addr___width-1:0] RTL___near_mem___icache___master_xactor_f_rd_addr___D_OUT;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___CLK;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RST;
    wire[RTL___near_mem___icache___master_xactor_f_rd_data___width-1:0] RTL___near_mem___icache___master_xactor_f_rd_data___D_IN;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___ENQ;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___DEQ;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___CLR;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___FULL_N;
    wire RTL___near_mem___icache___master_xactor_f_rd_data___EMPTY_N;
    wire[RTL___near_mem___icache___master_xactor_f_rd_data___width-1:0] RTL___near_mem___icache___master_xactor_f_rd_data___D_OUT;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___CLK;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RST;
    wire[RTL___near_mem___icache___master_xactor_f_wr_addr___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_addr___D_IN;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___CLR;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___FULL_N;
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___EMPTY_N;
    wire[RTL___near_mem___icache___master_xactor_f_wr_addr___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_addr___D_OUT;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___CLK;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RST;
    wire[RTL___near_mem___icache___master_xactor_f_wr_data___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_data___D_IN;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___ENQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___DEQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___CLR;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___FULL_N;
    wire RTL___near_mem___icache___master_xactor_f_wr_data___EMPTY_N;
    wire[RTL___near_mem___icache___master_xactor_f_wr_data___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_data___D_OUT;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___CLK;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RST;
    wire[RTL___near_mem___icache___master_xactor_f_wr_resp___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_resp___D_IN;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___CLR;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___FULL_N;
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___EMPTY_N;
    wire[RTL___near_mem___icache___master_xactor_f_wr_resp___width-1:0] RTL___near_mem___icache___master_xactor_f_wr_resp___D_OUT;

    reg RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
    reg RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; reg[ RTL___near_mem___dcache___f_fabric_write_reqs___width -1:0] RTL___near_mem___dcache___f_fabric_write_reqs___data0_reg ; reg[ RTL___near_mem___dcache___f_fabric_write_reqs___width -1:0] RTL___near_mem___dcache___f_fabric_write_reqs___data1_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___FULL_N = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___EMPTY_N = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___D_OUT = RTL___near_mem___dcache___f_fabric_write_reqs___data0_reg ; 
    wire RTL___near_mem___dcache___f_fabric_write_reqs___d0di =( RTL___near_mem___dcache___f_fabric_write_reqs___ENQ &&! RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg )||( RTL___near_mem___dcache___f_fabric_write_reqs___ENQ && RTL___near_mem___dcache___f_fabric_write_reqs___DEQ && RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ); 
    wire RTL___near_mem___dcache___f_fabric_write_reqs___d0d1 = RTL___near_mem___dcache___f_fabric_write_reqs___DEQ &&! RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
    wire RTL___near_mem___dcache___f_fabric_write_reqs___d0h =((! RTL___near_mem___dcache___f_fabric_write_reqs___DEQ )&&(! RTL___near_mem___dcache___f_fabric_write_reqs___ENQ ))||(! RTL___near_mem___dcache___f_fabric_write_reqs___DEQ && RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg )||(! RTL___near_mem___dcache___f_fabric_write_reqs___ENQ && RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ); 
    wire RTL___near_mem___dcache___f_fabric_write_reqs___d1di = RTL___near_mem___dcache___f_fabric_write_reqs___ENQ & RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___f_fabric_write_reqs___CLK )
         begin 
             if ( RTL___near_mem___dcache___f_fabric_write_reqs___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___f_fabric_write_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___f_fabric_write_reqs___CLR )
                         begin  
                             RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___f_fabric_write_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___f_fabric_write_reqs___ENQ &&! RTL___near_mem___dcache___f_fabric_write_reqs___DEQ )
                             begin  
                                 RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___f_fabric_write_reqs___full_reg  <=! RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___f_fabric_write_reqs___DEQ &&! RTL___near_mem___dcache___f_fabric_write_reqs___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___f_fabric_write_reqs___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg  <=! RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___f_fabric_write_reqs___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___f_fabric_write_reqs___data0_reg  <={ RTL___near_mem___dcache___f_fabric_write_reqs___width { RTL___near_mem___dcache___f_fabric_write_reqs___d0di }}& RTL___near_mem___dcache___f_fabric_write_reqs___D_IN |{ RTL___near_mem___dcache___f_fabric_write_reqs___width { RTL___near_mem___dcache___f_fabric_write_reqs___d0d1 }}& RTL___near_mem___dcache___f_fabric_write_reqs___data1_reg |{ RTL___near_mem___dcache___f_fabric_write_reqs___width { RTL___near_mem___dcache___f_fabric_write_reqs___d0h }}& RTL___near_mem___dcache___f_fabric_write_reqs___data0_reg ; 
                 RTL___near_mem___dcache___f_fabric_write_reqs___data1_reg  <= RTL___near_mem___dcache___f_fabric_write_reqs___d1di  ?  RTL___near_mem___dcache___f_fabric_write_reqs___D_IN : RTL___near_mem___dcache___f_fabric_write_reqs___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___f_fabric_write_reqs___CLK )
         begin : RTL___near_mem___dcache___f_fabric_write_reqs___error_checks 
           reg RTL___near_mem___dcache___f_fabric_write_reqs___deqerror , RTL___near_mem___dcache___f_fabric_write_reqs___enqerror ; 
             RTL___near_mem___dcache___f_fabric_write_reqs___deqerror  =0; 
             RTL___near_mem___dcache___f_fabric_write_reqs___enqerror  =0;
             if ( RTL___near_mem___dcache___f_fabric_write_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg && RTL___near_mem___dcache___f_fabric_write_reqs___DEQ )
                         begin  
                             RTL___near_mem___dcache___f_fabric_write_reqs___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___f_fabric_write_reqs___full_reg && RTL___near_mem___dcache___f_fabric_write_reqs___ENQ &&(! RTL___near_mem___dcache___f_fabric_write_reqs___DEQ || RTL___near_mem___dcache___f_fabric_write_reqs___guarded ))
                         begin  
                             RTL___near_mem___dcache___f_fabric_write_reqs___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___empty_reg ;
    reg RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
    reg RTL___near_mem___dcache___f_reset_reqs___empty_reg ; reg[ RTL___near_mem___dcache___f_reset_reqs___width -1:0] RTL___near_mem___dcache___f_reset_reqs___data0_reg ; reg[ RTL___near_mem___dcache___f_reset_reqs___width -1:0] RTL___near_mem___dcache___f_reset_reqs___data1_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___FULL_N = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___EMPTY_N = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___D_OUT = RTL___near_mem___dcache___f_reset_reqs___data0_reg ; 
    wire RTL___near_mem___dcache___f_reset_reqs___d0di =( RTL___near_mem___dcache___f_reset_reqs___ENQ &&! RTL___near_mem___dcache___f_reset_reqs___empty_reg )||( RTL___near_mem___dcache___f_reset_reqs___ENQ && RTL___near_mem___dcache___f_reset_reqs___DEQ && RTL___near_mem___dcache___f_reset_reqs___full_reg ); 
    wire RTL___near_mem___dcache___f_reset_reqs___d0d1 = RTL___near_mem___dcache___f_reset_reqs___DEQ &&! RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
    wire RTL___near_mem___dcache___f_reset_reqs___d0h =((! RTL___near_mem___dcache___f_reset_reqs___DEQ )&&(! RTL___near_mem___dcache___f_reset_reqs___ENQ ))||(! RTL___near_mem___dcache___f_reset_reqs___DEQ && RTL___near_mem___dcache___f_reset_reqs___empty_reg )||(! RTL___near_mem___dcache___f_reset_reqs___ENQ && RTL___near_mem___dcache___f_reset_reqs___full_reg ); 
    wire RTL___near_mem___dcache___f_reset_reqs___d1di = RTL___near_mem___dcache___f_reset_reqs___ENQ & RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___f_reset_reqs___CLK )
         begin 
             if ( RTL___near_mem___dcache___f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___f_reset_reqs___CLR )
                         begin  
                             RTL___near_mem___dcache___f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___f_reset_reqs___ENQ &&! RTL___near_mem___dcache___f_reset_reqs___DEQ )
                             begin  
                                 RTL___near_mem___dcache___f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___f_reset_reqs___full_reg  <=! RTL___near_mem___dcache___f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___f_reset_reqs___DEQ &&! RTL___near_mem___dcache___f_reset_reqs___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___f_reset_reqs___empty_reg  <=! RTL___near_mem___dcache___f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___f_reset_reqs___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___f_reset_reqs___data0_reg  <={ RTL___near_mem___dcache___f_reset_reqs___width { RTL___near_mem___dcache___f_reset_reqs___d0di }}& RTL___near_mem___dcache___f_reset_reqs___D_IN |{ RTL___near_mem___dcache___f_reset_reqs___width { RTL___near_mem___dcache___f_reset_reqs___d0d1 }}& RTL___near_mem___dcache___f_reset_reqs___data1_reg |{ RTL___near_mem___dcache___f_reset_reqs___width { RTL___near_mem___dcache___f_reset_reqs___d0h }}& RTL___near_mem___dcache___f_reset_reqs___data0_reg ; 
                 RTL___near_mem___dcache___f_reset_reqs___data1_reg  <= RTL___near_mem___dcache___f_reset_reqs___d1di  ?  RTL___near_mem___dcache___f_reset_reqs___D_IN : RTL___near_mem___dcache___f_reset_reqs___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___f_reset_reqs___CLK )
         begin : RTL___near_mem___dcache___f_reset_reqs___error_checks 
           reg RTL___near_mem___dcache___f_reset_reqs___deqerror , RTL___near_mem___dcache___f_reset_reqs___enqerror ; 
             RTL___near_mem___dcache___f_reset_reqs___deqerror  =0; 
             RTL___near_mem___dcache___f_reset_reqs___enqerror  =0;
             if ( RTL___near_mem___dcache___f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___f_reset_reqs___empty_reg && RTL___near_mem___dcache___f_reset_reqs___DEQ )
                         begin  
                             RTL___near_mem___dcache___f_reset_reqs___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___f_reset_reqs___full_reg && RTL___near_mem___dcache___f_reset_reqs___ENQ &&(! RTL___near_mem___dcache___f_reset_reqs___DEQ || RTL___near_mem___dcache___f_reset_reqs___guarded ))
                         begin  
                             RTL___near_mem___dcache___f_reset_reqs___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___empty_reg ;
    reg RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
    reg RTL___near_mem___dcache___f_reset_rsps___empty_reg ; reg[ RTL___near_mem___dcache___f_reset_rsps___width -1:0] RTL___near_mem___dcache___f_reset_rsps___data0_reg ; reg[ RTL___near_mem___dcache___f_reset_rsps___width -1:0] RTL___near_mem___dcache___f_reset_rsps___data1_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___FULL_N = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___EMPTY_N = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___D_OUT = RTL___near_mem___dcache___f_reset_rsps___data0_reg ; 
    wire RTL___near_mem___dcache___f_reset_rsps___d0di =( RTL___near_mem___dcache___f_reset_rsps___ENQ &&! RTL___near_mem___dcache___f_reset_rsps___empty_reg )||( RTL___near_mem___dcache___f_reset_rsps___ENQ && RTL___near_mem___dcache___f_reset_rsps___DEQ && RTL___near_mem___dcache___f_reset_rsps___full_reg ); 
    wire RTL___near_mem___dcache___f_reset_rsps___d0d1 = RTL___near_mem___dcache___f_reset_rsps___DEQ &&! RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
    wire RTL___near_mem___dcache___f_reset_rsps___d0h =((! RTL___near_mem___dcache___f_reset_rsps___DEQ )&&(! RTL___near_mem___dcache___f_reset_rsps___ENQ ))||(! RTL___near_mem___dcache___f_reset_rsps___DEQ && RTL___near_mem___dcache___f_reset_rsps___empty_reg )||(! RTL___near_mem___dcache___f_reset_rsps___ENQ && RTL___near_mem___dcache___f_reset_rsps___full_reg ); 
    wire RTL___near_mem___dcache___f_reset_rsps___d1di = RTL___near_mem___dcache___f_reset_rsps___ENQ & RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___f_reset_rsps___CLK )
         begin 
             if ( RTL___near_mem___dcache___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___f_reset_rsps___CLR )
                         begin  
                             RTL___near_mem___dcache___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___f_reset_rsps___ENQ &&! RTL___near_mem___dcache___f_reset_rsps___DEQ )
                             begin  
                                 RTL___near_mem___dcache___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___f_reset_rsps___full_reg  <=! RTL___near_mem___dcache___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___f_reset_rsps___DEQ &&! RTL___near_mem___dcache___f_reset_rsps___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___f_reset_rsps___empty_reg  <=! RTL___near_mem___dcache___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___f_reset_rsps___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___f_reset_rsps___data0_reg  <={ RTL___near_mem___dcache___f_reset_rsps___width { RTL___near_mem___dcache___f_reset_rsps___d0di }}& RTL___near_mem___dcache___f_reset_rsps___D_IN |{ RTL___near_mem___dcache___f_reset_rsps___width { RTL___near_mem___dcache___f_reset_rsps___d0d1 }}& RTL___near_mem___dcache___f_reset_rsps___data1_reg |{ RTL___near_mem___dcache___f_reset_rsps___width { RTL___near_mem___dcache___f_reset_rsps___d0h }}& RTL___near_mem___dcache___f_reset_rsps___data0_reg ; 
                 RTL___near_mem___dcache___f_reset_rsps___data1_reg  <= RTL___near_mem___dcache___f_reset_rsps___d1di  ?  RTL___near_mem___dcache___f_reset_rsps___D_IN : RTL___near_mem___dcache___f_reset_rsps___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___f_reset_rsps___CLK )
         begin : RTL___near_mem___dcache___f_reset_rsps___error_checks 
           reg RTL___near_mem___dcache___f_reset_rsps___deqerror , RTL___near_mem___dcache___f_reset_rsps___enqerror ; 
             RTL___near_mem___dcache___f_reset_rsps___deqerror  =0; 
             RTL___near_mem___dcache___f_reset_rsps___enqerror  =0;
             if ( RTL___near_mem___dcache___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___f_reset_rsps___empty_reg && RTL___near_mem___dcache___f_reset_rsps___DEQ )
                         begin  
                             RTL___near_mem___dcache___f_reset_rsps___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___f_reset_rsps___full_reg && RTL___near_mem___dcache___f_reset_rsps___ENQ &&(! RTL___near_mem___dcache___f_reset_rsps___DEQ || RTL___near_mem___dcache___f_reset_rsps___guarded ))
                         begin  
                             RTL___near_mem___dcache___f_reset_rsps___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___empty_reg ;
    reg RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
    reg RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_rd_addr___width -1:0] RTL___near_mem___dcache___master_xactor_f_rd_addr___data0_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_rd_addr___width -1:0] RTL___near_mem___dcache___master_xactor_f_rd_addr___data1_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___FULL_N = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___EMPTY_N = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___D_OUT = RTL___near_mem___dcache___master_xactor_f_rd_addr___data0_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___d0di =( RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ &&! RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg )||( RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ && RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ && RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___d0d1 = RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ &&! RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___d0h =((! RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ )&&(! RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ ))||(! RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ && RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg )||(! RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ && RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_rd_addr___d1di = RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ & RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_addr___CLK )
         begin 
             if ( RTL___near_mem___dcache___master_xactor_f_rd_addr___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___master_xactor_f_rd_addr___CLR )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ &&! RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ )
                             begin  
                                 RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg  <=! RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ &&! RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg  <=! RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_addr___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___master_xactor_f_rd_addr___data0_reg  <={ RTL___near_mem___dcache___master_xactor_f_rd_addr___width { RTL___near_mem___dcache___master_xactor_f_rd_addr___d0di }}& RTL___near_mem___dcache___master_xactor_f_rd_addr___D_IN |{ RTL___near_mem___dcache___master_xactor_f_rd_addr___width { RTL___near_mem___dcache___master_xactor_f_rd_addr___d0d1 }}& RTL___near_mem___dcache___master_xactor_f_rd_addr___data1_reg |{ RTL___near_mem___dcache___master_xactor_f_rd_addr___width { RTL___near_mem___dcache___master_xactor_f_rd_addr___d0h }}& RTL___near_mem___dcache___master_xactor_f_rd_addr___data0_reg ; 
                 RTL___near_mem___dcache___master_xactor_f_rd_addr___data1_reg  <= RTL___near_mem___dcache___master_xactor_f_rd_addr___d1di  ?  RTL___near_mem___dcache___master_xactor_f_rd_addr___D_IN : RTL___near_mem___dcache___master_xactor_f_rd_addr___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_addr___CLK )
         begin : RTL___near_mem___dcache___master_xactor_f_rd_addr___error_checks 
           reg RTL___near_mem___dcache___master_xactor_f_rd_addr___deqerror , RTL___near_mem___dcache___master_xactor_f_rd_addr___enqerror ; 
             RTL___near_mem___dcache___master_xactor_f_rd_addr___deqerror  =0; 
             RTL___near_mem___dcache___master_xactor_f_rd_addr___enqerror  =0;
             if ( RTL___near_mem___dcache___master_xactor_f_rd_addr___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg && RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_addr___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg && RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ &&(! RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ || RTL___near_mem___dcache___master_xactor_f_rd_addr___guarded ))
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_addr___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___empty_reg ;
    reg RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
    reg RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_rd_data___width -1:0] RTL___near_mem___dcache___master_xactor_f_rd_data___data0_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_rd_data___width -1:0] RTL___near_mem___dcache___master_xactor_f_rd_data___data1_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___FULL_N = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___EMPTY_N = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___D_OUT = RTL___near_mem___dcache___master_xactor_f_rd_data___data0_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___d0di =( RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ &&! RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg )||( RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ && RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ && RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___d0d1 = RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ &&! RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___d0h =((! RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ )&&(! RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ ))||(! RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ && RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg )||(! RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ && RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_rd_data___d1di = RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ & RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_data___CLK )
         begin 
             if ( RTL___near_mem___dcache___master_xactor_f_rd_data___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___master_xactor_f_rd_data___CLR )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ &&! RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ )
                             begin  
                                 RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg  <=! RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ &&! RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg  <=! RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_data___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___master_xactor_f_rd_data___data0_reg  <={ RTL___near_mem___dcache___master_xactor_f_rd_data___width { RTL___near_mem___dcache___master_xactor_f_rd_data___d0di }}& RTL___near_mem___dcache___master_xactor_f_rd_data___D_IN |{ RTL___near_mem___dcache___master_xactor_f_rd_data___width { RTL___near_mem___dcache___master_xactor_f_rd_data___d0d1 }}& RTL___near_mem___dcache___master_xactor_f_rd_data___data1_reg |{ RTL___near_mem___dcache___master_xactor_f_rd_data___width { RTL___near_mem___dcache___master_xactor_f_rd_data___d0h }}& RTL___near_mem___dcache___master_xactor_f_rd_data___data0_reg ; 
                 RTL___near_mem___dcache___master_xactor_f_rd_data___data1_reg  <= RTL___near_mem___dcache___master_xactor_f_rd_data___d1di  ?  RTL___near_mem___dcache___master_xactor_f_rd_data___D_IN : RTL___near_mem___dcache___master_xactor_f_rd_data___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_rd_data___CLK )
         begin : RTL___near_mem___dcache___master_xactor_f_rd_data___error_checks 
           reg RTL___near_mem___dcache___master_xactor_f_rd_data___deqerror , RTL___near_mem___dcache___master_xactor_f_rd_data___enqerror ; 
             RTL___near_mem___dcache___master_xactor_f_rd_data___deqerror  =0; 
             RTL___near_mem___dcache___master_xactor_f_rd_data___enqerror  =0;
             if ( RTL___near_mem___dcache___master_xactor_f_rd_data___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg && RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_data___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg && RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ &&(! RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ || RTL___near_mem___dcache___master_xactor_f_rd_data___guarded ))
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_rd_data___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___empty_reg ;
    reg RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
    reg RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_addr___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_addr___data0_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_addr___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_addr___data1_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_addr___data0_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___d0di =( RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg )||( RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___d0d1 = RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___d0h =((! RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ )&&(! RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ ))||(! RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg )||(! RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_addr___d1di = RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ & RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_addr___CLK )
         begin 
             if ( RTL___near_mem___dcache___master_xactor_f_wr_addr___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___master_xactor_f_wr_addr___CLR )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ )
                             begin  
                                 RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_addr___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___master_xactor_f_wr_addr___data0_reg  <={ RTL___near_mem___dcache___master_xactor_f_wr_addr___width { RTL___near_mem___dcache___master_xactor_f_wr_addr___d0di }}& RTL___near_mem___dcache___master_xactor_f_wr_addr___D_IN |{ RTL___near_mem___dcache___master_xactor_f_wr_addr___width { RTL___near_mem___dcache___master_xactor_f_wr_addr___d0d1 }}& RTL___near_mem___dcache___master_xactor_f_wr_addr___data1_reg |{ RTL___near_mem___dcache___master_xactor_f_wr_addr___width { RTL___near_mem___dcache___master_xactor_f_wr_addr___d0h }}& RTL___near_mem___dcache___master_xactor_f_wr_addr___data0_reg ; 
                 RTL___near_mem___dcache___master_xactor_f_wr_addr___data1_reg  <= RTL___near_mem___dcache___master_xactor_f_wr_addr___d1di  ?  RTL___near_mem___dcache___master_xactor_f_wr_addr___D_IN : RTL___near_mem___dcache___master_xactor_f_wr_addr___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_addr___CLK )
         begin : RTL___near_mem___dcache___master_xactor_f_wr_addr___error_checks 
           reg RTL___near_mem___dcache___master_xactor_f_wr_addr___deqerror , RTL___near_mem___dcache___master_xactor_f_wr_addr___enqerror ; 
             RTL___near_mem___dcache___master_xactor_f_wr_addr___deqerror  =0; 
             RTL___near_mem___dcache___master_xactor_f_wr_addr___enqerror  =0;
             if ( RTL___near_mem___dcache___master_xactor_f_wr_addr___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg && RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_addr___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg && RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ &&(! RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ || RTL___near_mem___dcache___master_xactor_f_wr_addr___guarded ))
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_addr___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___empty_reg ;
    reg RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
    reg RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_data___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_data___data0_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_data___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_data___data1_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_data___data0_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___d0di =( RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg )||( RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___d0d1 = RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___d0h =((! RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ )&&(! RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ ))||(! RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg )||(! RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_data___d1di = RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ & RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_data___CLK )
         begin 
             if ( RTL___near_mem___dcache___master_xactor_f_wr_data___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___master_xactor_f_wr_data___CLR )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ )
                             begin  
                                 RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_data___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___master_xactor_f_wr_data___data0_reg  <={ RTL___near_mem___dcache___master_xactor_f_wr_data___width { RTL___near_mem___dcache___master_xactor_f_wr_data___d0di }}& RTL___near_mem___dcache___master_xactor_f_wr_data___D_IN |{ RTL___near_mem___dcache___master_xactor_f_wr_data___width { RTL___near_mem___dcache___master_xactor_f_wr_data___d0d1 }}& RTL___near_mem___dcache___master_xactor_f_wr_data___data1_reg |{ RTL___near_mem___dcache___master_xactor_f_wr_data___width { RTL___near_mem___dcache___master_xactor_f_wr_data___d0h }}& RTL___near_mem___dcache___master_xactor_f_wr_data___data0_reg ; 
                 RTL___near_mem___dcache___master_xactor_f_wr_data___data1_reg  <= RTL___near_mem___dcache___master_xactor_f_wr_data___d1di  ?  RTL___near_mem___dcache___master_xactor_f_wr_data___D_IN : RTL___near_mem___dcache___master_xactor_f_wr_data___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_data___CLK )
         begin : RTL___near_mem___dcache___master_xactor_f_wr_data___error_checks 
           reg RTL___near_mem___dcache___master_xactor_f_wr_data___deqerror , RTL___near_mem___dcache___master_xactor_f_wr_data___enqerror ; 
             RTL___near_mem___dcache___master_xactor_f_wr_data___deqerror  =0; 
             RTL___near_mem___dcache___master_xactor_f_wr_data___enqerror  =0;
             if ( RTL___near_mem___dcache___master_xactor_f_wr_data___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg && RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_data___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg && RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ &&(! RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ || RTL___near_mem___dcache___master_xactor_f_wr_data___guarded ))
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_data___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___empty_reg ;
    reg RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
    reg RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_resp___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_resp___data0_reg ; reg[ RTL___near_mem___dcache___master_xactor_f_wr_resp___width -1:0] RTL___near_mem___dcache___master_xactor_f_wr_resp___data1_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_resp___data0_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___d0di =( RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg )||( RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___d0d1 = RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___d0h =((! RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ )&&(! RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ ))||(! RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ && RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg )||(! RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ && RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ); 
    wire RTL___near_mem___dcache___master_xactor_f_wr_resp___d1di = RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ & RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_resp___CLK )
         begin 
             if ( RTL___near_mem___dcache___master_xactor_f_wr_resp___RST ==1'b0)
                 begin  
                     RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg  <=1'b0; 
                     RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___master_xactor_f_wr_resp___CLR )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg  <=1'b0; 
                             RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ &&! RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ )
                             begin  
                                 RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg  <=1'b1; 
                                 RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ &&! RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ )
                                 begin  
                                     RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg  <=1'b1; 
                                     RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg  <=! RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_resp___CLK )
         begin 
             begin  
                 RTL___near_mem___dcache___master_xactor_f_wr_resp___data0_reg  <={ RTL___near_mem___dcache___master_xactor_f_wr_resp___width { RTL___near_mem___dcache___master_xactor_f_wr_resp___d0di }}& RTL___near_mem___dcache___master_xactor_f_wr_resp___D_IN |{ RTL___near_mem___dcache___master_xactor_f_wr_resp___width { RTL___near_mem___dcache___master_xactor_f_wr_resp___d0d1 }}& RTL___near_mem___dcache___master_xactor_f_wr_resp___data1_reg |{ RTL___near_mem___dcache___master_xactor_f_wr_resp___width { RTL___near_mem___dcache___master_xactor_f_wr_resp___d0h }}& RTL___near_mem___dcache___master_xactor_f_wr_resp___data0_reg ; 
                 RTL___near_mem___dcache___master_xactor_f_wr_resp___data1_reg  <= RTL___near_mem___dcache___master_xactor_f_wr_resp___d1di  ?  RTL___near_mem___dcache___master_xactor_f_wr_resp___D_IN : RTL___near_mem___dcache___master_xactor_f_wr_resp___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___dcache___master_xactor_f_wr_resp___CLK )
         begin : RTL___near_mem___dcache___master_xactor_f_wr_resp___error_checks 
           reg RTL___near_mem___dcache___master_xactor_f_wr_resp___deqerror , RTL___near_mem___dcache___master_xactor_f_wr_resp___enqerror ; 
             RTL___near_mem___dcache___master_xactor_f_wr_resp___deqerror  =0; 
             RTL___near_mem___dcache___master_xactor_f_wr_resp___enqerror  =0;
             if ( RTL___near_mem___dcache___master_xactor_f_wr_resp___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg && RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ )
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_resp___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg && RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ &&(! RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ || RTL___near_mem___dcache___master_xactor_f_wr_resp___guarded ))
                         begin  
                             RTL___near_mem___dcache___master_xactor_f_wr_resp___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___empty_reg ;
      
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKA;
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___ENA;
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___WEA;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDR_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDRA;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DIA;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA;
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKB;
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___ENB;
    wire RTL___near_mem___dcache___ram_state_and_ctag_cset___WEB;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDR_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDRB;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DIB;
    wire[RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB;
    wire RTL___near_mem___dcache___ram_word64_set___CLKA;
    wire RTL___near_mem___dcache___ram_word64_set___ENA;
    wire RTL___near_mem___dcache___ram_word64_set___WEA;
    wire[RTL___near_mem___dcache___ram_word64_set___ADDR_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___ADDRA;
    wire[RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___DIA;
    wire[RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___DOA;
    wire RTL___near_mem___dcache___ram_word64_set___CLKB;
    wire RTL___near_mem___dcache___ram_word64_set___ENB;
    wire RTL___near_mem___dcache___ram_word64_set___WEB;
    wire[RTL___near_mem___dcache___ram_word64_set___ADDR_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___ADDRB;
    wire[RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___DIB;
    wire[RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___dcache___ram_word64_set___DOB;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___CLKA;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___ENA;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___WEA;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___ADDR_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___ADDRA;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DIA;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOA;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___CLKB;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___ENB;
    wire RTL___near_mem___icache___ram_state_and_ctag_cset___WEB;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___ADDR_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___ADDRB;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DIB;
    wire[RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOB;
    wire RTL___near_mem___icache___ram_word64_set___CLKA;
    wire RTL___near_mem___icache___ram_word64_set___ENA;
    wire RTL___near_mem___icache___ram_word64_set___WEA;
    wire[RTL___near_mem___icache___ram_word64_set___ADDR_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___ADDRA;
    wire[RTL___near_mem___icache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___DIA;
    wire[RTL___near_mem___icache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___DOA;
    wire RTL___near_mem___icache___ram_word64_set___CLKB;
    wire RTL___near_mem___icache___ram_word64_set___ENB;
    wire RTL___near_mem___icache___ram_word64_set___WEB;
    wire[RTL___near_mem___icache___ram_word64_set___ADDR_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___ADDRB;
    wire[RTL___near_mem___icache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___DIB;
    wire[RTL___near_mem___icache___ram_word64_set___DATA_WIDTH-1:0] RTL___near_mem___icache___ram_word64_set___DOB;

    reg[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R ; reg[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R ; reg[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R2 ; reg[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R2 ; 
    wire[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___arb1 ; 
    wire[ RTL___near_mem___dcache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_state_and_ctag_cset___arb2 ; 
  always @( posedge  RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKA )
         begin 
             if ( RTL___near_mem___dcache___ram_state_and_ctag_cset___ENA )
                 begin 
                     if ( RTL___near_mem___dcache___ram_state_and_ctag_cset___WEA )
                         begin  
                             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___DIA ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___arb1 ;
                         end 
                 end  
             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R2  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R ;
         end
  always @( posedge  RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKB )
         begin 
             if ( RTL___near_mem___dcache___ram_state_and_ctag_cset___ENB )
                 begin 
                     if ( RTL___near_mem___dcache___ram_state_and_ctag_cset___WEB )
                         begin  
                             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___DIB ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___arb2 ;
                         end 
                 end  
             RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R2  <= RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R ;
         end
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA =( RTL___near_mem___dcache___ram_state_and_ctag_cset___PIPELINED ) ?  RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R2 : RTL___near_mem___dcache___ram_state_and_ctag_cset___DOA_R ; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB =( RTL___near_mem___dcache___ram_state_and_ctag_cset___PIPELINED ) ?  RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R2 : RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB_R ;
    reg[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___DOA_R ; reg[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___DOB_R ; reg[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___DOA_R2 ; reg[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___DOB_R2 ; 
    wire[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___arb1 ; 
    wire[ RTL___near_mem___dcache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___dcache___ram_word64_set___arb2 ; 
  always @( posedge  RTL___near_mem___dcache___ram_word64_set___CLKA )
         begin 
             if ( RTL___near_mem___dcache___ram_word64_set___ENA )
                 begin 
                     if ( RTL___near_mem___dcache___ram_word64_set___WEA )
                         begin  
                             RTL___near_mem___dcache___ram_word64_set___DOA_R  <= RTL___near_mem___dcache___ram_word64_set___DIA ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___dcache___ram_word64_set___DOA_R  <= RTL___near_mem___dcache___ram_word64_set___arb1 ;
                         end 
                 end  
             RTL___near_mem___dcache___ram_word64_set___DOA_R2  <= RTL___near_mem___dcache___ram_word64_set___DOA_R ;
         end
  always @( posedge  RTL___near_mem___dcache___ram_word64_set___CLKB )
         begin 
             if ( RTL___near_mem___dcache___ram_word64_set___ENB )
                 begin 
                     if ( RTL___near_mem___dcache___ram_word64_set___WEB )
                         begin  
                             RTL___near_mem___dcache___ram_word64_set___DOB_R  <= RTL___near_mem___dcache___ram_word64_set___DIB ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___dcache___ram_word64_set___DOB_R  <= RTL___near_mem___dcache___ram_word64_set___arb2 ;
                         end 
                 end  
             RTL___near_mem___dcache___ram_word64_set___DOB_R2  <= RTL___near_mem___dcache___ram_word64_set___DOB_R ;
         end
  assign  RTL___near_mem___dcache___ram_word64_set___DOA =( RTL___near_mem___dcache___ram_word64_set___PIPELINED ) ?  RTL___near_mem___dcache___ram_word64_set___DOA_R2 : RTL___near_mem___dcache___ram_word64_set___DOA_R ; 
  assign  RTL___near_mem___dcache___ram_word64_set___DOB =( RTL___near_mem___dcache___ram_word64_set___PIPELINED ) ?  RTL___near_mem___dcache___ram_word64_set___DOB_R2 : RTL___near_mem___dcache___ram_word64_set___DOB_R ;
      
    wire RTL___near_mem___dcache___soc_map___CLK;
    wire RTL___near_mem___dcache___soc_map___RST_N;
    wire[63:0] RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr;
    wire[63:0] RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr;
    wire[63:0] RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr_addr;
    wire RTL___near_mem___icache___soc_map___CLK;
    wire RTL___near_mem___icache___soc_map___RST_N;
    wire[63:0] RTL___near_mem___icache___soc_map___m_is_mem_addr_addr;
    wire[63:0] RTL___near_mem___icache___soc_map___m_is_IO_addr_addr;
    wire[63:0] RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr_addr;
    wire RTL___near_mem___soc_map___CLK;
    wire RTL___near_mem___soc_map___RST_N;
    wire[63:0] RTL___near_mem___soc_map___m_is_mem_addr_addr;
    wire[63:0] RTL___near_mem___soc_map___m_is_IO_addr_addr;
    wire[63:0] RTL___near_mem___soc_map___m_is_near_mem_IO_addr_addr;

    wire[63:0] RTL___near_mem___dcache___soc_map___m_boot_rom_addr_base , RTL___near_mem___dcache___soc_map___m_boot_rom_addr_lim , RTL___near_mem___dcache___soc_map___m_boot_rom_addr_size , RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_base , RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_lim , RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_size , RTL___near_mem___dcache___soc_map___m_mtvec_reset_value , RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_base , RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_lim , RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_size , RTL___near_mem___dcache___soc_map___m_nmivec_reset_value , RTL___near_mem___dcache___soc_map___m_pc_reset_value , RTL___near_mem___dcache___soc_map___m_plic_addr_base , RTL___near_mem___dcache___soc_map___m_plic_addr_lim , RTL___near_mem___dcache___soc_map___m_plic_addr_size , RTL___near_mem___dcache___soc_map___m_tcm_addr_base , RTL___near_mem___dcache___soc_map___m_tcm_addr_lim , RTL___near_mem___dcache___soc_map___m_tcm_addr_size , RTL___near_mem___dcache___soc_map___m_uart0_addr_base , RTL___near_mem___dcache___soc_map___m_uart0_addr_lim , RTL___near_mem___dcache___soc_map___m_uart0_addr_size ; 
    wire RTL___near_mem___dcache___soc_map___m_is_IO_addr , RTL___near_mem___dcache___soc_map___m_is_mem_addr , RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr ; 
  assign  RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL___near_mem___dcache___soc_map___m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL___near_mem___dcache___soc_map___m_plic_addr_base =64'h000000000C000000; 
  assign  RTL___near_mem___dcache___soc_map___m_plic_addr_size =64'h0000000000400000; 
  assign  RTL___near_mem___dcache___soc_map___m_plic_addr_lim =64'd205520896; 
  assign  RTL___near_mem___dcache___soc_map___m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL___near_mem___dcache___soc_map___m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL___near_mem___dcache___soc_map___m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL___near_mem___dcache___soc_map___m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL___near_mem___dcache___soc_map___m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL___near_mem___dcache___soc_map___m_boot_rom_addr_lim =64'd8192; 
  assign  RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL___near_mem___dcache___soc_map___m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL___near_mem___dcache___soc_map___m_tcm_addr_base =64'h0; 
  assign  RTL___near_mem___dcache___soc_map___m_tcm_addr_size =64'd0; 
  assign  RTL___near_mem___dcache___soc_map___m_tcm_addr_lim =64'd0; 
  assign  RTL___near_mem___dcache___soc_map___m_is_mem_addr = RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr >=64'h0000000000001000&& RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr <64'd8192|| RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr >=64'h0000000080000000&& RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL___near_mem___dcache___soc_map___m_is_IO_addr = RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr <64'd33603584|| RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr >=64'h000000000C000000&& RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr <64'd205520896|| RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr >=64'h00000000C0000000&& RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr = RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL___near_mem___dcache___soc_map___m_pc_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___dcache___soc_map___m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___dcache___soc_map___m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req = RTL___near_mem___dcache___f_fabric_write_reqs$EMPTY_N && RTL___near_mem___dcache___master_xactor_f_wr_addr$FULL_N && RTL___near_mem___dcache___master_xactor_f_wr_data$FULL_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req = RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_reset =( RTL___near_mem___dcache___rg_cset_in_cache !=7'd127|| RTL___near_mem___dcache___f_reset_reqs$EMPTY_N && RTL___near_mem___dcache___f_reset_rsps$FULL_N )&& RTL___near_mem___dcache___rg_state ==4'd1; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset = RTL___near_mem___dcache___CAN_FIRE_RL_rl_reset ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_probe_and_immed_rsp =( RTL___near_mem___dcache___dmem_not_imem &&! RTL___near_mem___dcache___soc_map$m_is_mem_addr ||! RTL___near_mem___dcache___rg_op || RTL___near_mem___dcache___f_fabric_write_reqs$FULL_N )&& RTL___near_mem___dcache___rg_state ==4'd3; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp = RTL___near_mem___dcache___CAN_FIRE_RL_rl_probe_and_immed_rsp &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_start_cache_refill = RTL___near_mem___dcache___master_xactor_f_rd_addr$FULL_N && RTL___near_mem___dcache___rg_state ==4'd8&& RTL___near_mem___dcache___b__h14485 ==4'd0; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill = RTL___near_mem___dcache___CAN_FIRE_RL_rl_start_cache_refill &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_cache_refill_rsps_loop = RTL___near_mem___dcache___master_xactor_f_rd_data$EMPTY_N && RTL___near_mem___dcache___rg_state ==4'd9; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop = RTL___near_mem___dcache___CAN_FIRE_RL_rl_cache_refill_rsps_loop &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_rereq = RTL___near_mem___dcache___rg_state ==4'd10; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq = RTL___near_mem___dcache___CAN_FIRE_RL_rl_rereq &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_ST_AMO_response = RTL___near_mem___dcache___rg_state ==4'd11; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_ST_AMO_response = RTL___near_mem___dcache___CAN_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_req = RTL___near_mem___dcache___master_xactor_f_rd_addr$FULL_N && RTL___near_mem___dcache___rg_state ==4'd12&&! RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___b__h14485 ==4'd0; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req = RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_req &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_rsp = RTL___near_mem___dcache___master_xactor_f_rd_data$EMPTY_N && RTL___near_mem___dcache___rg_state ==4'd13; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp = RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_read_rsp &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_maintain_io_read_rsp = RTL___near_mem___dcache___rg_state ==4'd14; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp = RTL___near_mem___dcache___CAN_FIRE_RL_rl_maintain_io_read_rsp ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_write_req = RTL___near_mem___dcache___f_fabric_write_reqs$FULL_N && RTL___near_mem___dcache___rg_state ==4'd12&& RTL___near_mem___dcache___rg_op ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req = RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_discard_write_rsp = RTL___near_mem___dcache___b__h14485 !=4'd0&& RTL___near_mem___dcache___master_xactor_f_wr_resp$EMPTY_N ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp = RTL___near_mem___dcache___CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_drive_exception_rsp = RTL___near_mem___dcache___rg_state ==4'd4; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_drive_exception_rsp = RTL___near_mem___dcache___rg_state ==4'd4; 
  assign  RTL___near_mem___dcache___CAN_FIRE_RL_rl_start_reset = RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset = RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_1 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_2 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 ; 
  assign  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__SEL_3 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL___near_mem___dcache___WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__SEL_1 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op ; 
  assign  RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 = RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 ; 
  assign  RTL___near_mem___dcache___MUX_ram_word64_set$a_put_1__SEL_1 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]!=2'd3; 
  assign  RTL___near_mem___dcache___MUX_rg_error_during_refill$write_1__SEL_1 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_1 = RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_2 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_2 = RTL___near_mem___dcache___f_reset_reqs$EMPTY_N && RTL___near_mem___dcache___rg_state !=4'd1; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_3 = RTL___near_mem___dcache___CAN_FIRE_RL_rl_io_write_req &&! RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_7 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]==2'd3; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_9 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 ; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_10 = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127; 
  always @(          RTL___near_mem___dcache___rg_f3                          or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247                 or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276                or   RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32               or   RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___word64__h5094             or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264            or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285           or   RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  )
         begin 
             case ( RTL___near_mem___dcache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 ;
              3 'b001: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 ;
              3 'b010: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 ;
              3 'b011: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  =( RTL___near_mem___dcache___rg_addr [2:0]==3'h0) ?  RTL___near_mem___dcache___word64__h5094 :64'd0;
              3 'b100: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 ;
              3 'b101: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 ;
              3 'b110: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 ;
              3 'd7: 
                  RTL___near_mem___dcache___MUX_dw_output_ld_val$wset_1__VAL_2  =64'd0;endcase
         end
  assign  RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_1 ={ RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_st_amo_val }; 
  assign  RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ={ RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_pa , RTL___near_mem___dcache___rg_st_amo_val }; 
  assign  RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 ={4'd0, RTL___near_mem___dcache___cline_fabric_addr__h14584 ,29'd7143424}; 
  assign  RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ={4'd0, RTL___near_mem___dcache___fabric_addr__h17243 ,8'd0, RTL___near_mem___dcache___value__h17372 ,18'd65536}; 
  assign  RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ={3'd4, RTL___near_mem___dcache___rg_pa [31:12]}; 
  assign  RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_2 = RTL___near_mem___dcache___rg_word64_set_in_cache +9'd1; 
  assign  RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_4 ={ RTL___near_mem___dcache___rg_addr [11:5],2'd0}; 
  assign  RTL___near_mem___dcache___MUX_rg_cset_in_cache$write_1__VAL_1 = RTL___near_mem___dcache___rg_cset_in_cache +7'd1; 
  assign  RTL___near_mem___dcache___MUX_rg_exc_code$write_1__VAL_1 = RTL___near_mem___dcache___req_op  ? 4'd6:4'd4; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_1 = RTL___near_mem___dcache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539  ? 4'd4:4'd3; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_4 =( RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0) ? 4'd14:4'd4; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_7 =( RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___dcache___rg_error_during_refill ) ? 4'd4:4'd10; 
  assign  RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_9 =( RTL___near_mem___dcache___dmem_not_imem &&! RTL___near_mem___dcache___soc_map$m_is_mem_addr ) ? 4'd12:( RTL___near_mem___dcache___rg_op  ? 4'd11:4'd8); 
  assign  RTL___near_mem___dcache___dw_valid$whas = RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 || RTL___near_mem___dcache___WILL_FIRE_RL_rl_drive_exception_rsp || RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL___near_mem___dcache___WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port0__write_1 = RTL___near_mem___dcache___ctr_wr_rsps_pending_crg +4'd1; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port1__write_1 = RTL___near_mem___dcache___b__h14485 -4'd1; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port2__read = RTL___near_mem___dcache___CAN_FIRE_RL_rl_discard_write_rsp  ?  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port1__write_1 : RTL___near_mem___dcache___b__h14485 ; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN_port2__write = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port3__read = RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN_port2__write  ? 4'd0: RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port2__read ; 
  assign  RTL___near_mem___dcache___cfg_verbosity$D_IN = RTL___near_mem___dcache___set_verbosity_verbosity ; 
  assign  RTL___near_mem___dcache___cfg_verbosity$EN = RTL___near_mem___dcache___EN_set_verbosity ; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$D_IN = RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port3__read ; 
  assign  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN =1'b1; 
  assign  RTL___near_mem___dcache___rg_addr$D_IN = RTL___near_mem___dcache___req_addr ; 
  assign  RTL___near_mem___dcache___rg_addr$EN = RTL___near_mem___dcache___EN_req ; 
    wire[6:0] RTL___near_mem___dcache___MUX_rg_cset_in_cache$write_1__VAL_1_any_val ; 
  assign  RTL___near_mem___dcache___rg_cset_in_cache$D_IN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset  ?  RTL___near_mem___dcache___MUX_rg_cset_in_cache$write_1__VAL_1_any_val :7'd0; 
  assign  RTL___near_mem___dcache___rg_cset_in_cache$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset || RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___rg_error_during_refill$D_IN = RTL___near_mem___dcache___MUX_rg_error_during_refill$write_1__SEL_1 ; 
  assign  RTL___near_mem___dcache___rg_error_during_refill$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill ; 
  always @(      RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_1                  or   RTL___near_mem___dcache___MUX_rg_exc_code$write_1__VAL_1             or   RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_2            or   RTL___near_mem___dcache___MUX_rg_error_during_refill$write_1__SEL_1           or   RTL___near_mem___dcache___access_exc_code__h2256  )
         case (1'b1) 
          RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_1  : 
              RTL___near_mem___dcache___rg_exc_code$D_IN  = RTL___near_mem___dcache___MUX_rg_exc_code$write_1__VAL_1 ; 
          RTL___near_mem___dcache___MUX_rg_exc_code$write_1__SEL_2  : 
              RTL___near_mem___dcache___rg_exc_code$D_IN  =4'd5; 
          RTL___near_mem___dcache___MUX_rg_error_during_refill$write_1__SEL_1  : 
              RTL___near_mem___dcache___rg_exc_code$D_IN  = RTL___near_mem___dcache___access_exc_code__h2256 ;
          default : 
              RTL___near_mem___dcache___rg_exc_code$D_IN  =4'b1010;endcase
  assign  RTL___near_mem___dcache___rg_exc_code$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL___near_mem___dcache___rg_f3$D_IN = RTL___near_mem___dcache___req_f3 ; 
  assign  RTL___near_mem___dcache___rg_f3$EN = RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___rg_ld_val$D_IN = RTL___near_mem___dcache___ld_val__h17594 ; 
  assign  RTL___near_mem___dcache___rg_ld_val$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp ; 
  assign  RTL___near_mem___dcache___rg_lower_word32$D_IN =32'h0; 
  assign  RTL___near_mem___dcache___rg_lower_word32$EN =1'b0; 
  assign  RTL___near_mem___dcache___rg_lower_word32_full$D_IN =1'd0; 
  assign  RTL___near_mem___dcache___rg_lower_word32_full$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___dcache___rg_op$D_IN = RTL___near_mem___dcache___req_op ; 
  assign  RTL___near_mem___dcache___rg_op$EN = RTL___near_mem___dcache___EN_req ; 
  assign  RTL___near_mem___dcache___rg_pa$D_IN = RTL___near_mem___dcache___EN_req  ?  RTL___near_mem___dcache___req_addr : RTL___near_mem___dcache___rg_addr ; 
  assign  RTL___near_mem___dcache___rg_pa$EN = RTL___near_mem___dcache___EN_req || RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp ; 
  assign  RTL___near_mem___dcache___rg_pte_pa$D_IN =32'h0; 
  assign  RTL___near_mem___dcache___rg_pte_pa$EN =1'b0; 
  assign  RTL___near_mem___dcache___rg_st_amo_val$D_IN = RTL___near_mem___dcache___req_st_value ; 
  assign  RTL___near_mem___dcache___rg_st_amo_val$EN = RTL___near_mem___dcache___EN_req ; 
  always @(               RTL___near_mem___dcache___EN_req                                    or   RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_1                      or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset                     or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req                    or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp                   or   RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_4                  or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req                 or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq                or   RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_7               or   RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_7              or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill             or   RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_9            or   RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_9           or   RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_10  )
         case (1'b1) 
          RTL___near_mem___dcache___EN_req  : 
              RTL___near_mem___dcache___rg_state$D_IN  = RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_1 ; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd1; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd11; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp  : 
              RTL___near_mem___dcache___rg_state$D_IN  = RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_4 ; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd13; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd3; 
          RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_7  : 
              RTL___near_mem___dcache___rg_state$D_IN  = RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_7 ; 
          RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd9; 
          RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_9  : 
              RTL___near_mem___dcache___rg_state$D_IN  = RTL___near_mem___dcache___MUX_rg_state$write_1__VAL_9 ; 
          RTL___near_mem___dcache___MUX_rg_state$write_1__SEL_10  : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'd2;
          default : 
              RTL___near_mem___dcache___rg_state$D_IN  =4'b1010;endcase
  assign  RTL___near_mem___dcache___rg_state$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]==2'd3|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 || RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp || RTL___near_mem___dcache___EN_req || RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset || RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq || RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req || RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL___near_mem___dcache___rg_word64_set_in_cache$D_IN = RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2  ?  RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_2 : RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_4 ; 
  assign  RTL___near_mem___dcache___rg_word64_set_in_cache$EN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]!=2'd3|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs$D_IN = RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__SEL_1  ?  RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_1 : RTL___near_mem___dcache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs$ENQ = RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op || RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs$DEQ = RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___dcache___f_fabric_write_reqs$CLR =1'b0; 
  assign  RTL___near_mem___dcache___f_reset_reqs$D_IN =! RTL___near_mem___dcache___EN_server_reset_request_put ; 
  assign  RTL___near_mem___dcache___f_reset_reqs$ENQ = RTL___near_mem___dcache___EN_server_reset_request_put || RTL___near_mem___dcache___EN_server_flush_request_put ; 
  assign  RTL___near_mem___dcache___f_reset_reqs$DEQ = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127; 
  assign  RTL___near_mem___dcache___f_reset_reqs$CLR =1'b0; 
  assign  RTL___near_mem___dcache___f_reset_rsps$D_IN = RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___f_reset_rsps$ENQ = RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127; 
  assign  RTL___near_mem___dcache___f_reset_rsps$DEQ = RTL___near_mem___dcache___EN_server_flush_response_get || RTL___near_mem___dcache___EN_server_reset_response_get ; 
  assign  RTL___near_mem___dcache___f_reset_rsps$CLR =1'b0; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr$D_IN = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 : RTL___near_mem___dcache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr$ENQ = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr$DEQ = RTL___near_mem___dcache___master_xactor_f_rd_addr$EMPTY_N && RTL___near_mem___dcache___mem_master_arready ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_addr$CLR = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data$D_IN ={ RTL___near_mem___dcache___mem_master_rid , RTL___near_mem___dcache___mem_master_rdata , RTL___near_mem___dcache___mem_master_rresp , RTL___near_mem___dcache___mem_master_rlast }; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data$ENQ = RTL___near_mem___dcache___mem_master_rvalid && RTL___near_mem___dcache___master_xactor_f_rd_data$FULL_N ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data$DEQ = RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp || RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop ; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_data$CLR = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr$D_IN ={4'd0, RTL___near_mem___dcache___mem_req_wr_addr_awaddr__h2473 ,8'd0, RTL___near_mem___dcache___x__h2520 ,18'd65536}; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr$ENQ = RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr$DEQ = RTL___near_mem___dcache___master_xactor_f_wr_addr$EMPTY_N && RTL___near_mem___dcache___mem_master_awready ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_addr$CLR = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data$D_IN ={ RTL___near_mem___dcache___mem_req_wr_data_wdata__h2699 , RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700 ,1'd1}; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data$ENQ = RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data$DEQ = RTL___near_mem___dcache___master_xactor_f_wr_data$EMPTY_N && RTL___near_mem___dcache___mem_master_wready ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_data$CLR = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp$D_IN ={ RTL___near_mem___dcache___mem_master_bid , RTL___near_mem___dcache___mem_master_bresp }; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp$ENQ = RTL___near_mem___dcache___mem_master_bvalid && RTL___near_mem___dcache___master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp$DEQ = RTL___near_mem___dcache___CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL___near_mem___dcache___master_xactor_f_wr_resp$CLR = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___dcache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRA = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___dcache___rg_addr [11:5]: RTL___near_mem___dcache___rg_cset_in_cache ; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRB = RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ?  RTL___near_mem___dcache___req_addr [11:5]: RTL___near_mem___dcache___rg_addr [11:5]; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$DIA = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 :23'd2796202; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$DIB = RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ? 23'b01010101010101010101010:23'b01010101010101010101010; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$WEA =1'd1; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$WEB =1'd0; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$ENA = RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset ; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset$ENB = RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq ; 
  assign  RTL___near_mem___dcache___ram_word64_set$ADDRA = RTL___near_mem___dcache___MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL___near_mem___dcache___rg_word64_set_in_cache : RTL___near_mem___dcache___rg_addr [11:3]; 
  always @(         RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                        or   RTL___near_mem___dcache___req_addr                or   RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2               or   RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_2              or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq             or   RTL___near_mem___dcache___rg_addr            or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill           or   RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_4  )
         begin 
             case (1'b1) 
              RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL___near_mem___dcache___ram_word64_set$ADDRB  = RTL___near_mem___dcache___req_addr [11:3]; 
              RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL___near_mem___dcache___ram_word64_set$ADDRB  = RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_2 ; 
              RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq  : 
                  RTL___near_mem___dcache___ram_word64_set$ADDRB  = RTL___near_mem___dcache___rg_addr [11:3]; 
              RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL___near_mem___dcache___ram_word64_set$ADDRB  = RTL___near_mem___dcache___MUX_ram_word64_set$b_put_2__VAL_4 ;
              default : 
                  RTL___near_mem___dcache___ram_word64_set$ADDRB  =9'b010101010;endcase
         end
  assign  RTL___near_mem___dcache___ram_word64_set$DIA = RTL___near_mem___dcache___MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:3]: RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 ; 
  always @(     RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                or   RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2            or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq           or   RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  )
         begin 
             case (1'b1) 
              RTL___near_mem___dcache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL___near_mem___dcache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___dcache___MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL___near_mem___dcache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq  : 
                  RTL___near_mem___dcache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL___near_mem___dcache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;
              default : 
                  RTL___near_mem___dcache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL___near_mem___dcache___ram_word64_set$WEA =1'd1; 
  assign  RTL___near_mem___dcache___ram_word64_set$WEB =1'd0; 
  assign  RTL___near_mem___dcache___ram_word64_set$ENA = RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 ; 
  assign  RTL___near_mem___dcache___ram_word64_set$ENB = RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]!=2'd3|| RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq || RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL___near_mem___dcache___soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___dcache___soc_map$m_is_mem_addr_addr ={32'd0, RTL___near_mem___dcache___rg_addr }; 
  assign  RTL___near_mem___dcache___soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 = RTL___near_mem___dcache___cfg_verbosity >4'd1; 
  assign  RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 = RTL___near_mem___dcache___cfg_verbosity >4'd2; 
  assign  RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 =(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___dcache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 =(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&&! RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___dcache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 = RTL___near_mem___dcache___req_f3 [1:0]!=2'b0&&( RTL___near_mem___dcache___req_f3 [1:0]!=2'b01|| RTL___near_mem___dcache___req_addr [0])&&( RTL___near_mem___dcache___req_f3 [1:0]!=2'b10|| RTL___near_mem___dcache___req_addr [1:0]!=2'b0)&&( RTL___near_mem___dcache___req_f3 [1:0]!=2'b11|| RTL___near_mem___dcache___req_addr [2:0]!=3'b0); 
  assign  RTL___near_mem___dcache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 =! RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL___near_mem___dcache____theResult___snd_fst__h2707 = RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [63:0]<< RTL___near_mem___dcache___shift_bits__h2487 ; 
  assign  RTL___near_mem___dcache___access_exc_code__h2256 = RTL___near_mem___dcache___dmem_not_imem  ? ( RTL___near_mem___dcache___rg_op  ? 4'd7:4'd5):4'd1; 
  assign  RTL___near_mem___dcache___b__h14485 = RTL___near_mem___dcache___CAN_FIRE_RL_rl_fabric_send_write_req  ?  RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$port0__write_1 : RTL___near_mem___dcache___ctr_wr_rsps_pending_crg ; 
  assign  RTL___near_mem___dcache___cline_addr__h14583 ={ RTL___near_mem___dcache___rg_pa [31:5],5'd0}; 
  assign  RTL___near_mem___dcache___cline_fabric_addr__h14584 ={32'd0, RTL___near_mem___dcache___cline_addr__h14583 }; 
  assign  RTL___near_mem___dcache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 = RTL___near_mem___dcache___dmem_not_imem &&! RTL___near_mem___dcache___soc_map$m_is_mem_addr || RTL___near_mem___dcache___rg_op ||! RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___dcache___fabric_addr__h17243 ={32'd0, RTL___near_mem___dcache___rg_pa }; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [10:3]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [18:11]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [18:3]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [26:19]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:19]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:27]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:3]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [42:35]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [50:35]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [50:43]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [58:51]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:35]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:51]; 
  assign  RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 = RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:59]; 
  assign  RTL___near_mem___dcache___mem_req_wr_addr_awaddr__h2473 ={32'd0, RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [95:64]}; 
  assign  RTL___near_mem___dcache___pa_ctag__h4952 ={2'd0, RTL___near_mem___dcache___rg_addr [31:12]}; 
  assign  RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 = RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [21:0]== RTL___near_mem___dcache___pa_ctag__h4952 ; 
  assign  RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 = RTL___near_mem___dcache___req_f3 [1:0]==2'b0|| RTL___near_mem___dcache___req_f3 [1:0]==2'b01&&! RTL___near_mem___dcache___req_addr [0]|| RTL___near_mem___dcache___req_f3 [1:0]==2'b10&& RTL___near_mem___dcache___req_addr [1:0]==2'b0|| RTL___near_mem___dcache___req_f3 [1:0]==2'b11&& RTL___near_mem___dcache___req_addr [2:0]==3'b0; 
  assign  RTL___near_mem___dcache___result__h11657 ={{56{ RTL___near_mem___dcache___word64094_BITS_15_TO_8__q18 [7]}}, RTL___near_mem___dcache___word64094_BITS_15_TO_8__q18 }; 
  assign  RTL___near_mem___dcache___result__h11685 ={{56{ RTL___near_mem___dcache___word64094_BITS_23_TO_16__q19 [7]}}, RTL___near_mem___dcache___word64094_BITS_23_TO_16__q19 }; 
  assign  RTL___near_mem___dcache___result__h11713 ={{56{ RTL___near_mem___dcache___word64094_BITS_31_TO_24__q21 [7]}}, RTL___near_mem___dcache___word64094_BITS_31_TO_24__q21 }; 
  assign  RTL___near_mem___dcache___result__h11741 ={{56{ RTL___near_mem___dcache___word64094_BITS_39_TO_32__q22 [7]}}, RTL___near_mem___dcache___word64094_BITS_39_TO_32__q22 }; 
  assign  RTL___near_mem___dcache___result__h11769 ={{56{ RTL___near_mem___dcache___word64094_BITS_47_TO_40__q25 [7]}}, RTL___near_mem___dcache___word64094_BITS_47_TO_40__q25 }; 
  assign  RTL___near_mem___dcache___result__h11797 ={{56{ RTL___near_mem___dcache___word64094_BITS_55_TO_48__q26 [7]}}, RTL___near_mem___dcache___word64094_BITS_55_TO_48__q26 }; 
  assign  RTL___near_mem___dcache___result__h11825 ={{56{ RTL___near_mem___dcache___word64094_BITS_63_TO_56__q28 [7]}}, RTL___near_mem___dcache___word64094_BITS_63_TO_56__q28 }; 
  assign  RTL___near_mem___dcache___result__h11870 ={56'd0, RTL___near_mem___dcache___word64__h5094 [7:0]}; 
  assign  RTL___near_mem___dcache___result__h11898 ={56'd0, RTL___near_mem___dcache___word64__h5094 [15:8]}; 
  assign  RTL___near_mem___dcache___result__h11926 ={56'd0, RTL___near_mem___dcache___word64__h5094 [23:16]}; 
  assign  RTL___near_mem___dcache___result__h11954 ={56'd0, RTL___near_mem___dcache___word64__h5094 [31:24]}; 
  assign  RTL___near_mem___dcache___result__h11982 ={56'd0, RTL___near_mem___dcache___word64__h5094 [39:32]}; 
  assign  RTL___near_mem___dcache___result__h12010 ={56'd0, RTL___near_mem___dcache___word64__h5094 [47:40]}; 
  assign  RTL___near_mem___dcache___result__h12038 ={56'd0, RTL___near_mem___dcache___word64__h5094 [55:48]}; 
  assign  RTL___near_mem___dcache___result__h12066 ={56'd0, RTL___near_mem___dcache___word64__h5094 [63:56]}; 
  assign  RTL___near_mem___dcache___result__h12111 ={{48{ RTL___near_mem___dcache___word64094_BITS_15_TO_0__q16 [15]}}, RTL___near_mem___dcache___word64094_BITS_15_TO_0__q16 }; 
  assign  RTL___near_mem___dcache___result__h12139 ={{48{ RTL___near_mem___dcache___word64094_BITS_31_TO_16__q20 [15]}}, RTL___near_mem___dcache___word64094_BITS_31_TO_16__q20 }; 
  assign  RTL___near_mem___dcache___result__h12167 ={{48{ RTL___near_mem___dcache___word64094_BITS_47_TO_32__q23 [15]}}, RTL___near_mem___dcache___word64094_BITS_47_TO_32__q23 }; 
  assign  RTL___near_mem___dcache___result__h12195 ={{48{ RTL___near_mem___dcache___word64094_BITS_63_TO_48__q27 [15]}}, RTL___near_mem___dcache___word64094_BITS_63_TO_48__q27 }; 
  assign  RTL___near_mem___dcache___result__h12236 ={48'd0, RTL___near_mem___dcache___word64__h5094 [15:0]}; 
  assign  RTL___near_mem___dcache___result__h12264 ={48'd0, RTL___near_mem___dcache___word64__h5094 [31:16]}; 
  assign  RTL___near_mem___dcache___result__h12292 ={48'd0, RTL___near_mem___dcache___word64__h5094 [47:32]}; 
  assign  RTL___near_mem___dcache___result__h12320 ={48'd0, RTL___near_mem___dcache___word64__h5094 [63:48]}; 
  assign  RTL___near_mem___dcache___result__h12361 ={{32{ RTL___near_mem___dcache___word64094_BITS_31_TO_0__q17 [31]}}, RTL___near_mem___dcache___word64094_BITS_31_TO_0__q17 }; 
  assign  RTL___near_mem___dcache___result__h12389 ={{32{ RTL___near_mem___dcache___word64094_BITS_63_TO_32__q24 [31]}}, RTL___near_mem___dcache___word64094_BITS_63_TO_32__q24 }; 
  assign  RTL___near_mem___dcache___result__h12428 ={32'd0, RTL___near_mem___dcache___word64__h5094 [31:0]}; 
  assign  RTL___near_mem___dcache___result__h12456 ={32'd0, RTL___near_mem___dcache___word64__h5094 [63:32]}; 
  assign  RTL___near_mem___dcache___result__h17654 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 }; 
  assign  RTL___near_mem___dcache___result__h17684 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 }; 
  assign  RTL___near_mem___dcache___result__h17711 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 }; 
  assign  RTL___near_mem___dcache___result__h17738 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 }; 
  assign  RTL___near_mem___dcache___result__h17765 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 }; 
  assign  RTL___near_mem___dcache___result__h17792 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 }; 
  assign  RTL___near_mem___dcache___result__h17819 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 }; 
  assign  RTL___near_mem___dcache___result__h17846 ={{56{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 [7]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 }; 
  assign  RTL___near_mem___dcache___result__h17890 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [10:3]}; 
  assign  RTL___near_mem___dcache___result__h17917 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [18:11]}; 
  assign  RTL___near_mem___dcache___result__h17944 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [26:19]}; 
  assign  RTL___near_mem___dcache___result__h17971 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:27]}; 
  assign  RTL___near_mem___dcache___result__h17998 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [42:35]}; 
  assign  RTL___near_mem___dcache___result__h18025 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [50:43]}; 
  assign  RTL___near_mem___dcache___result__h18052 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [58:51]}; 
  assign  RTL___near_mem___dcache___result__h18079 ={56'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:59]}; 
  assign  RTL___near_mem___dcache___result__h18123 ={{48{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 [15]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 }; 
  assign  RTL___near_mem___dcache___result__h18150 ={{48{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 [15]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 }; 
  assign  RTL___near_mem___dcache___result__h18177 ={{48{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 [15]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 }; 
  assign  RTL___near_mem___dcache___result__h18204 ={{48{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 [15]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 }; 
  assign  RTL___near_mem___dcache___result__h18244 ={48'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [18:3]}; 
  assign  RTL___near_mem___dcache___result__h18271 ={48'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:19]}; 
  assign  RTL___near_mem___dcache___result__h18298 ={48'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [50:35]}; 
  assign  RTL___near_mem___dcache___result__h18325 ={48'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:51]}; 
  assign  RTL___near_mem___dcache___result__h18365 ={{32{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 [31]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 }; 
  assign  RTL___near_mem___dcache___result__h18392 ={{32{ RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 [31]}}, RTL___near_mem___dcache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 }; 
  assign  RTL___near_mem___dcache___result__h18430 ={32'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [34:3]}; 
  assign  RTL___near_mem___dcache___result__h18457 ={32'd0, RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:35]}; 
  assign  RTL___near_mem___dcache___result__h5301 ={{56{ RTL___near_mem___dcache___word64094_BITS_7_TO_0__q15 [7]}}, RTL___near_mem___dcache___word64094_BITS_7_TO_0__q15 }; 
  assign  RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 = RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL___near_mem___dcache___shift_bits__h2487 ={ RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [66:64],3'b0}; 
  assign  RTL___near_mem___dcache___strobe64__h2637 =8'b00000001<< RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___dcache___strobe64__h2639 =8'b00000011<< RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___dcache___strobe64__h2641 =8'b00001111<< RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___dcache___word64094_BITS_15_TO_0__q16 = RTL___near_mem___dcache___word64__h5094 [15:0]; 
  assign  RTL___near_mem___dcache___word64094_BITS_15_TO_8__q18 = RTL___near_mem___dcache___word64__h5094 [15:8]; 
  assign  RTL___near_mem___dcache___word64094_BITS_23_TO_16__q19 = RTL___near_mem___dcache___word64__h5094 [23:16]; 
  assign  RTL___near_mem___dcache___word64094_BITS_31_TO_0__q17 = RTL___near_mem___dcache___word64__h5094 [31:0]; 
  assign  RTL___near_mem___dcache___word64094_BITS_31_TO_16__q20 = RTL___near_mem___dcache___word64__h5094 [31:16]; 
  assign  RTL___near_mem___dcache___word64094_BITS_31_TO_24__q21 = RTL___near_mem___dcache___word64__h5094 [31:24]; 
  assign  RTL___near_mem___dcache___word64094_BITS_39_TO_32__q22 = RTL___near_mem___dcache___word64__h5094 [39:32]; 
  assign  RTL___near_mem___dcache___word64094_BITS_47_TO_32__q23 = RTL___near_mem___dcache___word64__h5094 [47:32]; 
  assign  RTL___near_mem___dcache___word64094_BITS_47_TO_40__q25 = RTL___near_mem___dcache___word64__h5094 [47:40]; 
  assign  RTL___near_mem___dcache___word64094_BITS_55_TO_48__q26 = RTL___near_mem___dcache___word64__h5094 [55:48]; 
  assign  RTL___near_mem___dcache___word64094_BITS_63_TO_32__q24 = RTL___near_mem___dcache___word64__h5094 [63:32]; 
  assign  RTL___near_mem___dcache___word64094_BITS_63_TO_48__q27 = RTL___near_mem___dcache___word64__h5094 [63:48]; 
  assign  RTL___near_mem___dcache___word64094_BITS_63_TO_56__q28 = RTL___near_mem___dcache___word64__h5094 [63:56]; 
  assign  RTL___near_mem___dcache___word64094_BITS_7_TO_0__q15 = RTL___near_mem___dcache___word64__h5094 [7:0]; 
  assign  RTL___near_mem___dcache___word64__h5094 = RTL___near_mem___dcache___ram_word64_set$DOB & RTL___near_mem___dcache___y__h5337 ; 
  assign  RTL___near_mem___dcache___y__h5337 ={64{ RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 }}; 
  always @(  RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT  )
         begin 
             case ( RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL___near_mem___dcache___x__h2520  =3'b0;
              2 'b01: 
                  RTL___near_mem___dcache___x__h2520  =3'b001;
              2 'b10: 
                  RTL___near_mem___dcache___x__h2520  =3'b010;
              2 'b11: 
                  RTL___near_mem___dcache___x__h2520  =3'b011;endcase
         end
  always @(  RTL___near_mem___dcache___rg_f3  )
         begin 
             case ( RTL___near_mem___dcache___rg_f3 [1:0])
              2 'b0: 
                  RTL___near_mem___dcache___value__h17372  =3'b0;
              2 'b01: 
                  RTL___near_mem___dcache___value__h17372  =3'b001;
              2 'b10: 
                  RTL___near_mem___dcache___value__h17372  =3'b010;
              2 'd3: 
                  RTL___near_mem___dcache___value__h17372  =3'b011;endcase
         end
  always @(     RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT                or   RTL___near_mem___dcache___strobe64__h2637            or   RTL___near_mem___dcache___strobe64__h2639           or   RTL___near_mem___dcache___strobe64__h2641  )
         begin 
             case ( RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___dcache___strobe64__h2637 ;
              2 'b01: 
                  RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___dcache___strobe64__h2639 ;
              2 'b10: 
                  RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___dcache___strobe64__h2641 ;
              2 'b11: 
                  RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700  =8'b11111111;endcase
         end
  always @(   RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT            or   RTL___near_mem___dcache____theResult___snd_fst__h2707  )
         begin 
             case ( RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0,2'b01,2'b10: 
                  RTL___near_mem___dcache___mem_req_wr_data_wdata__h2699  = RTL___near_mem___dcache____theResult___snd_fst__h2707 ;
              2 'd3: 
                  RTL___near_mem___dcache___mem_req_wr_data_wdata__h2699  = RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT [63:0];endcase
         end
  always @(      RTL___near_mem___dcache___rg_addr                  or   RTL___near_mem___dcache___result__h12111             or   RTL___near_mem___dcache___result__h12139            or   RTL___near_mem___dcache___result__h12167           or   RTL___near_mem___dcache___result__h12195  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___dcache___result__h12111 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___dcache___result__h12139 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___dcache___result__h12167 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___dcache___result__h12195 ;
              default : 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  =64'd0;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___ram_word64_set$DOB           or   RTL___near_mem___dcache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:16], RTL___near_mem___dcache___rg_st_amo_val [15:0]};
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:32], RTL___near_mem___dcache___rg_st_amo_val [15:0], RTL___near_mem___dcache___ram_word64_set$DOB [15:0]};
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:48], RTL___near_mem___dcache___rg_st_amo_val [15:0], RTL___near_mem___dcache___ram_word64_set$DOB [31:0]};
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___dcache___rg_st_amo_val [15:0], RTL___near_mem___dcache___ram_word64_set$DOB [47:0]};
              default : 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  = RTL___near_mem___dcache___ram_word64_set$DOB ;endcase
         end
  always @(          RTL___near_mem___dcache___rg_addr                          or   RTL___near_mem___dcache___result__h5301                 or   RTL___near_mem___dcache___result__h11657                or   RTL___near_mem___dcache___result__h11685               or   RTL___near_mem___dcache___result__h11713              or   RTL___near_mem___dcache___result__h11741             or   RTL___near_mem___dcache___result__h11769            or   RTL___near_mem___dcache___result__h11797           or   RTL___near_mem___dcache___result__h11825  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h5301 ;
              3 'h1: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11657 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11685 ;
              3 'h3: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11713 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11741 ;
              3 'h5: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11769 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11797 ;
              3 'h7: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___dcache___result__h11825 ;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___ram_word64_set$DOB           or   RTL___near_mem___dcache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:8], RTL___near_mem___dcache___rg_st_amo_val [7:0]};
              3 'h1: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:16], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [7:0]};
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:24], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [15:0]};
              3 'h3: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:32], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [23:0]};
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:40], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [31:0]};
              3 'h5: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:48], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [39:0]};
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:56], RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [47:0]};
              3 'h7: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___dcache___rg_st_amo_val [7:0], RTL___near_mem___dcache___ram_word64_set$DOB [55:0]};endcase
         end
  always @(      RTL___near_mem___dcache___rg_addr                  or   RTL___near_mem___dcache___result__h18244             or   RTL___near_mem___dcache___result__h18271            or   RTL___near_mem___dcache___result__h18298           or   RTL___near_mem___dcache___result__h18325  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___dcache___result__h18244 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___dcache___result__h18271 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___dcache___result__h18298 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___dcache___result__h18325 ;
              default : 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  =64'd0;endcase
         end
  always @(      RTL___near_mem___dcache___rg_addr                  or   RTL___near_mem___dcache___result__h12236             or   RTL___near_mem___dcache___result__h12264            or   RTL___near_mem___dcache___result__h12292           or   RTL___near_mem___dcache___result__h12320  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___dcache___result__h12236 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___dcache___result__h12264 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___dcache___result__h12292 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___dcache___result__h12320 ;
              default : 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  =64'd0;endcase
         end
  always @(      RTL___near_mem___dcache___rg_addr                  or   RTL___near_mem___dcache___result__h18123             or   RTL___near_mem___dcache___result__h18150            or   RTL___near_mem___dcache___result__h18177           or   RTL___near_mem___dcache___result__h18204  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___dcache___result__h18123 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___dcache___result__h18150 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___dcache___result__h18177 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___dcache___result__h18204 ;
              default : 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  =64'd0;endcase
         end
  always @(          RTL___near_mem___dcache___rg_addr                          or   RTL___near_mem___dcache___result__h17890                 or   RTL___near_mem___dcache___result__h17917                or   RTL___near_mem___dcache___result__h17944               or   RTL___near_mem___dcache___result__h17971              or   RTL___near_mem___dcache___result__h17998             or   RTL___near_mem___dcache___result__h18025            or   RTL___near_mem___dcache___result__h18052           or   RTL___near_mem___dcache___result__h18079  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h17890 ;
              3 'h1: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h17917 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h17944 ;
              3 'h3: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h17971 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h17998 ;
              3 'h5: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h18025 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h18052 ;
              3 'h7: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___dcache___result__h18079 ;endcase
         end
  always @(          RTL___near_mem___dcache___rg_addr                          or   RTL___near_mem___dcache___result__h11870                 or   RTL___near_mem___dcache___result__h11898                or   RTL___near_mem___dcache___result__h11926               or   RTL___near_mem___dcache___result__h11954              or   RTL___near_mem___dcache___result__h11982             or   RTL___near_mem___dcache___result__h12010            or   RTL___near_mem___dcache___result__h12038           or   RTL___near_mem___dcache___result__h12066  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h11870 ;
              3 'h1: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h11898 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h11926 ;
              3 'h3: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h11954 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h11982 ;
              3 'h5: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h12010 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h12038 ;
              3 'h7: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___dcache___result__h12066 ;endcase
         end
  always @(          RTL___near_mem___dcache___rg_addr                          or   RTL___near_mem___dcache___result__h17654                 or   RTL___near_mem___dcache___result__h17684                or   RTL___near_mem___dcache___result__h17711               or   RTL___near_mem___dcache___result__h17738              or   RTL___near_mem___dcache___result__h17765             or   RTL___near_mem___dcache___result__h17792            or   RTL___near_mem___dcache___result__h17819           or   RTL___near_mem___dcache___result__h17846  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17654 ;
              3 'h1: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17684 ;
              3 'h2: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17711 ;
              3 'h3: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17738 ;
              3 'h4: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17765 ;
              3 'h5: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17792 ;
              3 'h6: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17819 ;
              3 'h7: 
                  RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___dcache___result__h17846 ;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___result__h18365           or   RTL___near_mem___dcache___result__h18392  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL___near_mem___dcache___result__h18365 ;
              3 'h4: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL___near_mem___dcache___result__h18392 ;
              default : 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  =64'd0;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___result__h18430           or   RTL___near_mem___dcache___result__h18457  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL___near_mem___dcache___result__h18430 ;
              3 'h4: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL___near_mem___dcache___result__h18457 ;
              default : 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  =64'd0;endcase
         end
  always @(          RTL___near_mem___dcache___rg_f3                          or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411                 or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439                or   RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29               or   RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT             or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427            or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447           or   RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  )
         begin 
             case ( RTL___near_mem___dcache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 ;
              3 'b001: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 ;
              3 'b010: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 ;
              3 'b011: 
                  RTL___near_mem___dcache___ld_val__h17594  =( RTL___near_mem___dcache___rg_addr [2:0]==3'h0) ?  RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:3]:64'd0;
              3 'b100: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 ;
              3 'b101: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 ;
              3 'b110: 
                  RTL___near_mem___dcache___ld_val__h17594  = RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 ;
              3 'd7: 
                  RTL___near_mem___dcache___ld_val__h17594  =64'd0;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___ram_word64_set$DOB           or   RTL___near_mem___dcache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL___near_mem___dcache___ram_word64_set$DOB [63:32], RTL___near_mem___dcache___rg_st_amo_val [31:0]};
              3 'h4: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL___near_mem___dcache___rg_st_amo_val [31:0], RTL___near_mem___dcache___ram_word64_set$DOB [31:0]};
              default : 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  = RTL___near_mem___dcache___ram_word64_set$DOB ;endcase
         end
  always @(       RTL___near_mem___dcache___rg_f3                    or   RTL___near_mem___dcache___ram_word64_set$DOB              or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157             or   RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167            or   RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31           or   RTL___near_mem___dcache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___dcache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 ;
              3 'b001: 
                  RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___dcache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 ;
              3 'b010: 
                  RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 ;
              3 'b011: 
                  RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___dcache___rg_st_amo_val ;
              default : 
                  RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___dcache___ram_word64_set$DOB ;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___result__h12361           or   RTL___near_mem___dcache___result__h12389  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL___near_mem___dcache___result__h12361 ;
              3 'h4: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL___near_mem___dcache___result__h12389 ;
              default : 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  =64'd0;endcase
         end
  always @(    RTL___near_mem___dcache___rg_addr              or   RTL___near_mem___dcache___result__h12428           or   RTL___near_mem___dcache___result__h12456  )
         begin 
             case ( RTL___near_mem___dcache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL___near_mem___dcache___result__h12428 ;
              3 'h4: 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL___near_mem___dcache___result__h12456 ;
              default : 
                  RTL___near_mem___dcache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  =64'd0;endcase
         end
  always @( posedge  RTL___near_mem___dcache___CLK )
         begin 
             if ( RTL___near_mem___dcache___RST_N ==1'b0)
                 begin  
                     RTL___near_mem___dcache___cfg_verbosity  <=4'd0; 
                     RTL___near_mem___dcache___ctr_wr_rsps_pending_crg  <=4'd0; 
                     RTL___near_mem___dcache___rg_cset_in_cache  <=7'd0; 
                     RTL___near_mem___dcache___rg_lower_word32_full  <=1'd0; 
                     RTL___near_mem___dcache___rg_state  <=4'd0;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___dcache___cfg_verbosity$EN ) 
                         RTL___near_mem___dcache___cfg_verbosity  <= RTL___near_mem___dcache___cfg_verbosity$D_IN ;
                     if ( RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$EN ) 
                         RTL___near_mem___dcache___ctr_wr_rsps_pending_crg  <= RTL___near_mem___dcache___ctr_wr_rsps_pending_crg$D_IN ;
                     if ( RTL___near_mem___dcache___rg_cset_in_cache$EN ) 
                         RTL___near_mem___dcache___rg_cset_in_cache  <= RTL___near_mem___dcache___rg_cset_in_cache$D_IN ;
                     if ( RTL___near_mem___dcache___rg_lower_word32_full$EN ) 
                         RTL___near_mem___dcache___rg_lower_word32_full  <= RTL___near_mem___dcache___rg_lower_word32_full$D_IN ;
                     if ( RTL___near_mem___dcache___rg_state$EN ) 
                         RTL___near_mem___dcache___rg_state  <= RTL___near_mem___dcache___rg_state$D_IN ;
                 end 
             if ( RTL___near_mem___dcache___rg_addr$EN ) 
                 RTL___near_mem___dcache___rg_addr  <= RTL___near_mem___dcache___rg_addr$D_IN ;
             if ( RTL___near_mem___dcache___rg_error_during_refill$EN ) 
                 RTL___near_mem___dcache___rg_error_during_refill  <= RTL___near_mem___dcache___rg_error_during_refill$D_IN ;
             if ( RTL___near_mem___dcache___rg_exc_code$EN ) 
                 RTL___near_mem___dcache___rg_exc_code  <= RTL___near_mem___dcache___rg_exc_code$D_IN ;
             if ( RTL___near_mem___dcache___rg_f3$EN ) 
                 RTL___near_mem___dcache___rg_f3  <= RTL___near_mem___dcache___rg_f3$D_IN ;
             if ( RTL___near_mem___dcache___rg_ld_val$EN ) 
                 RTL___near_mem___dcache___rg_ld_val  <= RTL___near_mem___dcache___rg_ld_val$D_IN ;
             if ( RTL___near_mem___dcache___rg_lower_word32$EN ) 
                 RTL___near_mem___dcache___rg_lower_word32  <= RTL___near_mem___dcache___rg_lower_word32$D_IN ;
             if ( RTL___near_mem___dcache___rg_op$EN ) 
                 RTL___near_mem___dcache___rg_op  <= RTL___near_mem___dcache___rg_op$D_IN ;
             if ( RTL___near_mem___dcache___rg_pa$EN ) 
                 RTL___near_mem___dcache___rg_pa  <= RTL___near_mem___dcache___rg_pa$D_IN ;
             if ( RTL___near_mem___dcache___rg_pte_pa$EN ) 
                 RTL___near_mem___dcache___rg_pte_pa  <= RTL___near_mem___dcache___rg_pte_pa$D_IN ;
             if ( RTL___near_mem___dcache___rg_st_amo_val$EN ) 
                 RTL___near_mem___dcache___rg_st_amo_val  <= RTL___near_mem___dcache___rg_st_amo_val$D_IN ;
             if ( RTL___near_mem___dcache___rg_word64_set_in_cache$EN ) 
                 RTL___near_mem___dcache___rg_word64_set_in_cache  <= RTL___near_mem___dcache___rg_word64_set_in_cache$D_IN ;
         end
  always @( negedge  RTL___near_mem___dcache___CLK )
         begin #0;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___ctr_wr_rsps_pending_crg ==4'd15)
                     begin  
                         RTL___near_mem___dcache___v__h2948  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h2942  = RTL___near_mem___dcache___v__h2948 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___ctr_wr_rsps_pending_crg ==4'd15)$display("%0d: ERROR: CreditCounter: overflow", RTL___near_mem___dcache___v__h2942 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___ctr_wr_rsps_pending_crg ==4'd15)$finish(32'd1);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Addr { ","awid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awaddr: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___mem_req_wr_addr_awaddr__h2473 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlen: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awsize: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___x__h2520 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awburst: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlock: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awcache: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awprot: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awqos: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awregion: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awuser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("                       ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Data { ","wdata: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___mem_req_wr_data_wdata__h2699 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wstrb: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___mem_req_wr_data_wstrb__h2700 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wlast: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("True");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wuser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127&& RTL___near_mem___dcache___cfg_verbosity !=4'd0&&! RTL___near_mem___dcache___f_reset_reqs$D_OUT )
                     begin  
                         RTL___near_mem___dcache___v__h3848  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h3842  = RTL___near_mem___dcache___v__h3848 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127&& RTL___near_mem___dcache___cfg_verbosity !=4'd0&&! RTL___near_mem___dcache___f_reset_reqs$D_OUT )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL___near_mem___dcache___v__h3842 ,"D_MMU_Cache",$signed(32'd128),$signed(32'd1));
                      else $display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL___near_mem___dcache___v__h3842 ,"I_MMU_Cache",$signed(32'd128),$signed(32'd1));
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___f_reset_reqs$D_OUT )
                     begin  
                         RTL___near_mem___dcache___v__h3949  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h3943  = RTL___near_mem___dcache___v__h3949 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_reset && RTL___near_mem___dcache___rg_cset_in_cache ==7'd127&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___f_reset_reqs$D_OUT )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_reset: Flushed", RTL___near_mem___dcache___v__h3943 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_reset: Flushed", RTL___near_mem___dcache___v__h3943 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h4098  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h4092  = RTL___near_mem___dcache___v__h4098 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL___near_mem___dcache___v__h4092 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_addr );
                      else $display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL___near_mem___dcache___v__h4092 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_addr );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        eaddr = {CTag 0x%0h  CSet 0x%0h  Word64 0x%0h  Byte 0x%0h}", RTL___near_mem___dcache___pa_ctag__h4952 , RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_addr [4:3], RTL___near_mem___dcache___rg_addr [2:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x: (state, tag):", RTL___near_mem___dcache___rg_addr [11:5]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" (");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22])$write("CTAG_CLEAN");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22])$write("CTAG_EMPTY");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22])$write(", 0x%0x", RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [21:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22])$write(", --");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(")");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_addr [4:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" 0x%0x", RTL___near_mem___dcache___ram_word64_set$DOB );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    TLB result: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_Xlate_Result { ","outcome: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_XLATE_OK");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","pa: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___rg_addr );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","exc_code: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'hA," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___dcache___dmem_not_imem &&! RTL___near_mem___dcache___soc_map$m_is_mem_addr && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => IO_REQ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$display("        Write-Cache-Hit: pa 0x%0h word64 0x%0h", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_st_amo_val );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        New Word64_Set:");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_addr [4:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write(" 0x%0x", RTL___near_mem___dcache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op &&(! RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Miss: pa 0x%0h word64 0x%0h", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_st_amo_val );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Hit/Miss: eaddr 0x%0h word64 0x%0h", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_st_amo_val );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___rg_op && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        => rl_write_response");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     begin  
                         RTL___near_mem___dcache___v__h12540  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h12534  = RTL___near_mem___dcache___v__h12540 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL___near_mem___dcache___v__h12534 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___word64__h5094 ,64'd0);
                      else $display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL___near_mem___dcache___v__h12534 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___word64__h5094 ,64'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&& RTL___near_mem___dcache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )$display("        Read-hit: addr 0x%0h word64 0x%0h", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___word64__h5094 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___dcache___dmem_not_imem || RTL___near_mem___dcache___soc_map$m_is_mem_addr )&&! RTL___near_mem___dcache___rg_op &&(! RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___dcache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Read Miss: -> CACHE_START_REFILL.");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h14531  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h14525  = RTL___near_mem___dcache___v__h14531 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_start_cache_refill: ", RTL___near_mem___dcache___v__h14525 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_cache_refill: ", RTL___near_mem___dcache___v__h14525 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    To fabric: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___cline_fabric_addr__h14584 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd3);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'b011);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    Victim way %0d; => CACHE_REFILL",1'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     begin  
                         RTL___near_mem___dcache___v__h15336  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h15330  = RTL___near_mem___dcache___v__h15336 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop:", RTL___near_mem___dcache___v__h15330 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_cache_refill_rsps_loop:", RTL___near_mem___dcache___v__h15330 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rdata: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rresp: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rlast: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 &&! RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","ruser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h15578  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h15572  = RTL___near_mem___dcache___v__h15578 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL___near_mem___dcache___v__h15572 ,"D_MMU_Cache", RTL___near_mem___dcache___access_exc_code__h2256 );
                      else $display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL___near_mem___dcache___v__h15572 ,"I_MMU_Cache", RTL___near_mem___dcache___access_exc_code__h2256 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]==2'd3&&( RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___dcache___rg_error_during_refill )&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => MODULE_EXCEPTION_RSP");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]==2'd3&& RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&&! RTL___near_mem___dcache___rg_error_during_refill && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => CACHE_REREQ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$display("        Updating Cache word64_set 0x%0h, word64_in_cline %0d) old => new", RTL___near_mem___dcache___rg_word64_set_in_cache , RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL___near_mem___dcache___ram_word64_set$DOB );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_rereq && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL___near_mem___dcache___rg_addr [11:5], RTL___near_mem___dcache___rg_addr [11:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h17191  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h17185  = RTL___near_mem___dcache___v__h17191 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL___near_mem___dcache___v__h17185 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa );
                      else $display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL___near_mem___dcache___v__h17185 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___fabric_addr__h17243 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___value__h17372 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h17485  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h17479  = RTL___near_mem___dcache___v__h17485 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL___near_mem___dcache___v__h17479 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa );
                      else $display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL___near_mem___dcache___v__h17479 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rdata: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rresp: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rlast: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","ruser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h18585  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h18579  = RTL___near_mem___dcache___v__h18585 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___dcache___v__h18579 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___ld_val__h17594 );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___dcache___v__h18579 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___ld_val__h17594 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h18692  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h18686  = RTL___near_mem___dcache___v__h18692 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL___near_mem___dcache___v__h18686 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL___near_mem___dcache___v__h18686 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h18797  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h18791  = RTL___near_mem___dcache___v__h18797 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___dcache___v__h18791 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_ld_val );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___dcache___v__h18791 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_ld_val );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h18877  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h18871  = RTL___near_mem___dcache___v__h18877 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL___near_mem___dcache___v__h18871 ,"D_MMU_Cache", RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa , RTL___near_mem___dcache___rg_st_amo_val );
                      else $display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL___near_mem___dcache___v__h18871 ,"I_MMU_Cache", RTL___near_mem___dcache___rg_f3 , RTL___near_mem___dcache___rg_addr , RTL___near_mem___dcache___rg_pa , RTL___near_mem___dcache___rg_st_amo_val );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => rl_ST_AMO_response");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h19505  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h19499  = RTL___near_mem___dcache___v__h19505 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL___near_mem___dcache___v__h19499 ,"D_MMU_Cache",$unsigned( RTL___near_mem___dcache___b__h14485 ));
                      else $write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL___near_mem___dcache___v__h19499 ,"I_MMU_Cache",$unsigned( RTL___near_mem___dcache___b__h14485 ));
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","bresp: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","buser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     begin  
                         RTL___near_mem___dcache___v__h19466  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h19460  = RTL___near_mem___dcache___v__h19466 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL___near_mem___dcache___v__h19460 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL___near_mem___dcache___v__h19460 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("    ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","bresp: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","buser: ");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h",1'd0," }");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h3483  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h3477  = RTL___near_mem___dcache___v__h3483 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___WILL_FIRE_RL_rl_start_reset && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___dcache___dmem_not_imem )$display("%0d: %s.rl_start_reset", RTL___near_mem___dcache___v__h3477 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_reset", RTL___near_mem___dcache___v__h3477 ,"I_MMU_Cache");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___dcache___v__h19852  =$stime;#0;
                     end  
             RTL___near_mem___dcache___v__h19846  = RTL___near_mem___dcache___v__h19852 /32'd10;
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("%0d: %m.req: op:", RTL___near_mem___dcache___v__h19846 );
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___req_op )$write("CACHE_ST");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___dcache___req_op )$write("CACHE_LD");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" f3:%0d addr:0x%0h st_value:0x%0h", RTL___near_mem___dcache___req_f3 , RTL___near_mem___dcache___req_addr , RTL___near_mem___dcache___req_st_value ,"\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    priv:");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___req_priv ==2'b0)$write("U");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___req_priv ==2'b01)$write("S");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___req_priv ==2'b11)$write("M");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___dcache___req_priv !=2'b0&& RTL___near_mem___dcache___req_priv !=2'b01&& RTL___near_mem___dcache___req_priv !=2'b11)$write("RESERVED");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" sstatus_SUM:%0d mstatus_MXR:%0d satp:0x%0h", RTL___near_mem___dcache___req_sstatus_SUM , RTL___near_mem___dcache___req_mstatus_MXR , RTL___near_mem___dcache___req_satp ,"\n");
             if ( RTL___near_mem___dcache___RST_N !=1'b0)
                 if ( RTL___near_mem___dcache___EN_req && RTL___near_mem___dcache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 && RTL___near_mem___dcache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL___near_mem___dcache___req_addr [11:5], RTL___near_mem___dcache___req_addr [11:3]);
         end
  assign  RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL___near_mem___dcache___rg_addr ; 
  assign  RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL___near_mem___dcache___rg_pa ;
      
    wire RTL___near_mem___f_reset_rsps___RST;
    wire RTL___near_mem___f_reset_rsps___CLK;
    wire RTL___near_mem___f_reset_rsps___ENQ;
    wire RTL___near_mem___f_reset_rsps___CLR;
    wire RTL___near_mem___f_reset_rsps___DEQ;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    wire RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    wire RTL___near_mem___f_reset_rsps___FULL_N;
    wire RTL___near_mem___f_reset_rsps___EMPTY_N;

    reg RTL___near_mem___f_reset_rsps___empty_reg ; 
    reg RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___FULL_N = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___EMPTY_N = RTL___near_mem___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___near_mem___f_reset_rsps___CLK )
         begin 
             if ( RTL___near_mem___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___near_mem___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___near_mem___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___f_reset_rsps___CLR )
                         begin  
                             RTL___near_mem___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___near_mem___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___f_reset_rsps___ENQ &&! RTL___near_mem___f_reset_rsps___DEQ )
                             begin  
                                 RTL___near_mem___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___near_mem___f_reset_rsps___full_reg  <=! RTL___near_mem___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___near_mem___f_reset_rsps___ENQ && RTL___near_mem___f_reset_rsps___DEQ )
                                 begin  
                                     RTL___near_mem___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___near_mem___f_reset_rsps___empty_reg  <=! RTL___near_mem___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___f_reset_rsps___CLK )
         begin : RTL___near_mem___f_reset_rsps___error_checks 
           reg RTL___near_mem___f_reset_rsps___deqerror , RTL___near_mem___f_reset_rsps___enqerror ; 
             RTL___near_mem___f_reset_rsps___deqerror  =0; 
             RTL___near_mem___f_reset_rsps___enqerror  =0;
             if ( RTL___near_mem___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___f_reset_rsps___empty_reg && RTL___near_mem___f_reset_rsps___DEQ )
                         begin  
                             RTL___near_mem___f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___f_reset_rsps___full_reg && RTL___near_mem___f_reset_rsps___ENQ &&(! RTL___near_mem___f_reset_rsps___DEQ || RTL___near_mem___f_reset_rsps___guarded ))
                         begin  
                             RTL___near_mem___f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___empty_reg ;
    assign RTL___near_mem___f_reset_rsps___RST = RTL___near_mem___RST_N;
    assign RTL___near_mem___f_reset_rsps___CLK = RTL___near_mem___CLK;
    assign RTL___near_mem___f_reset_rsps___ENQ = RTL___near_mem___f_reset_rsps$ENQ;
    assign RTL___near_mem___f_reset_rsps___CLR = RTL___near_mem___f_reset_rsps$CLR;
    assign RTL___near_mem___f_reset_rsps___DEQ = RTL___near_mem___f_reset_rsps$DEQ;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___f_reset_rsps$FULL_N = RTL___near_mem___f_reset_rsps___FULL_N;
    assign RTL___near_mem___f_reset_rsps$EMPTY_N = RTL___near_mem___f_reset_rsps___EMPTY_N;
      
    
    reg[63:0] RTL___near_mem___icache___word64 ; 
    wire[63:0] RTL___near_mem___icache___mem_master_araddr , RTL___near_mem___icache___mem_master_awaddr , RTL___near_mem___icache___mem_master_wdata , RTL___near_mem___icache___st_amo_val ; 
    wire[31:0] RTL___near_mem___icache___addr ; 
    wire[7:0] RTL___near_mem___icache___mem_master_arlen , RTL___near_mem___icache___mem_master_awlen , RTL___near_mem___icache___mem_master_wstrb ; 
    wire[3:0] RTL___near_mem___icache___exc_code , RTL___near_mem___icache___mem_master_arcache , RTL___near_mem___icache___mem_master_arid , RTL___near_mem___icache___mem_master_arqos , RTL___near_mem___icache___mem_master_arregion , RTL___near_mem___icache___mem_master_awcache , RTL___near_mem___icache___mem_master_awid , RTL___near_mem___icache___mem_master_awqos , RTL___near_mem___icache___mem_master_awregion ; 
    wire[2:0] RTL___near_mem___icache___mem_master_arprot , RTL___near_mem___icache___mem_master_arsize , RTL___near_mem___icache___mem_master_awprot , RTL___near_mem___icache___mem_master_awsize ; 
    wire[1:0] RTL___near_mem___icache___mem_master_arburst , RTL___near_mem___icache___mem_master_awburst ; 
    wire RTL___near_mem___icache___RDY_server_flush_request_put , RTL___near_mem___icache___RDY_server_flush_response_get , RTL___near_mem___icache___RDY_server_reset_request_put , RTL___near_mem___icache___RDY_server_reset_response_get , RTL___near_mem___icache___RDY_set_verbosity , RTL___near_mem___icache___RDY_tlb_flush , RTL___near_mem___icache___exc , RTL___near_mem___icache___mem_master_arlock , RTL___near_mem___icache___mem_master_arvalid , RTL___near_mem___icache___mem_master_awlock , RTL___near_mem___icache___mem_master_awvalid , RTL___near_mem___icache___mem_master_bready , RTL___near_mem___icache___mem_master_rready , RTL___near_mem___icache___mem_master_wlast , RTL___near_mem___icache___mem_master_wvalid , RTL___near_mem___icache___valid ; 
    wire[3:0] RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port0__write_1 , RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port1__write_1 , RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port2__read , RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port3__read ; 
    wire RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN_port2__write , RTL___near_mem___icache___dw_valid$whas ; reg[3:0] RTL___near_mem___icache___cfg_verbosity ; 
    wire[3:0] RTL___near_mem___icache___cfg_verbosity$D_IN ; 
    wire RTL___near_mem___icache___cfg_verbosity$EN ; reg[3:0] RTL___near_mem___icache___ctr_wr_rsps_pending_crg ; 
    wire[3:0] RTL___near_mem___icache___ctr_wr_rsps_pending_crg$D_IN ; 
    wire RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN ; reg[31:0] RTL___near_mem___icache___rg_addr ; 
    wire[31:0] RTL___near_mem___icache___rg_addr$D_IN ; 
    wire RTL___near_mem___icache___rg_addr$EN ; reg[6:0] RTL___near_mem___icache___rg_cset_in_cache ; 
    wire[6:0] RTL___near_mem___icache___rg_cset_in_cache$D_IN ; 
    wire RTL___near_mem___icache___rg_cset_in_cache$EN ; 
    reg RTL___near_mem___icache___rg_error_during_refill ; 
    wire RTL___near_mem___icache___rg_error_during_refill$D_IN , RTL___near_mem___icache___rg_error_during_refill$EN ; reg[3:0] RTL___near_mem___icache___rg_exc_code ; reg[3:0] RTL___near_mem___icache___rg_exc_code$D_IN ; 
    wire RTL___near_mem___icache___rg_exc_code$EN ; reg[2:0] RTL___near_mem___icache___rg_f3 ; 
    wire[2:0] RTL___near_mem___icache___rg_f3$D_IN ; 
    wire RTL___near_mem___icache___rg_f3$EN ; reg[63:0] RTL___near_mem___icache___rg_ld_val ; 
    wire[63:0] RTL___near_mem___icache___rg_ld_val$D_IN ; 
    wire RTL___near_mem___icache___rg_ld_val$EN ; reg[31:0] RTL___near_mem___icache___rg_lower_word32 ; 
    wire[31:0] RTL___near_mem___icache___rg_lower_word32$D_IN ; 
    wire RTL___near_mem___icache___rg_lower_word32$EN ; 
    reg RTL___near_mem___icache___rg_lower_word32_full ; 
    wire RTL___near_mem___icache___rg_lower_word32_full$D_IN , RTL___near_mem___icache___rg_lower_word32_full$EN ; 
    reg RTL___near_mem___icache___rg_op ; 
    wire RTL___near_mem___icache___rg_op$D_IN , RTL___near_mem___icache___rg_op$EN ; reg[31:0] RTL___near_mem___icache___rg_pa ; 
    wire[31:0] RTL___near_mem___icache___rg_pa$D_IN ; 
    wire RTL___near_mem___icache___rg_pa$EN ; reg[31:0] RTL___near_mem___icache___rg_pte_pa ; 
    wire[31:0] RTL___near_mem___icache___rg_pte_pa$D_IN ; 
    wire RTL___near_mem___icache___rg_pte_pa$EN ; reg[63:0] RTL___near_mem___icache___rg_st_amo_val ; 
    wire[63:0] RTL___near_mem___icache___rg_st_amo_val$D_IN ; 
    wire RTL___near_mem___icache___rg_st_amo_val$EN ; reg[3:0] RTL___near_mem___icache___rg_state ; reg[3:0] RTL___near_mem___icache___rg_state$D_IN ; 
    wire RTL___near_mem___icache___rg_state$EN ; reg[8:0] RTL___near_mem___icache___rg_word64_set_in_cache ; 
    wire[8:0] RTL___near_mem___icache___rg_word64_set_in_cache$D_IN ; 
    wire RTL___near_mem___icache___rg_word64_set_in_cache$EN ; 
    wire[98:0] RTL___near_mem___icache___f_fabric_write_reqs$D_IN , RTL___near_mem___icache___f_fabric_write_reqs$D_OUT ; 
    wire RTL___near_mem___icache___f_fabric_write_reqs$CLR , RTL___near_mem___icache___f_fabric_write_reqs$DEQ , RTL___near_mem___icache___f_fabric_write_reqs$EMPTY_N , RTL___near_mem___icache___f_fabric_write_reqs$ENQ , RTL___near_mem___icache___f_fabric_write_reqs$FULL_N ; 
    wire RTL___near_mem___icache___f_reset_reqs$CLR , RTL___near_mem___icache___f_reset_reqs$DEQ , RTL___near_mem___icache___f_reset_reqs$D_IN , RTL___near_mem___icache___f_reset_reqs$D_OUT , RTL___near_mem___icache___f_reset_reqs$EMPTY_N , RTL___near_mem___icache___f_reset_reqs$ENQ , RTL___near_mem___icache___f_reset_reqs$FULL_N ; 
    wire RTL___near_mem___icache___f_reset_rsps$CLR , RTL___near_mem___icache___f_reset_rsps$DEQ , RTL___near_mem___icache___f_reset_rsps$D_IN , RTL___near_mem___icache___f_reset_rsps$D_OUT , RTL___near_mem___icache___f_reset_rsps$EMPTY_N , RTL___near_mem___icache___f_reset_rsps$ENQ , RTL___near_mem___icache___f_reset_rsps$FULL_N ; 
    wire[96:0] RTL___near_mem___icache___master_xactor_f_rd_addr$D_IN , RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_addr$CLR , RTL___near_mem___icache___master_xactor_f_rd_addr$DEQ , RTL___near_mem___icache___master_xactor_f_rd_addr$EMPTY_N , RTL___near_mem___icache___master_xactor_f_rd_addr$ENQ , RTL___near_mem___icache___master_xactor_f_rd_addr$FULL_N ; 
    wire[70:0] RTL___near_mem___icache___master_xactor_f_rd_data$D_IN , RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_data$CLR , RTL___near_mem___icache___master_xactor_f_rd_data$DEQ , RTL___near_mem___icache___master_xactor_f_rd_data$EMPTY_N , RTL___near_mem___icache___master_xactor_f_rd_data$ENQ , RTL___near_mem___icache___master_xactor_f_rd_data$FULL_N ; 
    wire[96:0] RTL___near_mem___icache___master_xactor_f_wr_addr$D_IN , RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_addr$CLR , RTL___near_mem___icache___master_xactor_f_wr_addr$DEQ , RTL___near_mem___icache___master_xactor_f_wr_addr$EMPTY_N , RTL___near_mem___icache___master_xactor_f_wr_addr$ENQ , RTL___near_mem___icache___master_xactor_f_wr_addr$FULL_N ; 
    wire[72:0] RTL___near_mem___icache___master_xactor_f_wr_data$D_IN , RTL___near_mem___icache___master_xactor_f_wr_data$D_OUT ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_data$CLR , RTL___near_mem___icache___master_xactor_f_wr_data$DEQ , RTL___near_mem___icache___master_xactor_f_wr_data$EMPTY_N , RTL___near_mem___icache___master_xactor_f_wr_data$ENQ , RTL___near_mem___icache___master_xactor_f_wr_data$FULL_N ; 
    wire[5:0] RTL___near_mem___icache___master_xactor_f_wr_resp$D_IN , RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_resp$CLR , RTL___near_mem___icache___master_xactor_f_wr_resp$DEQ , RTL___near_mem___icache___master_xactor_f_wr_resp$EMPTY_N , RTL___near_mem___icache___master_xactor_f_wr_resp$ENQ , RTL___near_mem___icache___master_xactor_f_wr_resp$FULL_N ; 
    wire[22:0] RTL___near_mem___icache___ram_state_and_ctag_cset$DIA , RTL___near_mem___icache___ram_state_and_ctag_cset$DIB , RTL___near_mem___icache___ram_state_and_ctag_cset$DOB ; 
    wire[6:0] RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRA , RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRB ; 
    wire RTL___near_mem___icache___ram_state_and_ctag_cset$ENA , RTL___near_mem___icache___ram_state_and_ctag_cset$ENB , RTL___near_mem___icache___ram_state_and_ctag_cset$WEA , RTL___near_mem___icache___ram_state_and_ctag_cset$WEB ; reg[63:0] RTL___near_mem___icache___ram_word64_set$DIB ; reg[8:0] RTL___near_mem___icache___ram_word64_set$ADDRB ; 
    wire[63:0] RTL___near_mem___icache___ram_word64_set$DIA , RTL___near_mem___icache___ram_word64_set$DOB ; 
    wire[8:0] RTL___near_mem___icache___ram_word64_set$ADDRA ; 
    wire RTL___near_mem___icache___ram_word64_set$ENA , RTL___near_mem___icache___ram_word64_set$ENB , RTL___near_mem___icache___ram_word64_set$WEA , RTL___near_mem___icache___ram_word64_set$WEB ; 
    wire[63:0] RTL___near_mem___icache___soc_map$m_is_IO_addr_addr , RTL___near_mem___icache___soc_map$m_is_mem_addr_addr , RTL___near_mem___icache___soc_map$m_is_near_mem_IO_addr_addr ; 
    wire RTL___near_mem___icache___soc_map$m_is_mem_addr ; 
    wire RTL___near_mem___icache___CAN_FIRE_RL_rl_ST_AMO_response , RTL___near_mem___icache___CAN_FIRE_RL_rl_cache_refill_rsps_loop , RTL___near_mem___icache___CAN_FIRE_RL_rl_discard_write_rsp , RTL___near_mem___icache___CAN_FIRE_RL_rl_drive_exception_rsp , RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req , RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_req , RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_rsp , RTL___near_mem___icache___CAN_FIRE_RL_rl_io_write_req , RTL___near_mem___icache___CAN_FIRE_RL_rl_maintain_io_read_rsp , RTL___near_mem___icache___CAN_FIRE_RL_rl_probe_and_immed_rsp , RTL___near_mem___icache___CAN_FIRE_RL_rl_rereq , RTL___near_mem___icache___CAN_FIRE_RL_rl_reset , RTL___near_mem___icache___CAN_FIRE_RL_rl_start_cache_refill , RTL___near_mem___icache___CAN_FIRE_RL_rl_start_reset , RTL___near_mem___icache___CAN_FIRE_mem_master_m_arready , RTL___near_mem___icache___CAN_FIRE_mem_master_m_awready , RTL___near_mem___icache___CAN_FIRE_mem_master_m_bvalid , RTL___near_mem___icache___CAN_FIRE_mem_master_m_rvalid , RTL___near_mem___icache___CAN_FIRE_mem_master_m_wready , RTL___near_mem___icache___CAN_FIRE_req , RTL___near_mem___icache___CAN_FIRE_server_flush_request_put , RTL___near_mem___icache___CAN_FIRE_server_flush_response_get , RTL___near_mem___icache___CAN_FIRE_server_reset_request_put , RTL___near_mem___icache___CAN_FIRE_server_reset_response_get , RTL___near_mem___icache___CAN_FIRE_set_verbosity , RTL___near_mem___icache___CAN_FIRE_tlb_flush , RTL___near_mem___icache___WILL_FIRE_RL_rl_ST_AMO_response , RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop , RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp , RTL___near_mem___icache___WILL_FIRE_RL_rl_drive_exception_rsp , RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req , RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req , RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp , RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req , RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp , RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp , RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq , RTL___near_mem___icache___WILL_FIRE_RL_rl_reset , RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill , RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset , RTL___near_mem___icache___WILL_FIRE_mem_master_m_arready , RTL___near_mem___icache___WILL_FIRE_mem_master_m_awready , RTL___near_mem___icache___WILL_FIRE_mem_master_m_bvalid , RTL___near_mem___icache___WILL_FIRE_mem_master_m_rvalid , RTL___near_mem___icache___WILL_FIRE_mem_master_m_wready , RTL___near_mem___icache___WILL_FIRE_req , RTL___near_mem___icache___WILL_FIRE_server_flush_request_put , RTL___near_mem___icache___WILL_FIRE_server_flush_response_get , RTL___near_mem___icache___WILL_FIRE_server_reset_request_put , RTL___near_mem___icache___WILL_FIRE_server_reset_response_get , RTL___near_mem___icache___WILL_FIRE_set_verbosity , RTL___near_mem___icache___WILL_FIRE_tlb_flush ; reg[63:0] RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2 ; 
    wire[98:0] RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_1 , RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
    wire[96:0] RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 , RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
    wire[22:0] RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ; 
    wire[8:0] RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_2 , RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_4 ; 
    wire[6:0] RTL___near_mem___icache___MUX_rg_cset_in_cache$write_1__VAL_1 ; 
    wire[3:0] RTL___near_mem___icache___MUX_rg_exc_code$write_1__VAL_1 , RTL___near_mem___icache___MUX_rg_state$write_1__VAL_1 , RTL___near_mem___icache___MUX_rg_state$write_1__VAL_4 , RTL___near_mem___icache___MUX_rg_state$write_1__VAL_7 , RTL___near_mem___icache___MUX_rg_state$write_1__VAL_9 ; 
    wire RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_1 , RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_2 , RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_3 , RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__SEL_1 , RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 , RTL___near_mem___icache___MUX_ram_word64_set$a_put_1__SEL_1 , RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2 , RTL___near_mem___icache___MUX_rg_error_during_refill$write_1__SEL_1 , RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_1 , RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_2 , RTL___near_mem___icache___MUX_rg_state$write_1__SEL_10 , RTL___near_mem___icache___MUX_rg_state$write_1__SEL_2 , RTL___near_mem___icache___MUX_rg_state$write_1__SEL_3 , RTL___near_mem___icache___MUX_rg_state$write_1__SEL_7 , RTL___near_mem___icache___MUX_rg_state$write_1__SEL_9 ; reg[31:0] RTL___near_mem___icache___v__h2948 ; reg[31:0] RTL___near_mem___icache___v__h3848 ; reg[31:0] RTL___near_mem___icache___v__h3949 ; reg[31:0] RTL___near_mem___icache___v__h4098 ; reg[31:0] RTL___near_mem___icache___v__h12540 ; reg[31:0] RTL___near_mem___icache___v__h14531 ; reg[31:0] RTL___near_mem___icache___v__h15336 ; reg[31:0] RTL___near_mem___icache___v__h15578 ; reg[31:0] RTL___near_mem___icache___v__h17191 ; reg[31:0] RTL___near_mem___icache___v__h17485 ; reg[31:0] RTL___near_mem___icache___v__h18585 ; reg[31:0] RTL___near_mem___icache___v__h18692 ; reg[31:0] RTL___near_mem___icache___v__h18797 ; reg[31:0] RTL___near_mem___icache___v__h18877 ; reg[31:0] RTL___near_mem___icache___v__h19505 ; reg[31:0] RTL___near_mem___icache___v__h19466 ; reg[31:0] RTL___near_mem___icache___v__h3483 ; reg[31:0] RTL___near_mem___icache___v__h19852 ; reg[31:0] RTL___near_mem___icache___v__h2942 ; reg[31:0] RTL___near_mem___icache___v__h3477 ; reg[31:0] RTL___near_mem___icache___v__h3842 ; reg[31:0] RTL___near_mem___icache___v__h3943 ; reg[31:0] RTL___near_mem___icache___v__h4092 ; reg[31:0] RTL___near_mem___icache___v__h12534 ; reg[31:0] RTL___near_mem___icache___v__h14525 ; reg[31:0] RTL___near_mem___icache___v__h15330 ; reg[31:0] RTL___near_mem___icache___v__h15572 ; reg[31:0] RTL___near_mem___icache___v__h17185 ; reg[31:0] RTL___near_mem___icache___v__h17479 ; reg[31:0] RTL___near_mem___icache___v__h18579 ; reg[31:0] RTL___near_mem___icache___v__h18686 ; reg[31:0] RTL___near_mem___icache___v__h18791 ; reg[31:0] RTL___near_mem___icache___v__h18871 ; reg[31:0] RTL___near_mem___icache___v__h19460 ; reg[31:0] RTL___near_mem___icache___v__h19499 ; reg[31:0] RTL___near_mem___icache___v__h19846 ; reg[63:0] RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 , RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 , RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 , RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 , RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 , RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 , RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 , RTL___near_mem___icache___ld_val__h17594 , RTL___near_mem___icache___mem_req_wr_data_wdata__h2699 ; reg[7:0] RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700 ; reg[2:0] RTL___near_mem___icache___value__h17372 , RTL___near_mem___icache___x__h2520 ; 
    wire[63:0] RTL___near_mem___icache____theResult___snd_fst__h2707 , RTL___near_mem___icache___cline_fabric_addr__h14584 , RTL___near_mem___icache___fabric_addr__h17243 , RTL___near_mem___icache___mem_req_wr_addr_awaddr__h2473 , RTL___near_mem___icache___result__h11657 , RTL___near_mem___icache___result__h11685 , RTL___near_mem___icache___result__h11713 , RTL___near_mem___icache___result__h11741 , RTL___near_mem___icache___result__h11769 , RTL___near_mem___icache___result__h11797 , RTL___near_mem___icache___result__h11825 , RTL___near_mem___icache___result__h11870 , RTL___near_mem___icache___result__h11898 , RTL___near_mem___icache___result__h11926 , RTL___near_mem___icache___result__h11954 , RTL___near_mem___icache___result__h11982 , RTL___near_mem___icache___result__h12010 , RTL___near_mem___icache___result__h12038 , RTL___near_mem___icache___result__h12066 , RTL___near_mem___icache___result__h12111 , RTL___near_mem___icache___result__h12139 , RTL___near_mem___icache___result__h12167 , RTL___near_mem___icache___result__h12195 , RTL___near_mem___icache___result__h12236 , RTL___near_mem___icache___result__h12264 , RTL___near_mem___icache___result__h12292 , RTL___near_mem___icache___result__h12320 , RTL___near_mem___icache___result__h12361 , RTL___near_mem___icache___result__h12389 , RTL___near_mem___icache___result__h12428 , RTL___near_mem___icache___result__h12456 , RTL___near_mem___icache___result__h17654 , RTL___near_mem___icache___result__h17684 , RTL___near_mem___icache___result__h17711 , RTL___near_mem___icache___result__h17738 , RTL___near_mem___icache___result__h17765 , RTL___near_mem___icache___result__h17792 , RTL___near_mem___icache___result__h17819 , RTL___near_mem___icache___result__h17846 , RTL___near_mem___icache___result__h17890 , RTL___near_mem___icache___result__h17917 , RTL___near_mem___icache___result__h17944 , RTL___near_mem___icache___result__h17971 , RTL___near_mem___icache___result__h17998 , RTL___near_mem___icache___result__h18025 , RTL___near_mem___icache___result__h18052 , RTL___near_mem___icache___result__h18079 , RTL___near_mem___icache___result__h18123 , RTL___near_mem___icache___result__h18150 , RTL___near_mem___icache___result__h18177 , RTL___near_mem___icache___result__h18204 , RTL___near_mem___icache___result__h18244 , RTL___near_mem___icache___result__h18271 , RTL___near_mem___icache___result__h18298 , RTL___near_mem___icache___result__h18325 , RTL___near_mem___icache___result__h18365 , RTL___near_mem___icache___result__h18392 , RTL___near_mem___icache___result__h18430 , RTL___near_mem___icache___result__h18457 , RTL___near_mem___icache___result__h5301 , RTL___near_mem___icache___word64__h5094 , RTL___near_mem___icache___y__h5337 ; 
    wire[31:0] RTL___near_mem___icache___cline_addr__h14583 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 , RTL___near_mem___icache___word64094_BITS_31_TO_0__q17 , RTL___near_mem___icache___word64094_BITS_63_TO_32__q24 ; 
    wire[21:0] RTL___near_mem___icache___pa_ctag__h4952 ; 
    wire[15:0] RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 , RTL___near_mem___icache___word64094_BITS_15_TO_0__q16 , RTL___near_mem___icache___word64094_BITS_31_TO_16__q20 , RTL___near_mem___icache___word64094_BITS_47_TO_32__q23 , RTL___near_mem___icache___word64094_BITS_63_TO_48__q27 ; 
    wire[7:0] RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 , RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 , RTL___near_mem___icache___strobe64__h2637 , RTL___near_mem___icache___strobe64__h2639 , RTL___near_mem___icache___strobe64__h2641 , RTL___near_mem___icache___word64094_BITS_15_TO_8__q18 , RTL___near_mem___icache___word64094_BITS_23_TO_16__q19 , RTL___near_mem___icache___word64094_BITS_31_TO_24__q21 , RTL___near_mem___icache___word64094_BITS_39_TO_32__q22 , RTL___near_mem___icache___word64094_BITS_47_TO_40__q25 , RTL___near_mem___icache___word64094_BITS_55_TO_48__q26 , RTL___near_mem___icache___word64094_BITS_63_TO_56__q28 , RTL___near_mem___icache___word64094_BITS_7_TO_0__q15 ; 
    wire[5:0] RTL___near_mem___icache___shift_bits__h2487 ; 
    wire[3:0] RTL___near_mem___icache___access_exc_code__h2256 , RTL___near_mem___icache___b__h14485 ; 
    wire RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 , RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 , RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 , RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 , RTL___near_mem___icache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 , RTL___near_mem___icache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 , RTL___near_mem___icache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 , RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 , RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 , RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 ; 
  assign  RTL___near_mem___icache___RDY_set_verbosity =1'd1; 
  assign  RTL___near_mem___icache___CAN_FIRE_set_verbosity =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_set_verbosity = RTL___near_mem___icache___EN_set_verbosity ; 
  assign  RTL___near_mem___icache___RDY_server_reset_request_put = RTL___near_mem___icache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___icache___CAN_FIRE_server_reset_request_put = RTL___near_mem___icache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_server_reset_request_put = RTL___near_mem___icache___EN_server_reset_request_put ; 
  assign  RTL___near_mem___icache___RDY_server_reset_response_get =! RTL___near_mem___icache___f_reset_rsps$D_OUT && RTL___near_mem___icache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___icache___CAN_FIRE_server_reset_response_get =! RTL___near_mem___icache___f_reset_rsps$D_OUT && RTL___near_mem___icache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_server_reset_response_get = RTL___near_mem___icache___EN_server_reset_response_get ; 
  assign  RTL___near_mem___icache___CAN_FIRE_req =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_req = RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___valid = RTL___near_mem___icache___dw_valid$whas ; 
  assign  RTL___near_mem___icache___addr = RTL___near_mem___icache___rg_addr ; 
  always @(       RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_1                    or   RTL___near_mem___icache___ld_val__h17594              or   RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_2             or   RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2            or   RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_3           or   RTL___near_mem___icache___rg_ld_val  )
         begin 
             case (1'b1) 
              RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_1  : 
                  RTL___near_mem___icache___word64  = RTL___near_mem___icache___ld_val__h17594 ; 
              RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_2  : 
                  RTL___near_mem___icache___word64  = RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2 ; 
              RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_3  : 
                  RTL___near_mem___icache___word64  = RTL___near_mem___icache___rg_ld_val ;
              default : 
                  RTL___near_mem___icache___word64  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL___near_mem___icache___st_amo_val = RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_2  ? 64'd0: RTL___near_mem___icache___rg_st_amo_val ; 
  assign  RTL___near_mem___icache___exc = RTL___near_mem___icache___rg_state ==4'd4; 
  assign  RTL___near_mem___icache___exc_code = RTL___near_mem___icache___rg_exc_code ; 
  assign  RTL___near_mem___icache___RDY_server_flush_request_put = RTL___near_mem___icache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___icache___CAN_FIRE_server_flush_request_put = RTL___near_mem___icache___f_reset_reqs$FULL_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_server_flush_request_put = RTL___near_mem___icache___EN_server_flush_request_put ; 
  assign  RTL___near_mem___icache___RDY_server_flush_response_get = RTL___near_mem___icache___f_reset_rsps$D_OUT && RTL___near_mem___icache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___icache___CAN_FIRE_server_flush_response_get = RTL___near_mem___icache___f_reset_rsps$D_OUT && RTL___near_mem___icache___f_reset_rsps$EMPTY_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_server_flush_response_get = RTL___near_mem___icache___EN_server_flush_response_get ; 
  assign  RTL___near_mem___icache___RDY_tlb_flush =1'd1; 
  assign  RTL___near_mem___icache___CAN_FIRE_tlb_flush =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_tlb_flush = RTL___near_mem___icache___EN_tlb_flush ; 
  assign  RTL___near_mem___icache___mem_master_awvalid = RTL___near_mem___icache___master_xactor_f_wr_addr$EMPTY_N ; 
  assign  RTL___near_mem___icache___mem_master_awid = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [96:93]; 
  assign  RTL___near_mem___icache___mem_master_awaddr = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [92:29]; 
  assign  RTL___near_mem___icache___mem_master_awlen = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [28:21]; 
  assign  RTL___near_mem___icache___mem_master_awsize = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [20:18]; 
  assign  RTL___near_mem___icache___mem_master_awburst = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [17:16]; 
  assign  RTL___near_mem___icache___mem_master_awlock = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [15]; 
  assign  RTL___near_mem___icache___mem_master_awcache = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [14:11]; 
  assign  RTL___near_mem___icache___mem_master_awprot = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [10:8]; 
  assign  RTL___near_mem___icache___mem_master_awqos = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [7:4]; 
  assign  RTL___near_mem___icache___mem_master_awregion = RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT [3:0]; 
  assign  RTL___near_mem___icache___CAN_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_mem_master_m_awready =1'd1; 
  assign  RTL___near_mem___icache___mem_master_wvalid = RTL___near_mem___icache___master_xactor_f_wr_data$EMPTY_N ; 
  assign  RTL___near_mem___icache___mem_master_wdata = RTL___near_mem___icache___master_xactor_f_wr_data$D_OUT [72:9]; 
  assign  RTL___near_mem___icache___mem_master_wstrb = RTL___near_mem___icache___master_xactor_f_wr_data$D_OUT [8:1]; 
  assign  RTL___near_mem___icache___mem_master_wlast = RTL___near_mem___icache___master_xactor_f_wr_data$D_OUT [0]; 
  assign  RTL___near_mem___icache___CAN_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_mem_master_m_wready =1'd1; 
  assign  RTL___near_mem___icache___CAN_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_mem_master_m_bvalid =1'd1; 
  assign  RTL___near_mem___icache___mem_master_bready = RTL___near_mem___icache___master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL___near_mem___icache___mem_master_arvalid = RTL___near_mem___icache___master_xactor_f_rd_addr$EMPTY_N ; 
  assign  RTL___near_mem___icache___mem_master_arid = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [96:93]; 
  assign  RTL___near_mem___icache___mem_master_araddr = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [92:29]; 
  assign  RTL___near_mem___icache___mem_master_arlen = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [28:21]; 
  assign  RTL___near_mem___icache___mem_master_arsize = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [20:18]; 
  assign  RTL___near_mem___icache___mem_master_arburst = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [17:16]; 
  assign  RTL___near_mem___icache___mem_master_arlock = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [15]; 
  assign  RTL___near_mem___icache___mem_master_arcache = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [14:11]; 
  assign  RTL___near_mem___icache___mem_master_arprot = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [10:8]; 
  assign  RTL___near_mem___icache___mem_master_arqos = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [7:4]; 
  assign  RTL___near_mem___icache___mem_master_arregion = RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT [3:0]; 
  assign  RTL___near_mem___icache___CAN_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_mem_master_m_arready =1'd1; 
  assign  RTL___near_mem___icache___CAN_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_mem_master_m_rvalid =1'd1; 
  assign  RTL___near_mem___icache___mem_master_rready = RTL___near_mem___icache___master_xactor_f_rd_data$FULL_N ;  
    
    reg RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
    reg RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; reg[ RTL___near_mem___icache___f_fabric_write_reqs___width -1:0] RTL___near_mem___icache___f_fabric_write_reqs___data0_reg ; reg[ RTL___near_mem___icache___f_fabric_write_reqs___width -1:0] RTL___near_mem___icache___f_fabric_write_reqs___data1_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___FULL_N = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___EMPTY_N = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___D_OUT = RTL___near_mem___icache___f_fabric_write_reqs___data0_reg ; 
    wire RTL___near_mem___icache___f_fabric_write_reqs___d0di =( RTL___near_mem___icache___f_fabric_write_reqs___ENQ &&! RTL___near_mem___icache___f_fabric_write_reqs___empty_reg )||( RTL___near_mem___icache___f_fabric_write_reqs___ENQ && RTL___near_mem___icache___f_fabric_write_reqs___DEQ && RTL___near_mem___icache___f_fabric_write_reqs___full_reg ); 
    wire RTL___near_mem___icache___f_fabric_write_reqs___d0d1 = RTL___near_mem___icache___f_fabric_write_reqs___DEQ &&! RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
    wire RTL___near_mem___icache___f_fabric_write_reqs___d0h =((! RTL___near_mem___icache___f_fabric_write_reqs___DEQ )&&(! RTL___near_mem___icache___f_fabric_write_reqs___ENQ ))||(! RTL___near_mem___icache___f_fabric_write_reqs___DEQ && RTL___near_mem___icache___f_fabric_write_reqs___empty_reg )||(! RTL___near_mem___icache___f_fabric_write_reqs___ENQ && RTL___near_mem___icache___f_fabric_write_reqs___full_reg ); 
    wire RTL___near_mem___icache___f_fabric_write_reqs___d1di = RTL___near_mem___icache___f_fabric_write_reqs___ENQ & RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___f_fabric_write_reqs___CLK )
         begin 
             if ( RTL___near_mem___icache___f_fabric_write_reqs___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___f_fabric_write_reqs___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___f_fabric_write_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___f_fabric_write_reqs___CLR )
                         begin  
                             RTL___near_mem___icache___f_fabric_write_reqs___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___f_fabric_write_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___f_fabric_write_reqs___ENQ &&! RTL___near_mem___icache___f_fabric_write_reqs___DEQ )
                             begin  
                                 RTL___near_mem___icache___f_fabric_write_reqs___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___f_fabric_write_reqs___full_reg  <=! RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___f_fabric_write_reqs___DEQ &&! RTL___near_mem___icache___f_fabric_write_reqs___ENQ )
                                 begin  
                                     RTL___near_mem___icache___f_fabric_write_reqs___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___f_fabric_write_reqs___empty_reg  <=! RTL___near_mem___icache___f_fabric_write_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___f_fabric_write_reqs___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___f_fabric_write_reqs___data0_reg  <={ RTL___near_mem___icache___f_fabric_write_reqs___width { RTL___near_mem___icache___f_fabric_write_reqs___d0di }}& RTL___near_mem___icache___f_fabric_write_reqs___D_IN |{ RTL___near_mem___icache___f_fabric_write_reqs___width { RTL___near_mem___icache___f_fabric_write_reqs___d0d1 }}& RTL___near_mem___icache___f_fabric_write_reqs___data1_reg |{ RTL___near_mem___icache___f_fabric_write_reqs___width { RTL___near_mem___icache___f_fabric_write_reqs___d0h }}& RTL___near_mem___icache___f_fabric_write_reqs___data0_reg ; 
                 RTL___near_mem___icache___f_fabric_write_reqs___data1_reg  <= RTL___near_mem___icache___f_fabric_write_reqs___d1di  ?  RTL___near_mem___icache___f_fabric_write_reqs___D_IN : RTL___near_mem___icache___f_fabric_write_reqs___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___f_fabric_write_reqs___CLK )
         begin : RTL___near_mem___icache___f_fabric_write_reqs___error_checks 
           reg RTL___near_mem___icache___f_fabric_write_reqs___deqerror , RTL___near_mem___icache___f_fabric_write_reqs___enqerror ; 
             RTL___near_mem___icache___f_fabric_write_reqs___deqerror  =0; 
             RTL___near_mem___icache___f_fabric_write_reqs___enqerror  =0;
             if ( RTL___near_mem___icache___f_fabric_write_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___f_fabric_write_reqs___empty_reg && RTL___near_mem___icache___f_fabric_write_reqs___DEQ )
                         begin  
                             RTL___near_mem___icache___f_fabric_write_reqs___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___f_fabric_write_reqs___full_reg && RTL___near_mem___icache___f_fabric_write_reqs___ENQ &&(! RTL___near_mem___icache___f_fabric_write_reqs___DEQ || RTL___near_mem___icache___f_fabric_write_reqs___guarded ))
                         begin  
                             RTL___near_mem___icache___f_fabric_write_reqs___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___empty_reg ;
    reg RTL___near_mem___icache___f_reset_reqs___full_reg ; 
    reg RTL___near_mem___icache___f_reset_reqs___empty_reg ; reg[ RTL___near_mem___icache___f_reset_reqs___width -1:0] RTL___near_mem___icache___f_reset_reqs___data0_reg ; reg[ RTL___near_mem___icache___f_reset_reqs___width -1:0] RTL___near_mem___icache___f_reset_reqs___data1_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___FULL_N = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___EMPTY_N = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___D_OUT = RTL___near_mem___icache___f_reset_reqs___data0_reg ; 
    wire RTL___near_mem___icache___f_reset_reqs___d0di =( RTL___near_mem___icache___f_reset_reqs___ENQ &&! RTL___near_mem___icache___f_reset_reqs___empty_reg )||( RTL___near_mem___icache___f_reset_reqs___ENQ && RTL___near_mem___icache___f_reset_reqs___DEQ && RTL___near_mem___icache___f_reset_reqs___full_reg ); 
    wire RTL___near_mem___icache___f_reset_reqs___d0d1 = RTL___near_mem___icache___f_reset_reqs___DEQ &&! RTL___near_mem___icache___f_reset_reqs___full_reg ; 
    wire RTL___near_mem___icache___f_reset_reqs___d0h =((! RTL___near_mem___icache___f_reset_reqs___DEQ )&&(! RTL___near_mem___icache___f_reset_reqs___ENQ ))||(! RTL___near_mem___icache___f_reset_reqs___DEQ && RTL___near_mem___icache___f_reset_reqs___empty_reg )||(! RTL___near_mem___icache___f_reset_reqs___ENQ && RTL___near_mem___icache___f_reset_reqs___full_reg ); 
    wire RTL___near_mem___icache___f_reset_reqs___d1di = RTL___near_mem___icache___f_reset_reqs___ENQ & RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___f_reset_reqs___CLK )
         begin 
             if ( RTL___near_mem___icache___f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___f_reset_reqs___CLR )
                         begin  
                             RTL___near_mem___icache___f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___f_reset_reqs___ENQ &&! RTL___near_mem___icache___f_reset_reqs___DEQ )
                             begin  
                                 RTL___near_mem___icache___f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___f_reset_reqs___full_reg  <=! RTL___near_mem___icache___f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___f_reset_reqs___DEQ &&! RTL___near_mem___icache___f_reset_reqs___ENQ )
                                 begin  
                                     RTL___near_mem___icache___f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___f_reset_reqs___empty_reg  <=! RTL___near_mem___icache___f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___f_reset_reqs___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___f_reset_reqs___data0_reg  <={ RTL___near_mem___icache___f_reset_reqs___width { RTL___near_mem___icache___f_reset_reqs___d0di }}& RTL___near_mem___icache___f_reset_reqs___D_IN |{ RTL___near_mem___icache___f_reset_reqs___width { RTL___near_mem___icache___f_reset_reqs___d0d1 }}& RTL___near_mem___icache___f_reset_reqs___data1_reg |{ RTL___near_mem___icache___f_reset_reqs___width { RTL___near_mem___icache___f_reset_reqs___d0h }}& RTL___near_mem___icache___f_reset_reqs___data0_reg ; 
                 RTL___near_mem___icache___f_reset_reqs___data1_reg  <= RTL___near_mem___icache___f_reset_reqs___d1di  ?  RTL___near_mem___icache___f_reset_reqs___D_IN : RTL___near_mem___icache___f_reset_reqs___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___f_reset_reqs___CLK )
         begin : RTL___near_mem___icache___f_reset_reqs___error_checks 
           reg RTL___near_mem___icache___f_reset_reqs___deqerror , RTL___near_mem___icache___f_reset_reqs___enqerror ; 
             RTL___near_mem___icache___f_reset_reqs___deqerror  =0; 
             RTL___near_mem___icache___f_reset_reqs___enqerror  =0;
             if ( RTL___near_mem___icache___f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___f_reset_reqs___empty_reg && RTL___near_mem___icache___f_reset_reqs___DEQ )
                         begin  
                             RTL___near_mem___icache___f_reset_reqs___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___f_reset_reqs___full_reg && RTL___near_mem___icache___f_reset_reqs___ENQ &&(! RTL___near_mem___icache___f_reset_reqs___DEQ || RTL___near_mem___icache___f_reset_reqs___guarded ))
                         begin  
                             RTL___near_mem___icache___f_reset_reqs___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___empty_reg ;
    reg RTL___near_mem___icache___f_reset_rsps___full_reg ; 
    reg RTL___near_mem___icache___f_reset_rsps___empty_reg ; reg[ RTL___near_mem___icache___f_reset_rsps___width -1:0] RTL___near_mem___icache___f_reset_rsps___data0_reg ; reg[ RTL___near_mem___icache___f_reset_rsps___width -1:0] RTL___near_mem___icache___f_reset_rsps___data1_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___FULL_N = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___EMPTY_N = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___D_OUT = RTL___near_mem___icache___f_reset_rsps___data0_reg ; 
    wire RTL___near_mem___icache___f_reset_rsps___d0di =( RTL___near_mem___icache___f_reset_rsps___ENQ &&! RTL___near_mem___icache___f_reset_rsps___empty_reg )||( RTL___near_mem___icache___f_reset_rsps___ENQ && RTL___near_mem___icache___f_reset_rsps___DEQ && RTL___near_mem___icache___f_reset_rsps___full_reg ); 
    wire RTL___near_mem___icache___f_reset_rsps___d0d1 = RTL___near_mem___icache___f_reset_rsps___DEQ &&! RTL___near_mem___icache___f_reset_rsps___full_reg ; 
    wire RTL___near_mem___icache___f_reset_rsps___d0h =((! RTL___near_mem___icache___f_reset_rsps___DEQ )&&(! RTL___near_mem___icache___f_reset_rsps___ENQ ))||(! RTL___near_mem___icache___f_reset_rsps___DEQ && RTL___near_mem___icache___f_reset_rsps___empty_reg )||(! RTL___near_mem___icache___f_reset_rsps___ENQ && RTL___near_mem___icache___f_reset_rsps___full_reg ); 
    wire RTL___near_mem___icache___f_reset_rsps___d1di = RTL___near_mem___icache___f_reset_rsps___ENQ & RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___f_reset_rsps___CLK )
         begin 
             if ( RTL___near_mem___icache___f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___f_reset_rsps___CLR )
                         begin  
                             RTL___near_mem___icache___f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___f_reset_rsps___ENQ &&! RTL___near_mem___icache___f_reset_rsps___DEQ )
                             begin  
                                 RTL___near_mem___icache___f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___f_reset_rsps___full_reg  <=! RTL___near_mem___icache___f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___f_reset_rsps___DEQ &&! RTL___near_mem___icache___f_reset_rsps___ENQ )
                                 begin  
                                     RTL___near_mem___icache___f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___f_reset_rsps___empty_reg  <=! RTL___near_mem___icache___f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___f_reset_rsps___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___f_reset_rsps___data0_reg  <={ RTL___near_mem___icache___f_reset_rsps___width { RTL___near_mem___icache___f_reset_rsps___d0di }}& RTL___near_mem___icache___f_reset_rsps___D_IN |{ RTL___near_mem___icache___f_reset_rsps___width { RTL___near_mem___icache___f_reset_rsps___d0d1 }}& RTL___near_mem___icache___f_reset_rsps___data1_reg |{ RTL___near_mem___icache___f_reset_rsps___width { RTL___near_mem___icache___f_reset_rsps___d0h }}& RTL___near_mem___icache___f_reset_rsps___data0_reg ; 
                 RTL___near_mem___icache___f_reset_rsps___data1_reg  <= RTL___near_mem___icache___f_reset_rsps___d1di  ?  RTL___near_mem___icache___f_reset_rsps___D_IN : RTL___near_mem___icache___f_reset_rsps___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___f_reset_rsps___CLK )
         begin : RTL___near_mem___icache___f_reset_rsps___error_checks 
           reg RTL___near_mem___icache___f_reset_rsps___deqerror , RTL___near_mem___icache___f_reset_rsps___enqerror ; 
             RTL___near_mem___icache___f_reset_rsps___deqerror  =0; 
             RTL___near_mem___icache___f_reset_rsps___enqerror  =0;
             if ( RTL___near_mem___icache___f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___f_reset_rsps___empty_reg && RTL___near_mem___icache___f_reset_rsps___DEQ )
                         begin  
                             RTL___near_mem___icache___f_reset_rsps___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___f_reset_rsps___full_reg && RTL___near_mem___icache___f_reset_rsps___ENQ &&(! RTL___near_mem___icache___f_reset_rsps___DEQ || RTL___near_mem___icache___f_reset_rsps___guarded ))
                         begin  
                             RTL___near_mem___icache___f_reset_rsps___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___full_reg ; 
  assign  RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___empty_reg ;
    reg RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
    reg RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; reg[ RTL___near_mem___icache___master_xactor_f_rd_addr___width -1:0] RTL___near_mem___icache___master_xactor_f_rd_addr___data0_reg ; reg[ RTL___near_mem___icache___master_xactor_f_rd_addr___width -1:0] RTL___near_mem___icache___master_xactor_f_rd_addr___data1_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___FULL_N = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___EMPTY_N = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___D_OUT = RTL___near_mem___icache___master_xactor_f_rd_addr___data0_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___d0di =( RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ &&! RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg )||( RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ && RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ && RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___d0d1 = RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ &&! RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___d0h =((! RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ )&&(! RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ ))||(! RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ && RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg )||(! RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ && RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_rd_addr___d1di = RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ & RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_addr___CLK )
         begin 
             if ( RTL___near_mem___icache___master_xactor_f_rd_addr___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___master_xactor_f_rd_addr___CLR )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ &&! RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ )
                             begin  
                                 RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg  <=! RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ &&! RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ )
                                 begin  
                                     RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg  <=! RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_addr___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___master_xactor_f_rd_addr___data0_reg  <={ RTL___near_mem___icache___master_xactor_f_rd_addr___width { RTL___near_mem___icache___master_xactor_f_rd_addr___d0di }}& RTL___near_mem___icache___master_xactor_f_rd_addr___D_IN |{ RTL___near_mem___icache___master_xactor_f_rd_addr___width { RTL___near_mem___icache___master_xactor_f_rd_addr___d0d1 }}& RTL___near_mem___icache___master_xactor_f_rd_addr___data1_reg |{ RTL___near_mem___icache___master_xactor_f_rd_addr___width { RTL___near_mem___icache___master_xactor_f_rd_addr___d0h }}& RTL___near_mem___icache___master_xactor_f_rd_addr___data0_reg ; 
                 RTL___near_mem___icache___master_xactor_f_rd_addr___data1_reg  <= RTL___near_mem___icache___master_xactor_f_rd_addr___d1di  ?  RTL___near_mem___icache___master_xactor_f_rd_addr___D_IN : RTL___near_mem___icache___master_xactor_f_rd_addr___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_addr___CLK )
         begin : RTL___near_mem___icache___master_xactor_f_rd_addr___error_checks 
           reg RTL___near_mem___icache___master_xactor_f_rd_addr___deqerror , RTL___near_mem___icache___master_xactor_f_rd_addr___enqerror ; 
             RTL___near_mem___icache___master_xactor_f_rd_addr___deqerror  =0; 
             RTL___near_mem___icache___master_xactor_f_rd_addr___enqerror  =0;
             if ( RTL___near_mem___icache___master_xactor_f_rd_addr___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg && RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_addr___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg && RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ &&(! RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ || RTL___near_mem___icache___master_xactor_f_rd_addr___guarded ))
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_addr___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___empty_reg ;
    reg RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
    reg RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; reg[ RTL___near_mem___icache___master_xactor_f_rd_data___width -1:0] RTL___near_mem___icache___master_xactor_f_rd_data___data0_reg ; reg[ RTL___near_mem___icache___master_xactor_f_rd_data___width -1:0] RTL___near_mem___icache___master_xactor_f_rd_data___data1_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___FULL_N = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___EMPTY_N = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___D_OUT = RTL___near_mem___icache___master_xactor_f_rd_data___data0_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_data___d0di =( RTL___near_mem___icache___master_xactor_f_rd_data___ENQ &&! RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg )||( RTL___near_mem___icache___master_xactor_f_rd_data___ENQ && RTL___near_mem___icache___master_xactor_f_rd_data___DEQ && RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_rd_data___d0d1 = RTL___near_mem___icache___master_xactor_f_rd_data___DEQ &&! RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_rd_data___d0h =((! RTL___near_mem___icache___master_xactor_f_rd_data___DEQ )&&(! RTL___near_mem___icache___master_xactor_f_rd_data___ENQ ))||(! RTL___near_mem___icache___master_xactor_f_rd_data___DEQ && RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg )||(! RTL___near_mem___icache___master_xactor_f_rd_data___ENQ && RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_rd_data___d1di = RTL___near_mem___icache___master_xactor_f_rd_data___ENQ & RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_data___CLK )
         begin 
             if ( RTL___near_mem___icache___master_xactor_f_rd_data___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___master_xactor_f_rd_data___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___master_xactor_f_rd_data___CLR )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___master_xactor_f_rd_data___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___master_xactor_f_rd_data___ENQ &&! RTL___near_mem___icache___master_xactor_f_rd_data___DEQ )
                             begin  
                                 RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___master_xactor_f_rd_data___full_reg  <=! RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___master_xactor_f_rd_data___DEQ &&! RTL___near_mem___icache___master_xactor_f_rd_data___ENQ )
                                 begin  
                                     RTL___near_mem___icache___master_xactor_f_rd_data___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg  <=! RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_data___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___master_xactor_f_rd_data___data0_reg  <={ RTL___near_mem___icache___master_xactor_f_rd_data___width { RTL___near_mem___icache___master_xactor_f_rd_data___d0di }}& RTL___near_mem___icache___master_xactor_f_rd_data___D_IN |{ RTL___near_mem___icache___master_xactor_f_rd_data___width { RTL___near_mem___icache___master_xactor_f_rd_data___d0d1 }}& RTL___near_mem___icache___master_xactor_f_rd_data___data1_reg |{ RTL___near_mem___icache___master_xactor_f_rd_data___width { RTL___near_mem___icache___master_xactor_f_rd_data___d0h }}& RTL___near_mem___icache___master_xactor_f_rd_data___data0_reg ; 
                 RTL___near_mem___icache___master_xactor_f_rd_data___data1_reg  <= RTL___near_mem___icache___master_xactor_f_rd_data___d1di  ?  RTL___near_mem___icache___master_xactor_f_rd_data___D_IN : RTL___near_mem___icache___master_xactor_f_rd_data___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_rd_data___CLK )
         begin : RTL___near_mem___icache___master_xactor_f_rd_data___error_checks 
           reg RTL___near_mem___icache___master_xactor_f_rd_data___deqerror , RTL___near_mem___icache___master_xactor_f_rd_data___enqerror ; 
             RTL___near_mem___icache___master_xactor_f_rd_data___deqerror  =0; 
             RTL___near_mem___icache___master_xactor_f_rd_data___enqerror  =0;
             if ( RTL___near_mem___icache___master_xactor_f_rd_data___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg && RTL___near_mem___icache___master_xactor_f_rd_data___DEQ )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_data___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___master_xactor_f_rd_data___full_reg && RTL___near_mem___icache___master_xactor_f_rd_data___ENQ &&(! RTL___near_mem___icache___master_xactor_f_rd_data___DEQ || RTL___near_mem___icache___master_xactor_f_rd_data___guarded ))
                         begin  
                             RTL___near_mem___icache___master_xactor_f_rd_data___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___empty_reg ;
    reg RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
    reg RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_addr___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_addr___data0_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_addr___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_addr___data1_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___FULL_N = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___D_OUT = RTL___near_mem___icache___master_xactor_f_wr_addr___data0_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___d0di =( RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg )||( RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ && RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ && RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___d0d1 = RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___d0h =((! RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ )&&(! RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ ))||(! RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ && RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg )||(! RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ && RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_addr___d1di = RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ & RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_addr___CLK )
         begin 
             if ( RTL___near_mem___icache___master_xactor_f_wr_addr___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___master_xactor_f_wr_addr___CLR )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ )
                             begin  
                                 RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ )
                                 begin  
                                     RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_addr___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___master_xactor_f_wr_addr___data0_reg  <={ RTL___near_mem___icache___master_xactor_f_wr_addr___width { RTL___near_mem___icache___master_xactor_f_wr_addr___d0di }}& RTL___near_mem___icache___master_xactor_f_wr_addr___D_IN |{ RTL___near_mem___icache___master_xactor_f_wr_addr___width { RTL___near_mem___icache___master_xactor_f_wr_addr___d0d1 }}& RTL___near_mem___icache___master_xactor_f_wr_addr___data1_reg |{ RTL___near_mem___icache___master_xactor_f_wr_addr___width { RTL___near_mem___icache___master_xactor_f_wr_addr___d0h }}& RTL___near_mem___icache___master_xactor_f_wr_addr___data0_reg ; 
                 RTL___near_mem___icache___master_xactor_f_wr_addr___data1_reg  <= RTL___near_mem___icache___master_xactor_f_wr_addr___d1di  ?  RTL___near_mem___icache___master_xactor_f_wr_addr___D_IN : RTL___near_mem___icache___master_xactor_f_wr_addr___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_addr___CLK )
         begin : RTL___near_mem___icache___master_xactor_f_wr_addr___error_checks 
           reg RTL___near_mem___icache___master_xactor_f_wr_addr___deqerror , RTL___near_mem___icache___master_xactor_f_wr_addr___enqerror ; 
             RTL___near_mem___icache___master_xactor_f_wr_addr___deqerror  =0; 
             RTL___near_mem___icache___master_xactor_f_wr_addr___enqerror  =0;
             if ( RTL___near_mem___icache___master_xactor_f_wr_addr___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg && RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_addr___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg && RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ &&(! RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ || RTL___near_mem___icache___master_xactor_f_wr_addr___guarded ))
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_addr___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___empty_reg ;
    reg RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
    reg RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_data___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_data___data0_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_data___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_data___data1_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___FULL_N = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___D_OUT = RTL___near_mem___icache___master_xactor_f_wr_data___data0_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_data___d0di =( RTL___near_mem___icache___master_xactor_f_wr_data___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg )||( RTL___near_mem___icache___master_xactor_f_wr_data___ENQ && RTL___near_mem___icache___master_xactor_f_wr_data___DEQ && RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_data___d0d1 = RTL___near_mem___icache___master_xactor_f_wr_data___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_data___d0h =((! RTL___near_mem___icache___master_xactor_f_wr_data___DEQ )&&(! RTL___near_mem___icache___master_xactor_f_wr_data___ENQ ))||(! RTL___near_mem___icache___master_xactor_f_wr_data___DEQ && RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg )||(! RTL___near_mem___icache___master_xactor_f_wr_data___ENQ && RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_data___d1di = RTL___near_mem___icache___master_xactor_f_wr_data___ENQ & RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_data___CLK )
         begin 
             if ( RTL___near_mem___icache___master_xactor_f_wr_data___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___master_xactor_f_wr_data___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___master_xactor_f_wr_data___CLR )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___master_xactor_f_wr_data___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___master_xactor_f_wr_data___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_data___DEQ )
                             begin  
                                 RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___master_xactor_f_wr_data___full_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___master_xactor_f_wr_data___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_data___ENQ )
                                 begin  
                                     RTL___near_mem___icache___master_xactor_f_wr_data___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_data___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___master_xactor_f_wr_data___data0_reg  <={ RTL___near_mem___icache___master_xactor_f_wr_data___width { RTL___near_mem___icache___master_xactor_f_wr_data___d0di }}& RTL___near_mem___icache___master_xactor_f_wr_data___D_IN |{ RTL___near_mem___icache___master_xactor_f_wr_data___width { RTL___near_mem___icache___master_xactor_f_wr_data___d0d1 }}& RTL___near_mem___icache___master_xactor_f_wr_data___data1_reg |{ RTL___near_mem___icache___master_xactor_f_wr_data___width { RTL___near_mem___icache___master_xactor_f_wr_data___d0h }}& RTL___near_mem___icache___master_xactor_f_wr_data___data0_reg ; 
                 RTL___near_mem___icache___master_xactor_f_wr_data___data1_reg  <= RTL___near_mem___icache___master_xactor_f_wr_data___d1di  ?  RTL___near_mem___icache___master_xactor_f_wr_data___D_IN : RTL___near_mem___icache___master_xactor_f_wr_data___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_data___CLK )
         begin : RTL___near_mem___icache___master_xactor_f_wr_data___error_checks 
           reg RTL___near_mem___icache___master_xactor_f_wr_data___deqerror , RTL___near_mem___icache___master_xactor_f_wr_data___enqerror ; 
             RTL___near_mem___icache___master_xactor_f_wr_data___deqerror  =0; 
             RTL___near_mem___icache___master_xactor_f_wr_data___enqerror  =0;
             if ( RTL___near_mem___icache___master_xactor_f_wr_data___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg && RTL___near_mem___icache___master_xactor_f_wr_data___DEQ )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_data___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_data___full_reg && RTL___near_mem___icache___master_xactor_f_wr_data___ENQ &&(! RTL___near_mem___icache___master_xactor_f_wr_data___DEQ || RTL___near_mem___icache___master_xactor_f_wr_data___guarded ))
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_data___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___empty_reg ;
    reg RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
    reg RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_resp___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_resp___data0_reg ; reg[ RTL___near_mem___icache___master_xactor_f_wr_resp___width -1:0] RTL___near_mem___icache___master_xactor_f_wr_resp___data1_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___FULL_N = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___D_OUT = RTL___near_mem___icache___master_xactor_f_wr_resp___data0_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___d0di =( RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg )||( RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ && RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ && RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___d0d1 = RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___d0h =((! RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ )&&(! RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ ))||(! RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ && RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg )||(! RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ && RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ); 
    wire RTL___near_mem___icache___master_xactor_f_wr_resp___d1di = RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ & RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_resp___CLK )
         begin 
             if ( RTL___near_mem___icache___master_xactor_f_wr_resp___RST ==1'b0)
                 begin  
                     RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg  <=1'b0; 
                     RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___master_xactor_f_wr_resp___CLR )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg  <=1'b0; 
                             RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ &&! RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ )
                             begin  
                                 RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg  <=1'b1; 
                                 RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ;
                             end 
                          else 
                             if ( RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ &&! RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ )
                                 begin  
                                     RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg  <=1'b1; 
                                     RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg  <=! RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_resp___CLK )
         begin 
             begin  
                 RTL___near_mem___icache___master_xactor_f_wr_resp___data0_reg  <={ RTL___near_mem___icache___master_xactor_f_wr_resp___width { RTL___near_mem___icache___master_xactor_f_wr_resp___d0di }}& RTL___near_mem___icache___master_xactor_f_wr_resp___D_IN |{ RTL___near_mem___icache___master_xactor_f_wr_resp___width { RTL___near_mem___icache___master_xactor_f_wr_resp___d0d1 }}& RTL___near_mem___icache___master_xactor_f_wr_resp___data1_reg |{ RTL___near_mem___icache___master_xactor_f_wr_resp___width { RTL___near_mem___icache___master_xactor_f_wr_resp___d0h }}& RTL___near_mem___icache___master_xactor_f_wr_resp___data0_reg ; 
                 RTL___near_mem___icache___master_xactor_f_wr_resp___data1_reg  <= RTL___near_mem___icache___master_xactor_f_wr_resp___d1di  ?  RTL___near_mem___icache___master_xactor_f_wr_resp___D_IN : RTL___near_mem___icache___master_xactor_f_wr_resp___data1_reg ;
             end 
         end
  always @( posedge  RTL___near_mem___icache___master_xactor_f_wr_resp___CLK )
         begin : RTL___near_mem___icache___master_xactor_f_wr_resp___error_checks 
           reg RTL___near_mem___icache___master_xactor_f_wr_resp___deqerror , RTL___near_mem___icache___master_xactor_f_wr_resp___enqerror ; 
             RTL___near_mem___icache___master_xactor_f_wr_resp___deqerror  =0; 
             RTL___near_mem___icache___master_xactor_f_wr_resp___enqerror  =0;
             if ( RTL___near_mem___icache___master_xactor_f_wr_resp___RST ==!1'b0)
                 begin 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg && RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ )
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_resp___deqerror  =1;$display("Warning: FIFO2: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg && RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ &&(! RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ || RTL___near_mem___icache___master_xactor_f_wr_resp___guarded ))
                         begin  
                             RTL___near_mem___icache___master_xactor_f_wr_resp___enqerror  =1;$display("Warning: FIFO2: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___full_reg ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___empty_reg ;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___D_IN = RTL___near_mem___dcache___f_fabric_write_reqs$D_IN;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___ENQ = RTL___near_mem___dcache___f_fabric_write_reqs$ENQ;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___DEQ = RTL___near_mem___dcache___f_fabric_write_reqs$DEQ;
    assign RTL___near_mem___dcache___f_fabric_write_reqs___CLR = RTL___near_mem___dcache___f_fabric_write_reqs$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___f_fabric_write_reqs$FULL_N = RTL___near_mem___dcache___f_fabric_write_reqs___FULL_N;
    assign RTL___near_mem___dcache___f_fabric_write_reqs$EMPTY_N = RTL___near_mem___dcache___f_fabric_write_reqs___EMPTY_N;
    assign RTL___near_mem___dcache___f_fabric_write_reqs$D_OUT = RTL___near_mem___dcache___f_fabric_write_reqs___D_OUT;
    assign RTL___near_mem___dcache___f_reset_reqs___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___f_reset_reqs___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___f_reset_reqs___D_IN = RTL___near_mem___dcache___f_reset_reqs$D_IN;
    assign RTL___near_mem___dcache___f_reset_reqs___ENQ = RTL___near_mem___dcache___f_reset_reqs$ENQ;
    assign RTL___near_mem___dcache___f_reset_reqs___DEQ = RTL___near_mem___dcache___f_reset_reqs$DEQ;
    assign RTL___near_mem___dcache___f_reset_reqs___CLR = RTL___near_mem___dcache___f_reset_reqs$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___CLK = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___dcache___f_reset_rsps$D_IN = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___f_reset_rsps$CLR = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___dcache___f_reset_rsps$D_OUT = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___dcache___f_reset_rsps$EMPTY_N = RTL___near_mem___dcache___f_reset_reqs___RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___dcache___f_reset_reqs$FULL_N = RTL___near_mem___dcache___f_reset_reqs___FULL_N;
    assign RTL___near_mem___dcache___f_reset_reqs$EMPTY_N = RTL___near_mem___dcache___f_reset_reqs___EMPTY_N;
    assign RTL___near_mem___dcache___f_reset_reqs$D_OUT = RTL___near_mem___dcache___f_reset_reqs___D_OUT;
    assign RTL___near_mem___dcache___f_reset_rsps___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___f_reset_rsps___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___f_reset_rsps___D_IN = RTL___near_mem___dcache___f_reset_rsps$D_IN;
    assign RTL___near_mem___dcache___f_reset_rsps___ENQ = RTL___near_mem___dcache___f_reset_rsps$ENQ;
    assign RTL___near_mem___dcache___f_reset_rsps___DEQ = RTL___near_mem___dcache___f_reset_rsps$DEQ;
    assign RTL___near_mem___dcache___f_reset_rsps___CLR = RTL___near_mem___dcache___f_reset_rsps$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___dcache___f_reset_rsps$FULL_N = RTL___near_mem___dcache___f_reset_rsps___FULL_N;
    assign RTL___near_mem___dcache___f_reset_rsps$EMPTY_N = RTL___near_mem___dcache___f_reset_rsps___EMPTY_N;
    assign RTL___near_mem___dcache___f_reset_rsps$D_OUT = RTL___near_mem___dcache___f_reset_rsps___D_OUT;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___D_IN = RTL___near_mem___dcache___master_xactor_f_rd_addr$D_IN;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___ENQ = RTL___near_mem___dcache___master_xactor_f_rd_addr$ENQ;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___DEQ = RTL___near_mem___dcache___master_xactor_f_rd_addr$DEQ;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr___CLR = RTL___near_mem___dcache___master_xactor_f_rd_addr$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr$FULL_N = RTL___near_mem___dcache___master_xactor_f_rd_addr___FULL_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr$EMPTY_N = RTL___near_mem___dcache___master_xactor_f_rd_addr___EMPTY_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_addr$D_OUT = RTL___near_mem___dcache___master_xactor_f_rd_addr___D_OUT;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___D_IN = RTL___near_mem___dcache___master_xactor_f_rd_data$D_IN;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___ENQ = RTL___near_mem___dcache___master_xactor_f_rd_data$ENQ;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___DEQ = RTL___near_mem___dcache___master_xactor_f_rd_data$DEQ;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data___CLR = RTL___near_mem___dcache___master_xactor_f_rd_data$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data$FULL_N = RTL___near_mem___dcache___master_xactor_f_rd_data___FULL_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data$EMPTY_N = RTL___near_mem___dcache___master_xactor_f_rd_data___EMPTY_N;
    assign RTL___near_mem___dcache___master_xactor_f_rd_data$D_OUT = RTL___near_mem___dcache___master_xactor_f_rd_data___D_OUT;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___D_IN = RTL___near_mem___dcache___master_xactor_f_wr_addr$D_IN;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___ENQ = RTL___near_mem___dcache___master_xactor_f_wr_addr$ENQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___DEQ = RTL___near_mem___dcache___master_xactor_f_wr_addr$DEQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr___CLR = RTL___near_mem___dcache___master_xactor_f_wr_addr$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr$FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_addr___FULL_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr$EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_addr___EMPTY_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_addr$D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_addr___D_OUT;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___D_IN = RTL___near_mem___dcache___master_xactor_f_wr_data$D_IN;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___ENQ = RTL___near_mem___dcache___master_xactor_f_wr_data$ENQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___DEQ = RTL___near_mem___dcache___master_xactor_f_wr_data$DEQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data___CLR = RTL___near_mem___dcache___master_xactor_f_wr_data$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data$FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_data___FULL_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data$EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_data___EMPTY_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_data$D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_data___D_OUT;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___RST = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___D_IN = RTL___near_mem___dcache___master_xactor_f_wr_resp$D_IN;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___ENQ = RTL___near_mem___dcache___master_xactor_f_wr_resp$ENQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___DEQ = RTL___near_mem___dcache___master_xactor_f_wr_resp$DEQ;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp___CLR = RTL___near_mem___dcache___master_xactor_f_wr_resp$CLR;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp$FULL_N = RTL___near_mem___dcache___master_xactor_f_wr_resp___FULL_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp$EMPTY_N = RTL___near_mem___dcache___master_xactor_f_wr_resp___EMPTY_N;
    assign RTL___near_mem___dcache___master_xactor_f_wr_resp$D_OUT = RTL___near_mem___dcache___master_xactor_f_wr_resp___D_OUT;
    assign RTL___near_mem___icache___f_fabric_write_reqs___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___f_fabric_write_reqs___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___f_fabric_write_reqs___D_IN = RTL___near_mem___icache___f_fabric_write_reqs$D_IN;
    assign RTL___near_mem___icache___f_fabric_write_reqs___ENQ = RTL___near_mem___icache___f_fabric_write_reqs$ENQ;
    assign RTL___near_mem___icache___f_fabric_write_reqs___DEQ = RTL___near_mem___icache___f_fabric_write_reqs$DEQ;
    assign RTL___near_mem___icache___f_fabric_write_reqs___CLR = RTL___near_mem___icache___f_fabric_write_reqs$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___f_fabric_write_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___icache___f_fabric_write_reqs$FULL_N = RTL___near_mem___icache___f_fabric_write_reqs___FULL_N;
    assign RTL___near_mem___icache___f_fabric_write_reqs$EMPTY_N = RTL___near_mem___icache___f_fabric_write_reqs___EMPTY_N;
    assign RTL___near_mem___icache___f_fabric_write_reqs$D_OUT = RTL___near_mem___icache___f_fabric_write_reqs___D_OUT;
    assign RTL___near_mem___icache___f_reset_reqs___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___f_reset_reqs___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___f_reset_reqs___D_IN = RTL___near_mem___icache___f_reset_reqs$D_IN;
    assign RTL___near_mem___icache___f_reset_reqs___ENQ = RTL___near_mem___icache___f_reset_reqs$ENQ;
    assign RTL___near_mem___icache___f_reset_reqs___DEQ = RTL___near_mem___icache___f_reset_reqs$DEQ;
    assign RTL___near_mem___icache___f_reset_reqs___CLR = RTL___near_mem___icache___f_reset_reqs$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___icache___RST_N = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___f_reset_reqs___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___icache___f_reset_reqs$FULL_N = RTL___near_mem___icache___f_reset_reqs___FULL_N;
    assign RTL___near_mem___icache___f_reset_reqs$EMPTY_N = RTL___near_mem___icache___f_reset_reqs___EMPTY_N;
    assign RTL___near_mem___icache___f_reset_reqs$D_OUT = RTL___near_mem___icache___f_reset_reqs___D_OUT;
    assign RTL___near_mem___icache___f_reset_rsps___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___f_reset_rsps___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___f_reset_rsps___D_IN = RTL___near_mem___icache___f_reset_rsps$D_IN;
    assign RTL___near_mem___icache___f_reset_rsps___ENQ = RTL___near_mem___icache___f_reset_rsps$ENQ;
    assign RTL___near_mem___icache___f_reset_rsps___DEQ = RTL___near_mem___icache___f_reset_rsps$DEQ;
    assign RTL___near_mem___icache___f_reset_rsps___CLR = RTL___near_mem___icache___f_reset_rsps$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___f_reset_rsps___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___icache___f_reset_rsps$FULL_N = RTL___near_mem___icache___f_reset_rsps___FULL_N;
    assign RTL___near_mem___icache___f_reset_rsps$EMPTY_N = RTL___near_mem___icache___f_reset_rsps___EMPTY_N;
    assign RTL___near_mem___icache___f_reset_rsps$D_OUT = RTL___near_mem___icache___f_reset_rsps___D_OUT;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___D_IN = RTL___near_mem___icache___master_xactor_f_rd_addr$D_IN;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___ENQ = RTL___near_mem___icache___master_xactor_f_rd_addr$ENQ;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___DEQ = RTL___near_mem___icache___master_xactor_f_rd_addr$DEQ;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr___CLR = RTL___near_mem___icache___master_xactor_f_rd_addr$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr$FULL_N = RTL___near_mem___icache___master_xactor_f_rd_addr___FULL_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr$EMPTY_N = RTL___near_mem___icache___master_xactor_f_rd_addr___EMPTY_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_addr$D_OUT = RTL___near_mem___icache___master_xactor_f_rd_addr___D_OUT;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___D_IN = RTL___near_mem___icache___master_xactor_f_rd_data$D_IN;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___ENQ = RTL___near_mem___icache___master_xactor_f_rd_data$ENQ;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___DEQ = RTL___near_mem___icache___master_xactor_f_rd_data$DEQ;
    assign RTL___near_mem___icache___master_xactor_f_rd_data___CLR = RTL___near_mem___icache___master_xactor_f_rd_data$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_rd_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___icache___master_xactor_f_rd_data$FULL_N = RTL___near_mem___icache___master_xactor_f_rd_data___FULL_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_data$EMPTY_N = RTL___near_mem___icache___master_xactor_f_rd_data___EMPTY_N;
    assign RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT = RTL___near_mem___icache___master_xactor_f_rd_data___D_OUT;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___D_IN = RTL___near_mem___icache___master_xactor_f_wr_addr$D_IN;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___ENQ = RTL___near_mem___icache___master_xactor_f_wr_addr$ENQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___DEQ = RTL___near_mem___icache___master_xactor_f_wr_addr$DEQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr___CLR = RTL___near_mem___icache___master_xactor_f_wr_addr$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_addr___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr$FULL_N = RTL___near_mem___icache___master_xactor_f_wr_addr___FULL_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr$EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_addr___EMPTY_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_addr$D_OUT = RTL___near_mem___icache___master_xactor_f_wr_addr___D_OUT;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___D_IN = RTL___near_mem___icache___master_xactor_f_wr_data$D_IN;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___ENQ = RTL___near_mem___icache___master_xactor_f_wr_data$ENQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___DEQ = RTL___near_mem___icache___master_xactor_f_wr_data$DEQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_data___CLR = RTL___near_mem___icache___master_xactor_f_wr_data$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_data___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___icache___master_xactor_f_wr_data$FULL_N = RTL___near_mem___icache___master_xactor_f_wr_data___FULL_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_data$EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_data___EMPTY_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_data$D_OUT = RTL___near_mem___icache___master_xactor_f_wr_data___D_OUT;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___RST = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___D_IN = RTL___near_mem___icache___master_xactor_f_wr_resp$D_IN;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___ENQ = RTL___near_mem___icache___master_xactor_f_wr_resp$ENQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___DEQ = RTL___near_mem___icache___master_xactor_f_wr_resp$DEQ;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp___CLR = RTL___near_mem___icache___master_xactor_f_wr_resp$CLR;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___master_xactor_f_wr_resp___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp$FULL_N = RTL___near_mem___icache___master_xactor_f_wr_resp___FULL_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp$EMPTY_N = RTL___near_mem___icache___master_xactor_f_wr_resp___EMPTY_N;
    assign RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT = RTL___near_mem___icache___master_xactor_f_wr_resp___D_OUT;
      
    
    reg[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R ; reg[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R ; reg[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R2 ; reg[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R2 ; 
    wire[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___arb1 ; 
    wire[ RTL___near_mem___icache___ram_state_and_ctag_cset___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_state_and_ctag_cset___arb2 ; 
  always @( posedge  RTL___near_mem___icache___ram_state_and_ctag_cset___CLKA )
         begin 
             if ( RTL___near_mem___icache___ram_state_and_ctag_cset___ENA )
                 begin 
                     if ( RTL___near_mem___icache___ram_state_and_ctag_cset___WEA )
                         begin  
                             RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R  <= RTL___near_mem___icache___ram_state_and_ctag_cset___DIA ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R  <= RTL___near_mem___icache___ram_state_and_ctag_cset___arb1 ;
                         end 
                 end  
             RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R2  <= RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R ;
         end
  always @( posedge  RTL___near_mem___icache___ram_state_and_ctag_cset___CLKB )
         begin 
             if ( RTL___near_mem___icache___ram_state_and_ctag_cset___ENB )
                 begin 
                     if ( RTL___near_mem___icache___ram_state_and_ctag_cset___WEB )
                         begin  
                             RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R  <= RTL___near_mem___icache___ram_state_and_ctag_cset___DIB ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R  <= RTL___near_mem___icache___ram_state_and_ctag_cset___arb2 ;
                         end 
                 end  
             RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R2  <= RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R ;
         end
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset___DOA =( RTL___near_mem___icache___ram_state_and_ctag_cset___PIPELINED ) ?  RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R2 : RTL___near_mem___icache___ram_state_and_ctag_cset___DOA_R ; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset___DOB =( RTL___near_mem___icache___ram_state_and_ctag_cset___PIPELINED ) ?  RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R2 : RTL___near_mem___icache___ram_state_and_ctag_cset___DOB_R ;
    reg[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___DOA_R ; reg[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___DOB_R ; reg[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___DOA_R2 ; reg[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___DOB_R2 ; 
    wire[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___arb1 ; 
    wire[ RTL___near_mem___icache___ram_word64_set___DATA_WIDTH -1:0] RTL___near_mem___icache___ram_word64_set___arb2 ; 
  always @( posedge  RTL___near_mem___icache___ram_word64_set___CLKA )
         begin 
             if ( RTL___near_mem___icache___ram_word64_set___ENA )
                 begin 
                     if ( RTL___near_mem___icache___ram_word64_set___WEA )
                         begin  
                             RTL___near_mem___icache___ram_word64_set___DOA_R  <= RTL___near_mem___icache___ram_word64_set___DIA ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___icache___ram_word64_set___DOA_R  <= RTL___near_mem___icache___ram_word64_set___arb1 ;
                         end 
                 end  
             RTL___near_mem___icache___ram_word64_set___DOA_R2  <= RTL___near_mem___icache___ram_word64_set___DOA_R ;
         end
  always @( posedge  RTL___near_mem___icache___ram_word64_set___CLKB )
         begin 
             if ( RTL___near_mem___icache___ram_word64_set___ENB )
                 begin 
                     if ( RTL___near_mem___icache___ram_word64_set___WEB )
                         begin  
                             RTL___near_mem___icache___ram_word64_set___DOB_R  <= RTL___near_mem___icache___ram_word64_set___DIB ;
                         end 
                      else 
                         begin  
                             RTL___near_mem___icache___ram_word64_set___DOB_R  <= RTL___near_mem___icache___ram_word64_set___arb2 ;
                         end 
                 end  
             RTL___near_mem___icache___ram_word64_set___DOB_R2  <= RTL___near_mem___icache___ram_word64_set___DOB_R ;
         end
  assign  RTL___near_mem___icache___ram_word64_set___DOA =( RTL___near_mem___icache___ram_word64_set___PIPELINED ) ?  RTL___near_mem___icache___ram_word64_set___DOA_R2 : RTL___near_mem___icache___ram_word64_set___DOA_R ; 
  assign  RTL___near_mem___icache___ram_word64_set___DOB =( RTL___near_mem___icache___ram_word64_set___PIPELINED ) ?  RTL___near_mem___icache___ram_word64_set___DOB_R2 : RTL___near_mem___icache___ram_word64_set___DOB_R ;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKA = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___ENA = RTL___near_mem___dcache___ram_state_and_ctag_cset$ENA;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___WEA = RTL___near_mem___dcache___ram_state_and_ctag_cset$WEA;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDRA = RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRA;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___DIA = RTL___near_mem___dcache___ram_state_and_ctag_cset$DIA;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___CLKB = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___ENB = RTL___near_mem___dcache___ram_state_and_ctag_cset$ENB;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___WEB = RTL___near_mem___dcache___ram_state_and_ctag_cset$WEB;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___ADDRB = RTL___near_mem___dcache___ram_state_and_ctag_cset$ADDRB;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset___DIB = RTL___near_mem___dcache___ram_state_and_ctag_cset$DIB;
    assign RTL___near_mem___dcache___ram_state_and_ctag_cset$DOB = RTL___near_mem___dcache___ram_state_and_ctag_cset___DOB;
    assign RTL___near_mem___dcache___ram_word64_set___CLKA = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___ram_word64_set___ENA = RTL___near_mem___dcache___ram_word64_set$ENA;
    assign RTL___near_mem___dcache___ram_word64_set___WEA = RTL___near_mem___dcache___ram_word64_set$WEA;
    assign RTL___near_mem___dcache___ram_word64_set___ADDRA = RTL___near_mem___dcache___ram_word64_set$ADDRA;
    assign RTL___near_mem___dcache___ram_word64_set___DIA = RTL___near_mem___dcache___ram_word64_set$DIA;
    assign RTL___near_mem___dcache___ram_word64_set___CLKB = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___ram_word64_set___ENB = RTL___near_mem___dcache___ram_word64_set$ENB;
    assign RTL___near_mem___dcache___ram_word64_set___WEB = RTL___near_mem___dcache___ram_word64_set$WEB;
    assign RTL___near_mem___dcache___ram_word64_set___ADDRB = RTL___near_mem___dcache___ram_word64_set$ADDRB;
    assign RTL___near_mem___dcache___ram_word64_set___DIB = RTL___near_mem___dcache___ram_word64_set$DIB;
    assign RTL___near_mem___dcache___ram_word64_set$DOB = RTL___near_mem___dcache___ram_word64_set___DOB;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___CLKA = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___ENA = RTL___near_mem___icache___ram_state_and_ctag_cset$ENA;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___WEA = RTL___near_mem___icache___ram_state_and_ctag_cset$WEA;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___ADDRA = RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRA;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___DIA = RTL___near_mem___icache___ram_state_and_ctag_cset$DIA;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___CLKB = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___ENB = RTL___near_mem___icache___ram_state_and_ctag_cset$ENB;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___WEB = RTL___near_mem___icache___ram_state_and_ctag_cset$WEB;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___ADDRB = RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRB;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset___DIB = RTL___near_mem___icache___ram_state_and_ctag_cset$DIB;
    assign RTL___near_mem___icache___ram_state_and_ctag_cset$DOB = RTL___near_mem___icache___ram_state_and_ctag_cset___DOB;
    assign RTL___near_mem___icache___ram_word64_set___CLKA = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___ram_word64_set___ENA = RTL___near_mem___icache___ram_word64_set$ENA;
    assign RTL___near_mem___icache___ram_word64_set___WEA = RTL___near_mem___icache___ram_word64_set$WEA;
    assign RTL___near_mem___icache___ram_word64_set___ADDRA = RTL___near_mem___icache___ram_word64_set$ADDRA;
    assign RTL___near_mem___icache___ram_word64_set___DIA = RTL___near_mem___icache___ram_word64_set$DIA;
    assign RTL___near_mem___icache___ram_word64_set___CLKB = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___ram_word64_set___ENB = RTL___near_mem___icache___ram_word64_set$ENB;
    assign RTL___near_mem___icache___ram_word64_set___WEB = RTL___near_mem___icache___ram_word64_set$WEB;
    assign RTL___near_mem___icache___ram_word64_set___ADDRB = RTL___near_mem___icache___ram_word64_set$ADDRB;
    assign RTL___near_mem___icache___ram_word64_set___DIB = RTL___near_mem___icache___ram_word64_set$DIB;
    assign RTL___near_mem___icache___ram_word64_set$DOB = RTL___near_mem___icache___ram_word64_set___DOB;
      
    
    wire[63:0] RTL___near_mem___icache___soc_map___m_boot_rom_addr_base , RTL___near_mem___icache___soc_map___m_boot_rom_addr_lim , RTL___near_mem___icache___soc_map___m_boot_rom_addr_size , RTL___near_mem___icache___soc_map___m_mem0_controller_addr_base , RTL___near_mem___icache___soc_map___m_mem0_controller_addr_lim , RTL___near_mem___icache___soc_map___m_mem0_controller_addr_size , RTL___near_mem___icache___soc_map___m_mtvec_reset_value , RTL___near_mem___icache___soc_map___m_near_mem_io_addr_base , RTL___near_mem___icache___soc_map___m_near_mem_io_addr_lim , RTL___near_mem___icache___soc_map___m_near_mem_io_addr_size , RTL___near_mem___icache___soc_map___m_nmivec_reset_value , RTL___near_mem___icache___soc_map___m_pc_reset_value , RTL___near_mem___icache___soc_map___m_plic_addr_base , RTL___near_mem___icache___soc_map___m_plic_addr_lim , RTL___near_mem___icache___soc_map___m_plic_addr_size , RTL___near_mem___icache___soc_map___m_tcm_addr_base , RTL___near_mem___icache___soc_map___m_tcm_addr_lim , RTL___near_mem___icache___soc_map___m_tcm_addr_size , RTL___near_mem___icache___soc_map___m_uart0_addr_base , RTL___near_mem___icache___soc_map___m_uart0_addr_lim , RTL___near_mem___icache___soc_map___m_uart0_addr_size ; 
    wire RTL___near_mem___icache___soc_map___m_is_IO_addr , RTL___near_mem___icache___soc_map___m_is_mem_addr , RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr ; 
  assign  RTL___near_mem___icache___soc_map___m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL___near_mem___icache___soc_map___m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL___near_mem___icache___soc_map___m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL___near_mem___icache___soc_map___m_plic_addr_base =64'h000000000C000000; 
  assign  RTL___near_mem___icache___soc_map___m_plic_addr_size =64'h0000000000400000; 
  assign  RTL___near_mem___icache___soc_map___m_plic_addr_lim =64'd205520896; 
  assign  RTL___near_mem___icache___soc_map___m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL___near_mem___icache___soc_map___m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL___near_mem___icache___soc_map___m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL___near_mem___icache___soc_map___m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL___near_mem___icache___soc_map___m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL___near_mem___icache___soc_map___m_boot_rom_addr_lim =64'd8192; 
  assign  RTL___near_mem___icache___soc_map___m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL___near_mem___icache___soc_map___m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL___near_mem___icache___soc_map___m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL___near_mem___icache___soc_map___m_tcm_addr_base =64'h0; 
  assign  RTL___near_mem___icache___soc_map___m_tcm_addr_size =64'd0; 
  assign  RTL___near_mem___icache___soc_map___m_tcm_addr_lim =64'd0; 
  assign  RTL___near_mem___icache___soc_map___m_is_mem_addr = RTL___near_mem___icache___soc_map___m_is_mem_addr_addr >=64'h0000000000001000&& RTL___near_mem___icache___soc_map___m_is_mem_addr_addr <64'd8192|| RTL___near_mem___icache___soc_map___m_is_mem_addr_addr >=64'h0000000080000000&& RTL___near_mem___icache___soc_map___m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL___near_mem___icache___soc_map___m_is_IO_addr = RTL___near_mem___icache___soc_map___m_is_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___icache___soc_map___m_is_IO_addr_addr <64'd33603584|| RTL___near_mem___icache___soc_map___m_is_IO_addr_addr >=64'h000000000C000000&& RTL___near_mem___icache___soc_map___m_is_IO_addr_addr <64'd205520896|| RTL___near_mem___icache___soc_map___m_is_IO_addr_addr >=64'h00000000C0000000&& RTL___near_mem___icache___soc_map___m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr = RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL___near_mem___icache___soc_map___m_pc_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___icache___soc_map___m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___icache___soc_map___m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
     
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req = RTL___near_mem___icache___f_fabric_write_reqs$EMPTY_N && RTL___near_mem___icache___master_xactor_f_wr_addr$FULL_N && RTL___near_mem___icache___master_xactor_f_wr_data$FULL_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req = RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_reset =( RTL___near_mem___icache___rg_cset_in_cache !=7'd127|| RTL___near_mem___icache___f_reset_reqs$EMPTY_N && RTL___near_mem___icache___f_reset_rsps$FULL_N )&& RTL___near_mem___icache___rg_state ==4'd1; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_reset = RTL___near_mem___icache___CAN_FIRE_RL_rl_reset ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_probe_and_immed_rsp =( RTL___near_mem___icache___dmem_not_imem &&! RTL___near_mem___icache___soc_map$m_is_mem_addr ||! RTL___near_mem___icache___rg_op || RTL___near_mem___icache___f_fabric_write_reqs$FULL_N )&& RTL___near_mem___icache___rg_state ==4'd3; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp = RTL___near_mem___icache___CAN_FIRE_RL_rl_probe_and_immed_rsp &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_start_cache_refill = RTL___near_mem___icache___master_xactor_f_rd_addr$FULL_N && RTL___near_mem___icache___rg_state ==4'd8&& RTL___near_mem___icache___b__h14485 ==4'd0; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill = RTL___near_mem___icache___CAN_FIRE_RL_rl_start_cache_refill &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_cache_refill_rsps_loop = RTL___near_mem___icache___master_xactor_f_rd_data$EMPTY_N && RTL___near_mem___icache___rg_state ==4'd9; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop = RTL___near_mem___icache___CAN_FIRE_RL_rl_cache_refill_rsps_loop &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_rereq = RTL___near_mem___icache___rg_state ==4'd10; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq = RTL___near_mem___icache___CAN_FIRE_RL_rl_rereq &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_ST_AMO_response = RTL___near_mem___icache___rg_state ==4'd11; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_ST_AMO_response = RTL___near_mem___icache___CAN_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_req = RTL___near_mem___icache___master_xactor_f_rd_addr$FULL_N && RTL___near_mem___icache___rg_state ==4'd12&&! RTL___near_mem___icache___rg_op && RTL___near_mem___icache___b__h14485 ==4'd0; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req = RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_req &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_rsp = RTL___near_mem___icache___master_xactor_f_rd_data$EMPTY_N && RTL___near_mem___icache___rg_state ==4'd13; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp = RTL___near_mem___icache___CAN_FIRE_RL_rl_io_read_rsp &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_maintain_io_read_rsp = RTL___near_mem___icache___rg_state ==4'd14; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp = RTL___near_mem___icache___CAN_FIRE_RL_rl_maintain_io_read_rsp ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_io_write_req = RTL___near_mem___icache___f_fabric_write_reqs$FULL_N && RTL___near_mem___icache___rg_state ==4'd12&& RTL___near_mem___icache___rg_op ; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req = RTL___near_mem___icache___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_discard_write_rsp = RTL___near_mem___icache___b__h14485 !=4'd0&& RTL___near_mem___icache___master_xactor_f_wr_resp$EMPTY_N ; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp = RTL___near_mem___icache___CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_drive_exception_rsp = RTL___near_mem___icache___rg_state ==4'd4; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_drive_exception_rsp = RTL___near_mem___icache___rg_state ==4'd4; 
  assign  RTL___near_mem___icache___CAN_FIRE_RL_rl_start_reset = RTL___near_mem___icache___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset = RTL___near_mem___icache___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_1 = RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_2 = RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 ; 
  assign  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__SEL_3 = RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL___near_mem___icache___WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__SEL_1 = RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op ; 
  assign  RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1 = RTL___near_mem___icache___EN_req && RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 ; 
  assign  RTL___near_mem___icache___MUX_ram_word64_set$a_put_1__SEL_1 = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0; 
  assign  RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2 = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]!=2'd3; 
  assign  RTL___near_mem___icache___MUX_rg_error_during_refill$write_1__SEL_1 = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_1 = RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_2 = RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__SEL_2 = RTL___near_mem___icache___f_reset_reqs$EMPTY_N && RTL___near_mem___icache___rg_state !=4'd1; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__SEL_3 = RTL___near_mem___icache___CAN_FIRE_RL_rl_io_write_req &&! RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__SEL_7 = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]==2'd3; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__SEL_9 = RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 ; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__SEL_10 = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127; 
  always @(          RTL___near_mem___icache___rg_f3                          or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247                 or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276                or   RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32               or   RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___word64__h5094             or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264            or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285           or   RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  )
         begin 
             case ( RTL___near_mem___icache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247 ;
              3 'b001: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276 ;
              3 'b010: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32 ;
              3 'b011: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  =( RTL___near_mem___icache___rg_addr [2:0]==3'h0) ?  RTL___near_mem___icache___word64__h5094 :64'd0;
              3 'b100: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264 ;
              3 'b101: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285 ;
              3 'b110: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  = RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33 ;
              3 'd7: 
                  RTL___near_mem___icache___MUX_dw_output_ld_val$wset_1__VAL_2  =64'd0;endcase
         end
  assign  RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_1 ={ RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_st_amo_val }; 
  assign  RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ={ RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_pa , RTL___near_mem___icache___rg_st_amo_val }; 
  assign  RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 ={4'd0, RTL___near_mem___icache___cline_fabric_addr__h14584 ,29'd7143424}; 
  assign  RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ={4'd0, RTL___near_mem___icache___fabric_addr__h17243 ,8'd0, RTL___near_mem___icache___value__h17372 ,18'd65536}; 
  assign  RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 ={3'd4, RTL___near_mem___icache___rg_pa [31:12]}; 
  assign  RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_2 = RTL___near_mem___icache___rg_word64_set_in_cache +9'd1; 
  assign  RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_4 ={ RTL___near_mem___icache___rg_addr [11:5],2'd0}; 
  assign  RTL___near_mem___icache___MUX_rg_cset_in_cache$write_1__VAL_1 = RTL___near_mem___icache___rg_cset_in_cache +7'd1; 
  assign  RTL___near_mem___icache___MUX_rg_exc_code$write_1__VAL_1 = RTL___near_mem___icache___req_op  ? 4'd6:4'd4; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__VAL_1 = RTL___near_mem___icache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539  ? 4'd4:4'd3; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__VAL_4 =( RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0) ? 4'd14:4'd4; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__VAL_7 =( RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___icache___rg_error_during_refill ) ? 4'd4:4'd10; 
  assign  RTL___near_mem___icache___MUX_rg_state$write_1__VAL_9 =( RTL___near_mem___icache___dmem_not_imem &&! RTL___near_mem___icache___soc_map$m_is_mem_addr ) ? 4'd12:( RTL___near_mem___icache___rg_op  ? 4'd11:4'd8); 
  assign  RTL___near_mem___icache___dw_valid$whas = RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 || RTL___near_mem___icache___WILL_FIRE_RL_rl_drive_exception_rsp || RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp || RTL___near_mem___icache___WILL_FIRE_RL_rl_ST_AMO_response ; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port0__write_1 = RTL___near_mem___icache___ctr_wr_rsps_pending_crg +4'd1; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port1__write_1 = RTL___near_mem___icache___b__h14485 -4'd1; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port2__read = RTL___near_mem___icache___CAN_FIRE_RL_rl_discard_write_rsp  ?  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port1__write_1 : RTL___near_mem___icache___b__h14485 ; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN_port2__write = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port3__read = RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN_port2__write  ? 4'd0: RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port2__read ; 
  assign  RTL___near_mem___icache___cfg_verbosity$D_IN = RTL___near_mem___icache___set_verbosity_verbosity ; 
  assign  RTL___near_mem___icache___cfg_verbosity$EN = RTL___near_mem___icache___EN_set_verbosity ; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$D_IN = RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port3__read ; 
  assign  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN =1'b1; 
  assign  RTL___near_mem___icache___rg_addr$D_IN = RTL___near_mem___icache___req_addr ; 
  assign  RTL___near_mem___icache___rg_addr$EN = RTL___near_mem___icache___EN_req ; 
    wire[6:0] RTL___near_mem___icache___MUX_rg_cset_in_cache$write_1__VAL_1_any_val ; 
  assign  RTL___near_mem___icache___rg_cset_in_cache$D_IN = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset  ?  RTL___near_mem___icache___MUX_rg_cset_in_cache$write_1__VAL_1_any_val :7'd0; 
  assign  RTL___near_mem___icache___rg_cset_in_cache$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset || RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___rg_error_during_refill$D_IN = RTL___near_mem___icache___MUX_rg_error_during_refill$write_1__SEL_1 ; 
  assign  RTL___near_mem___icache___rg_error_during_refill$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill ; 
  always @(      RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_1                  or   RTL___near_mem___icache___MUX_rg_exc_code$write_1__VAL_1             or   RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_2            or   RTL___near_mem___icache___MUX_rg_error_during_refill$write_1__SEL_1           or   RTL___near_mem___icache___access_exc_code__h2256  )
         case (1'b1) 
          RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_1  : 
              RTL___near_mem___icache___rg_exc_code$D_IN  = RTL___near_mem___icache___MUX_rg_exc_code$write_1__VAL_1 ; 
          RTL___near_mem___icache___MUX_rg_exc_code$write_1__SEL_2  : 
              RTL___near_mem___icache___rg_exc_code$D_IN  =4'd5; 
          RTL___near_mem___icache___MUX_rg_error_during_refill$write_1__SEL_1  : 
              RTL___near_mem___icache___rg_exc_code$D_IN  = RTL___near_mem___icache___access_exc_code__h2256 ;
          default : 
              RTL___near_mem___icache___rg_exc_code$D_IN  =4'b1010;endcase
  assign  RTL___near_mem___icache___rg_exc_code$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 ; 
  assign  RTL___near_mem___icache___rg_f3$D_IN = RTL___near_mem___icache___req_f3 ; 
  assign  RTL___near_mem___icache___rg_f3$EN = RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___rg_ld_val$D_IN = RTL___near_mem___icache___ld_val__h17594 ; 
  assign  RTL___near_mem___icache___rg_ld_val$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp ; 
  assign  RTL___near_mem___icache___rg_lower_word32$D_IN =32'h0; 
  assign  RTL___near_mem___icache___rg_lower_word32$EN =1'b0; 
  assign  RTL___near_mem___icache___rg_lower_word32_full$D_IN =1'd0; 
  assign  RTL___near_mem___icache___rg_lower_word32_full$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset ; 
  assign  RTL___near_mem___icache___rg_op$D_IN = RTL___near_mem___icache___req_op ; 
  assign  RTL___near_mem___icache___rg_op$EN = RTL___near_mem___icache___EN_req ; 
  assign  RTL___near_mem___icache___rg_pa$D_IN = RTL___near_mem___icache___EN_req  ?  RTL___near_mem___icache___req_addr : RTL___near_mem___icache___rg_addr ; 
  assign  RTL___near_mem___icache___rg_pa$EN = RTL___near_mem___icache___EN_req || RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp ; 
  assign  RTL___near_mem___icache___rg_pte_pa$D_IN =32'h0; 
  assign  RTL___near_mem___icache___rg_pte_pa$EN =1'b0; 
  assign  RTL___near_mem___icache___rg_st_amo_val$D_IN = RTL___near_mem___icache___req_st_value ; 
  assign  RTL___near_mem___icache___rg_st_amo_val$EN = RTL___near_mem___icache___EN_req ; 
  always @(               RTL___near_mem___icache___EN_req                                    or   RTL___near_mem___icache___MUX_rg_state$write_1__VAL_1                      or   RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset                     or   RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req                    or   RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp                   or   RTL___near_mem___icache___MUX_rg_state$write_1__VAL_4                  or   RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req                 or   RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq                or   RTL___near_mem___icache___MUX_rg_state$write_1__SEL_7               or   RTL___near_mem___icache___MUX_rg_state$write_1__VAL_7              or   RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill             or   RTL___near_mem___icache___MUX_rg_state$write_1__SEL_9            or   RTL___near_mem___icache___MUX_rg_state$write_1__VAL_9           or   RTL___near_mem___icache___MUX_rg_state$write_1__SEL_10  )
         case (1'b1) 
          RTL___near_mem___icache___EN_req  : 
              RTL___near_mem___icache___rg_state$D_IN  = RTL___near_mem___icache___MUX_rg_state$write_1__VAL_1 ; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd1; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd11; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp  : 
              RTL___near_mem___icache___rg_state$D_IN  = RTL___near_mem___icache___MUX_rg_state$write_1__VAL_4 ; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd13; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd3; 
          RTL___near_mem___icache___MUX_rg_state$write_1__SEL_7  : 
              RTL___near_mem___icache___rg_state$D_IN  = RTL___near_mem___icache___MUX_rg_state$write_1__VAL_7 ; 
          RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd9; 
          RTL___near_mem___icache___MUX_rg_state$write_1__SEL_9  : 
              RTL___near_mem___icache___rg_state$D_IN  = RTL___near_mem___icache___MUX_rg_state$write_1__VAL_9 ; 
          RTL___near_mem___icache___MUX_rg_state$write_1__SEL_10  : 
              RTL___near_mem___icache___rg_state$D_IN  =4'd2;
          default : 
              RTL___near_mem___icache___rg_state$D_IN  =4'b1010;endcase
  assign  RTL___near_mem___icache___rg_state$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127|| RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]==2'd3|| RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 || RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp || RTL___near_mem___icache___EN_req || RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset || RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq || RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req || RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL___near_mem___icache___rg_word64_set_in_cache$D_IN = RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2  ?  RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_2 : RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_4 ; 
  assign  RTL___near_mem___icache___rg_word64_set_in_cache$EN = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]!=2'd3|| RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs$D_IN = RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__SEL_1  ?  RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_1 : RTL___near_mem___icache___MUX_f_fabric_write_reqs$enq_1__VAL_2 ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs$ENQ = RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op || RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs$DEQ = RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___icache___f_fabric_write_reqs$CLR =1'b0; 
  assign  RTL___near_mem___icache___f_reset_reqs$D_IN =! RTL___near_mem___icache___EN_server_reset_request_put ; 
  assign  RTL___near_mem___icache___f_reset_reqs$ENQ = RTL___near_mem___icache___EN_server_reset_request_put || RTL___near_mem___icache___EN_server_flush_request_put ; 
  assign  RTL___near_mem___icache___f_reset_reqs$DEQ = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127; 
  assign  RTL___near_mem___icache___f_reset_reqs$CLR =1'b0; 
  assign  RTL___near_mem___icache___f_reset_rsps$D_IN = RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___f_reset_rsps$ENQ = RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127; 
  assign  RTL___near_mem___icache___f_reset_rsps$DEQ = RTL___near_mem___icache___EN_server_flush_response_get || RTL___near_mem___icache___EN_server_reset_response_get ; 
  assign  RTL___near_mem___icache___f_reset_rsps$CLR =1'b0; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr$D_IN = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_1 : RTL___near_mem___icache___MUX_master_xactor_f_rd_addr$enq_1__VAL_2 ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr$ENQ = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr$DEQ = RTL___near_mem___icache___master_xactor_f_rd_addr$EMPTY_N && RTL___near_mem___icache___mem_master_arready ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_addr$CLR = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data$D_IN ={ RTL___near_mem___icache___mem_master_rid , RTL___near_mem___icache___mem_master_rdata , RTL___near_mem___icache___mem_master_rresp , RTL___near_mem___icache___mem_master_rlast }; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data$ENQ = RTL___near_mem___icache___mem_master_rvalid && RTL___near_mem___icache___master_xactor_f_rd_data$FULL_N ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data$DEQ = RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp || RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop ; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_data$CLR = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr$D_IN ={4'd0, RTL___near_mem___icache___mem_req_wr_addr_awaddr__h2473 ,8'd0, RTL___near_mem___icache___x__h2520 ,18'd65536}; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr$ENQ = RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr$DEQ = RTL___near_mem___icache___master_xactor_f_wr_addr$EMPTY_N && RTL___near_mem___icache___mem_master_awready ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_addr$CLR = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data$D_IN ={ RTL___near_mem___icache___mem_req_wr_data_wdata__h2699 , RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700 ,1'd1}; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data$ENQ = RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data$DEQ = RTL___near_mem___icache___master_xactor_f_wr_data$EMPTY_N && RTL___near_mem___icache___mem_master_wready ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_data$CLR = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp$D_IN ={ RTL___near_mem___icache___mem_master_bid , RTL___near_mem___icache___mem_master_bresp }; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp$ENQ = RTL___near_mem___icache___mem_master_bvalid && RTL___near_mem___icache___master_xactor_f_wr_resp$FULL_N ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp$DEQ = RTL___near_mem___icache___CAN_FIRE_RL_rl_discard_write_rsp ; 
  assign  RTL___near_mem___icache___master_xactor_f_wr_resp$CLR = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset &&! RTL___near_mem___icache___f_reset_reqs$D_OUT ; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRA = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___icache___rg_addr [11:5]: RTL___near_mem___icache___rg_cset_in_cache ; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$ADDRB = RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ?  RTL___near_mem___icache___req_addr [11:5]: RTL___near_mem___icache___rg_addr [11:5]; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$DIA = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  ?  RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$a_put_3__VAL_1 :23'd2796202; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$DIB = RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  ? 23'b01010101010101010101010:23'b01010101010101010101010; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$WEA =1'd1; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$WEB =1'd0; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$ENA = RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill || RTL___near_mem___icache___WILL_FIRE_RL_rl_reset ; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset$ENB = RTL___near_mem___icache___EN_req && RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq ; 
  assign  RTL___near_mem___icache___ram_word64_set$ADDRA = RTL___near_mem___icache___MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL___near_mem___icache___rg_word64_set_in_cache : RTL___near_mem___icache___rg_addr [11:3]; 
  always @(         RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                        or   RTL___near_mem___icache___req_addr                or   RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2               or   RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_2              or   RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq             or   RTL___near_mem___icache___rg_addr            or   RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill           or   RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_4  )
         begin 
             case (1'b1) 
              RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL___near_mem___icache___ram_word64_set$ADDRB  = RTL___near_mem___icache___req_addr [11:3]; 
              RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL___near_mem___icache___ram_word64_set$ADDRB  = RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_2 ; 
              RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq  : 
                  RTL___near_mem___icache___ram_word64_set$ADDRB  = RTL___near_mem___icache___rg_addr [11:3]; 
              RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL___near_mem___icache___ram_word64_set$ADDRB  = RTL___near_mem___icache___MUX_ram_word64_set$b_put_2__VAL_4 ;
              default : 
                  RTL___near_mem___icache___ram_word64_set$ADDRB  =9'b010101010;endcase
         end
  assign  RTL___near_mem___icache___ram_word64_set$DIA = RTL___near_mem___icache___MUX_ram_word64_set$a_put_1__SEL_1  ?  RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:3]: RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 ; 
  always @(     RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1                or   RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2            or   RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq           or   RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  )
         begin 
             case (1'b1) 
              RTL___near_mem___icache___MUX_ram_state_and_ctag_cset$b_put_1__SEL_1  : 
                  RTL___near_mem___icache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___icache___MUX_ram_word64_set$b_put_1__SEL_2  : 
                  RTL___near_mem___icache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq  : 
                  RTL___near_mem___icache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA; 
              RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill  : 
                  RTL___near_mem___icache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;
              default : 
                  RTL___near_mem___icache___ram_word64_set$DIB  =64'hAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL___near_mem___icache___ram_word64_set$WEA =1'd1; 
  assign  RTL___near_mem___icache___ram_word64_set$WEB =1'd0; 
  assign  RTL___near_mem___icache___ram_word64_set$ENA = RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0|| RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 ; 
  assign  RTL___near_mem___icache___ram_word64_set$ENB = RTL___near_mem___icache___EN_req && RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 || RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]!=2'd3|| RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq || RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill ; 
  assign  RTL___near_mem___icache___soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___icache___soc_map$m_is_mem_addr_addr ={32'd0, RTL___near_mem___icache___rg_addr }; 
  assign  RTL___near_mem___icache___soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 = RTL___near_mem___icache___cfg_verbosity >4'd1; 
  assign  RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 = RTL___near_mem___icache___cfg_verbosity >4'd2; 
  assign  RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d114 =(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___icache___NOT_dmem_not_imem_10_OR_soc_map_m_is_mem_addr__ETC___d190 =(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&&! RTL___near_mem___icache___rg_op && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___icache___NOT_req_f3_BITS_1_TO_0_18_EQ_0b0_19_20_AND_NOT_ETC___d539 = RTL___near_mem___icache___req_f3 [1:0]!=2'b0&&( RTL___near_mem___icache___req_f3 [1:0]!=2'b01|| RTL___near_mem___icache___req_addr [0])&&( RTL___near_mem___icache___req_f3 [1:0]!=2'b10|| RTL___near_mem___icache___req_addr [1:0]!=2'b0)&&( RTL___near_mem___icache___req_f3 [1:0]!=2'b11|| RTL___near_mem___icache___req_addr [2:0]!=3'b0); 
  assign  RTL___near_mem___icache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 =! RTL___near_mem___icache___rg_op && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL___near_mem___icache____theResult___snd_fst__h2707 = RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [63:0]<< RTL___near_mem___icache___shift_bits__h2487 ; 
  assign  RTL___near_mem___icache___access_exc_code__h2256 = RTL___near_mem___icache___dmem_not_imem  ? ( RTL___near_mem___icache___rg_op  ? 4'd7:4'd5):4'd1; 
  assign  RTL___near_mem___icache___b__h14485 = RTL___near_mem___icache___CAN_FIRE_RL_rl_fabric_send_write_req  ?  RTL___near_mem___icache___ctr_wr_rsps_pending_crg$port0__write_1 : RTL___near_mem___icache___ctr_wr_rsps_pending_crg ; 
  assign  RTL___near_mem___icache___cline_addr__h14583 ={ RTL___near_mem___icache___rg_pa [31:5],5'd0}; 
  assign  RTL___near_mem___icache___cline_fabric_addr__h14584 ={32'd0, RTL___near_mem___icache___cline_addr__h14583 }; 
  assign  RTL___near_mem___icache___dmem_not_imem_AND_NOT_soc_map_m_is_mem_addr_0__ETC___d106 = RTL___near_mem___icache___dmem_not_imem &&! RTL___near_mem___icache___soc_map$m_is_mem_addr || RTL___near_mem___icache___rg_op ||! RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 ; 
  assign  RTL___near_mem___icache___fabric_addr__h17243 ={32'd0, RTL___near_mem___icache___rg_pa }; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [10:3]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [18:11]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [18:3]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [26:19]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:19]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:27]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:3]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [42:35]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [50:35]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [50:43]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [58:51]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:35]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:51]; 
  assign  RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 = RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:59]; 
  assign  RTL___near_mem___icache___mem_req_wr_addr_awaddr__h2473 ={32'd0, RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [95:64]}; 
  assign  RTL___near_mem___icache___pa_ctag__h4952 ={2'd0, RTL___near_mem___icache___rg_addr [31:12]}; 
  assign  RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 = RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [21:0]== RTL___near_mem___icache___pa_ctag__h4952 ; 
  assign  RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 = RTL___near_mem___icache___req_f3 [1:0]==2'b0|| RTL___near_mem___icache___req_f3 [1:0]==2'b01&&! RTL___near_mem___icache___req_addr [0]|| RTL___near_mem___icache___req_f3 [1:0]==2'b10&& RTL___near_mem___icache___req_addr [1:0]==2'b0|| RTL___near_mem___icache___req_f3 [1:0]==2'b11&& RTL___near_mem___icache___req_addr [2:0]==3'b0; 
  assign  RTL___near_mem___icache___result__h11657 ={{56{ RTL___near_mem___icache___word64094_BITS_15_TO_8__q18 [7]}}, RTL___near_mem___icache___word64094_BITS_15_TO_8__q18 }; 
  assign  RTL___near_mem___icache___result__h11685 ={{56{ RTL___near_mem___icache___word64094_BITS_23_TO_16__q19 [7]}}, RTL___near_mem___icache___word64094_BITS_23_TO_16__q19 }; 
  assign  RTL___near_mem___icache___result__h11713 ={{56{ RTL___near_mem___icache___word64094_BITS_31_TO_24__q21 [7]}}, RTL___near_mem___icache___word64094_BITS_31_TO_24__q21 }; 
  assign  RTL___near_mem___icache___result__h11741 ={{56{ RTL___near_mem___icache___word64094_BITS_39_TO_32__q22 [7]}}, RTL___near_mem___icache___word64094_BITS_39_TO_32__q22 }; 
  assign  RTL___near_mem___icache___result__h11769 ={{56{ RTL___near_mem___icache___word64094_BITS_47_TO_40__q25 [7]}}, RTL___near_mem___icache___word64094_BITS_47_TO_40__q25 }; 
  assign  RTL___near_mem___icache___result__h11797 ={{56{ RTL___near_mem___icache___word64094_BITS_55_TO_48__q26 [7]}}, RTL___near_mem___icache___word64094_BITS_55_TO_48__q26 }; 
  assign  RTL___near_mem___icache___result__h11825 ={{56{ RTL___near_mem___icache___word64094_BITS_63_TO_56__q28 [7]}}, RTL___near_mem___icache___word64094_BITS_63_TO_56__q28 }; 
  assign  RTL___near_mem___icache___result__h11870 ={56'd0, RTL___near_mem___icache___word64__h5094 [7:0]}; 
  assign  RTL___near_mem___icache___result__h11898 ={56'd0, RTL___near_mem___icache___word64__h5094 [15:8]}; 
  assign  RTL___near_mem___icache___result__h11926 ={56'd0, RTL___near_mem___icache___word64__h5094 [23:16]}; 
  assign  RTL___near_mem___icache___result__h11954 ={56'd0, RTL___near_mem___icache___word64__h5094 [31:24]}; 
  assign  RTL___near_mem___icache___result__h11982 ={56'd0, RTL___near_mem___icache___word64__h5094 [39:32]}; 
  assign  RTL___near_mem___icache___result__h12010 ={56'd0, RTL___near_mem___icache___word64__h5094 [47:40]}; 
  assign  RTL___near_mem___icache___result__h12038 ={56'd0, RTL___near_mem___icache___word64__h5094 [55:48]}; 
  assign  RTL___near_mem___icache___result__h12066 ={56'd0, RTL___near_mem___icache___word64__h5094 [63:56]}; 
  assign  RTL___near_mem___icache___result__h12111 ={{48{ RTL___near_mem___icache___word64094_BITS_15_TO_0__q16 [15]}}, RTL___near_mem___icache___word64094_BITS_15_TO_0__q16 }; 
  assign  RTL___near_mem___icache___result__h12139 ={{48{ RTL___near_mem___icache___word64094_BITS_31_TO_16__q20 [15]}}, RTL___near_mem___icache___word64094_BITS_31_TO_16__q20 }; 
  assign  RTL___near_mem___icache___result__h12167 ={{48{ RTL___near_mem___icache___word64094_BITS_47_TO_32__q23 [15]}}, RTL___near_mem___icache___word64094_BITS_47_TO_32__q23 }; 
  assign  RTL___near_mem___icache___result__h12195 ={{48{ RTL___near_mem___icache___word64094_BITS_63_TO_48__q27 [15]}}, RTL___near_mem___icache___word64094_BITS_63_TO_48__q27 }; 
  assign  RTL___near_mem___icache___result__h12236 ={48'd0, RTL___near_mem___icache___word64__h5094 [15:0]}; 
  assign  RTL___near_mem___icache___result__h12264 ={48'd0, RTL___near_mem___icache___word64__h5094 [31:16]}; 
  assign  RTL___near_mem___icache___result__h12292 ={48'd0, RTL___near_mem___icache___word64__h5094 [47:32]}; 
  assign  RTL___near_mem___icache___result__h12320 ={48'd0, RTL___near_mem___icache___word64__h5094 [63:48]}; 
  assign  RTL___near_mem___icache___result__h12361 ={{32{ RTL___near_mem___icache___word64094_BITS_31_TO_0__q17 [31]}}, RTL___near_mem___icache___word64094_BITS_31_TO_0__q17 }; 
  assign  RTL___near_mem___icache___result__h12389 ={{32{ RTL___near_mem___icache___word64094_BITS_63_TO_32__q24 [31]}}, RTL___near_mem___icache___word64094_BITS_63_TO_32__q24 }; 
  assign  RTL___near_mem___icache___result__h12428 ={32'd0, RTL___near_mem___icache___word64__h5094 [31:0]}; 
  assign  RTL___near_mem___icache___result__h12456 ={32'd0, RTL___near_mem___icache___word64__h5094 [63:32]}; 
  assign  RTL___near_mem___icache___result__h17654 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_10_TO_3__q1 }; 
  assign  RTL___near_mem___icache___result__h17684 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_11__q4 }; 
  assign  RTL___near_mem___icache___result__h17711 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_26_TO_19__q5 }; 
  assign  RTL___near_mem___icache___result__h17738 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_27__q7 }; 
  assign  RTL___near_mem___icache___result__h17765 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_42_TO_35__q8 }; 
  assign  RTL___near_mem___icache___result__h17792 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_43__q11 }; 
  assign  RTL___near_mem___icache___result__h17819 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_58_TO_51__q12 }; 
  assign  RTL___near_mem___icache___result__h17846 ={{56{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 [7]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_59__q14 }; 
  assign  RTL___near_mem___icache___result__h17890 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [10:3]}; 
  assign  RTL___near_mem___icache___result__h17917 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [18:11]}; 
  assign  RTL___near_mem___icache___result__h17944 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [26:19]}; 
  assign  RTL___near_mem___icache___result__h17971 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:27]}; 
  assign  RTL___near_mem___icache___result__h17998 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [42:35]}; 
  assign  RTL___near_mem___icache___result__h18025 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [50:43]}; 
  assign  RTL___near_mem___icache___result__h18052 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [58:51]}; 
  assign  RTL___near_mem___icache___result__h18079 ={56'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:59]}; 
  assign  RTL___near_mem___icache___result__h18123 ={{48{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 [15]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_18_TO_3__q2 }; 
  assign  RTL___near_mem___icache___result__h18150 ={{48{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 [15]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_19__q6 }; 
  assign  RTL___near_mem___icache___result__h18177 ={{48{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 [15]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_50_TO_35__q9 }; 
  assign  RTL___near_mem___icache___result__h18204 ={{48{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 [15]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_51__q13 }; 
  assign  RTL___near_mem___icache___result__h18244 ={48'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [18:3]}; 
  assign  RTL___near_mem___icache___result__h18271 ={48'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:19]}; 
  assign  RTL___near_mem___icache___result__h18298 ={48'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [50:35]}; 
  assign  RTL___near_mem___icache___result__h18325 ={48'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:51]}; 
  assign  RTL___near_mem___icache___result__h18365 ={{32{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 [31]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_34_TO_3__q3 }; 
  assign  RTL___near_mem___icache___result__h18392 ={{32{ RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 [31]}}, RTL___near_mem___icache___master_xactor_f_rd_dataD_OUT_BITS_66_TO_35__q10 }; 
  assign  RTL___near_mem___icache___result__h18430 ={32'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [34:3]}; 
  assign  RTL___near_mem___icache___result__h18457 ={32'd0, RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:35]}; 
  assign  RTL___near_mem___icache___result__h5301 ={{56{ RTL___near_mem___icache___word64094_BITS_7_TO_0__q15 [7]}}, RTL___near_mem___icache___word64094_BITS_7_TO_0__q15 }; 
  assign  RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 = RTL___near_mem___icache___rg_op && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 ; 
  assign  RTL___near_mem___icache___shift_bits__h2487 ={ RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [66:64],3'b0}; 
  assign  RTL___near_mem___icache___strobe64__h2637 =8'b00000001<< RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___icache___strobe64__h2639 =8'b00000011<< RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___icache___strobe64__h2641 =8'b00001111<< RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [66:64]; 
  assign  RTL___near_mem___icache___word64094_BITS_15_TO_0__q16 = RTL___near_mem___icache___word64__h5094 [15:0]; 
  assign  RTL___near_mem___icache___word64094_BITS_15_TO_8__q18 = RTL___near_mem___icache___word64__h5094 [15:8]; 
  assign  RTL___near_mem___icache___word64094_BITS_23_TO_16__q19 = RTL___near_mem___icache___word64__h5094 [23:16]; 
  assign  RTL___near_mem___icache___word64094_BITS_31_TO_0__q17 = RTL___near_mem___icache___word64__h5094 [31:0]; 
  assign  RTL___near_mem___icache___word64094_BITS_31_TO_16__q20 = RTL___near_mem___icache___word64__h5094 [31:16]; 
  assign  RTL___near_mem___icache___word64094_BITS_31_TO_24__q21 = RTL___near_mem___icache___word64__h5094 [31:24]; 
  assign  RTL___near_mem___icache___word64094_BITS_39_TO_32__q22 = RTL___near_mem___icache___word64__h5094 [39:32]; 
  assign  RTL___near_mem___icache___word64094_BITS_47_TO_32__q23 = RTL___near_mem___icache___word64__h5094 [47:32]; 
  assign  RTL___near_mem___icache___word64094_BITS_47_TO_40__q25 = RTL___near_mem___icache___word64__h5094 [47:40]; 
  assign  RTL___near_mem___icache___word64094_BITS_55_TO_48__q26 = RTL___near_mem___icache___word64__h5094 [55:48]; 
  assign  RTL___near_mem___icache___word64094_BITS_63_TO_32__q24 = RTL___near_mem___icache___word64__h5094 [63:32]; 
  assign  RTL___near_mem___icache___word64094_BITS_63_TO_48__q27 = RTL___near_mem___icache___word64__h5094 [63:48]; 
  assign  RTL___near_mem___icache___word64094_BITS_63_TO_56__q28 = RTL___near_mem___icache___word64__h5094 [63:56]; 
  assign  RTL___near_mem___icache___word64094_BITS_7_TO_0__q15 = RTL___near_mem___icache___word64__h5094 [7:0]; 
  assign  RTL___near_mem___icache___word64__h5094 = RTL___near_mem___icache___ram_word64_set$DOB & RTL___near_mem___icache___y__h5337 ; 
  assign  RTL___near_mem___icache___y__h5337 ={64{ RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]&& RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 }}; 
  always @(  RTL___near_mem___icache___f_fabric_write_reqs$D_OUT  )
         begin 
             case ( RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL___near_mem___icache___x__h2520  =3'b0;
              2 'b01: 
                  RTL___near_mem___icache___x__h2520  =3'b001;
              2 'b10: 
                  RTL___near_mem___icache___x__h2520  =3'b010;
              2 'b11: 
                  RTL___near_mem___icache___x__h2520  =3'b011;endcase
         end
  always @(  RTL___near_mem___icache___rg_f3  )
         begin 
             case ( RTL___near_mem___icache___rg_f3 [1:0])
              2 'b0: 
                  RTL___near_mem___icache___value__h17372  =3'b0;
              2 'b01: 
                  RTL___near_mem___icache___value__h17372  =3'b001;
              2 'b10: 
                  RTL___near_mem___icache___value__h17372  =3'b010;
              2 'd3: 
                  RTL___near_mem___icache___value__h17372  =3'b011;endcase
         end
  always @(     RTL___near_mem___icache___f_fabric_write_reqs$D_OUT                or   RTL___near_mem___icache___strobe64__h2637            or   RTL___near_mem___icache___strobe64__h2639           or   RTL___near_mem___icache___strobe64__h2641  )
         begin 
             case ( RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0: 
                  RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___icache___strobe64__h2637 ;
              2 'b01: 
                  RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___icache___strobe64__h2639 ;
              2 'b10: 
                  RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700  = RTL___near_mem___icache___strobe64__h2641 ;
              2 'b11: 
                  RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700  =8'b11111111;endcase
         end
  always @(   RTL___near_mem___icache___f_fabric_write_reqs$D_OUT            or   RTL___near_mem___icache____theResult___snd_fst__h2707  )
         begin 
             case ( RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [97:96])
              2 'b0,2'b01,2'b10: 
                  RTL___near_mem___icache___mem_req_wr_data_wdata__h2699  = RTL___near_mem___icache____theResult___snd_fst__h2707 ;
              2 'd3: 
                  RTL___near_mem___icache___mem_req_wr_data_wdata__h2699  = RTL___near_mem___icache___f_fabric_write_reqs$D_OUT [63:0];endcase
         end
  always @(      RTL___near_mem___icache___rg_addr                  or   RTL___near_mem___icache___result__h12111             or   RTL___near_mem___icache___result__h12139            or   RTL___near_mem___icache___result__h12167           or   RTL___near_mem___icache___result__h12195  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___icache___result__h12111 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___icache___result__h12139 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___icache___result__h12167 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  = RTL___near_mem___icache___result__h12195 ;
              default : 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d276  =64'd0;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___ram_word64_set$DOB           or   RTL___near_mem___icache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:16], RTL___near_mem___icache___rg_st_amo_val [15:0]};
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:32], RTL___near_mem___icache___rg_st_amo_val [15:0], RTL___near_mem___icache___ram_word64_set$DOB [15:0]};
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:48], RTL___near_mem___icache___rg_st_amo_val [15:0], RTL___near_mem___icache___ram_word64_set$DOB [31:0]};
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  ={ RTL___near_mem___icache___rg_st_amo_val [15:0], RTL___near_mem___icache___ram_word64_set$DOB [47:0]};
              default : 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167  = RTL___near_mem___icache___ram_word64_set$DOB ;endcase
         end
  always @(          RTL___near_mem___icache___rg_addr                          or   RTL___near_mem___icache___result__h5301                 or   RTL___near_mem___icache___result__h11657                or   RTL___near_mem___icache___result__h11685               or   RTL___near_mem___icache___result__h11713              or   RTL___near_mem___icache___result__h11741             or   RTL___near_mem___icache___result__h11769            or   RTL___near_mem___icache___result__h11797           or   RTL___near_mem___icache___result__h11825  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h5301 ;
              3 'h1: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11657 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11685 ;
              3 'h3: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11713 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11741 ;
              3 'h5: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11769 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11797 ;
              3 'h7: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d247  = RTL___near_mem___icache___result__h11825 ;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___ram_word64_set$DOB           or   RTL___near_mem___icache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:8], RTL___near_mem___icache___rg_st_amo_val [7:0]};
              3 'h1: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:16], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [7:0]};
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:24], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [15:0]};
              3 'h3: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:32], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [23:0]};
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:40], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [31:0]};
              3 'h5: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:48], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [39:0]};
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:56], RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [47:0]};
              3 'h7: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157  ={ RTL___near_mem___icache___rg_st_amo_val [7:0], RTL___near_mem___icache___ram_word64_set$DOB [55:0]};endcase
         end
  always @(      RTL___near_mem___icache___rg_addr                  or   RTL___near_mem___icache___result__h18244             or   RTL___near_mem___icache___result__h18271            or   RTL___near_mem___icache___result__h18298           or   RTL___near_mem___icache___result__h18325  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___icache___result__h18244 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___icache___result__h18271 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___icache___result__h18298 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  = RTL___near_mem___icache___result__h18325 ;
              default : 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447  =64'd0;endcase
         end
  always @(      RTL___near_mem___icache___rg_addr                  or   RTL___near_mem___icache___result__h12236             or   RTL___near_mem___icache___result__h12264            or   RTL___near_mem___icache___result__h12292           or   RTL___near_mem___icache___result__h12320  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___icache___result__h12236 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___icache___result__h12264 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___icache___result__h12292 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  = RTL___near_mem___icache___result__h12320 ;
              default : 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d285  =64'd0;endcase
         end
  always @(      RTL___near_mem___icache___rg_addr                  or   RTL___near_mem___icache___result__h18123             or   RTL___near_mem___icache___result__h18150            or   RTL___near_mem___icache___result__h18177           or   RTL___near_mem___icache___result__h18204  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___icache___result__h18123 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___icache___result__h18150 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___icache___result__h18177 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  = RTL___near_mem___icache___result__h18204 ;
              default : 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439  =64'd0;endcase
         end
  always @(          RTL___near_mem___icache___rg_addr                          or   RTL___near_mem___icache___result__h17890                 or   RTL___near_mem___icache___result__h17917                or   RTL___near_mem___icache___result__h17944               or   RTL___near_mem___icache___result__h17971              or   RTL___near_mem___icache___result__h17998             or   RTL___near_mem___icache___result__h18025            or   RTL___near_mem___icache___result__h18052           or   RTL___near_mem___icache___result__h18079  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h17890 ;
              3 'h1: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h17917 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h17944 ;
              3 'h3: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h17971 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h17998 ;
              3 'h5: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h18025 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h18052 ;
              3 'h7: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427  = RTL___near_mem___icache___result__h18079 ;endcase
         end
  always @(          RTL___near_mem___icache___rg_addr                          or   RTL___near_mem___icache___result__h11870                 or   RTL___near_mem___icache___result__h11898                or   RTL___near_mem___icache___result__h11926               or   RTL___near_mem___icache___result__h11954              or   RTL___near_mem___icache___result__h11982             or   RTL___near_mem___icache___result__h12010            or   RTL___near_mem___icache___result__h12038           or   RTL___near_mem___icache___result__h12066  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h11870 ;
              3 'h1: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h11898 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h11926 ;
              3 'h3: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h11954 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h11982 ;
              3 'h5: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h12010 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h12038 ;
              3 'h7: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d264  = RTL___near_mem___icache___result__h12066 ;endcase
         end
  always @(          RTL___near_mem___icache___rg_addr                          or   RTL___near_mem___icache___result__h17654                 or   RTL___near_mem___icache___result__h17684                or   RTL___near_mem___icache___result__h17711               or   RTL___near_mem___icache___result__h17738              or   RTL___near_mem___icache___result__h17765             or   RTL___near_mem___icache___result__h17792            or   RTL___near_mem___icache___result__h17819           or   RTL___near_mem___icache___result__h17846  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17654 ;
              3 'h1: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17684 ;
              3 'h2: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17711 ;
              3 'h3: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17738 ;
              3 'h4: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17765 ;
              3 'h5: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17792 ;
              3 'h6: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17819 ;
              3 'h7: 
                  RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411  = RTL___near_mem___icache___result__h17846 ;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___result__h18365           or   RTL___near_mem___icache___result__h18392  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL___near_mem___icache___result__h18365 ;
              3 'h4: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  = RTL___near_mem___icache___result__h18392 ;
              default : 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29  =64'd0;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___result__h18430           or   RTL___near_mem___icache___result__h18457  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL___near_mem___icache___result__h18430 ;
              3 'h4: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  = RTL___near_mem___icache___result__h18457 ;
              default : 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  =64'd0;endcase
         end
  always @(          RTL___near_mem___icache___rg_f3                          or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411                 or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439                or   RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29               or   RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT             or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427            or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447           or   RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30  )
         begin 
             case ( RTL___near_mem___icache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d411 ;
              3 'b001: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_SEXT_ETC___d439 ;
              3 'b010: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8365_0x4_re_ETC__q29 ;
              3 'b011: 
                  RTL___near_mem___icache___ld_val__h17594  =( RTL___near_mem___icache___rg_addr [2:0]==3'h0) ?  RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:3]:64'd0;
              3 'b100: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d427 ;
              3 'b101: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_0_CO_ETC___d447 ;
              3 'b110: 
                  RTL___near_mem___icache___ld_val__h17594  = RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result8430_0x4_re_ETC__q30 ;
              3 'd7: 
                  RTL___near_mem___icache___ld_val__h17594  =64'd0;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___ram_word64_set$DOB           or   RTL___near_mem___icache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL___near_mem___icache___ram_word64_set$DOB [63:32], RTL___near_mem___icache___rg_st_amo_val [31:0]};
              3 'h4: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  ={ RTL___near_mem___icache___rg_st_amo_val [31:0], RTL___near_mem___icache___ram_word64_set$DOB [31:0]};
              default : 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31  = RTL___near_mem___icache___ram_word64_set$DOB ;endcase
         end
  always @(       RTL___near_mem___icache___rg_f3                    or   RTL___near_mem___icache___ram_word64_set$DOB              or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157             or   RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167            or   RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31           or   RTL___near_mem___icache___rg_st_amo_val  )
         begin 
             case ( RTL___near_mem___icache___rg_f3 )
              3 'b0: 
                  RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d157 ;
              3 'b001: 
                  RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___icache___IF_rg_addr_6_BITS_2_TO_0_4_EQ_0x0_18_THEN_ram__ETC___d167 ;
              3 'b010: 
                  RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_ram_word64_setDO_ETC__q31 ;
              3 'b011: 
                  RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___icache___rg_st_amo_val ;
              default : 
                  RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178  = RTL___near_mem___icache___ram_word64_set$DOB ;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___result__h12361           or   RTL___near_mem___icache___result__h12389  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL___near_mem___icache___result__h12361 ;
              3 'h4: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  = RTL___near_mem___icache___result__h12389 ;
              default : 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2361_0x4_re_ETC__q32  =64'd0;endcase
         end
  always @(    RTL___near_mem___icache___rg_addr              or   RTL___near_mem___icache___result__h12428           or   RTL___near_mem___icache___result__h12456  )
         begin 
             case ( RTL___near_mem___icache___rg_addr [2:0])
              3 'h0: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL___near_mem___icache___result__h12428 ;
              3 'h4: 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  = RTL___near_mem___icache___result__h12456 ;
              default : 
                  RTL___near_mem___icache___CASE_rg_addr_BITS_2_TO_0_0x0_result2428_0x4_re_ETC__q33  =64'd0;endcase
         end
  always @( posedge  RTL___near_mem___icache___CLK )
         begin 
             if ( RTL___near_mem___icache___RST_N ==1'b0)
                 begin  
                     RTL___near_mem___icache___cfg_verbosity  <=4'd0; 
                     RTL___near_mem___icache___ctr_wr_rsps_pending_crg  <=4'd0; 
                     RTL___near_mem___icache___rg_cset_in_cache  <=7'd0; 
                     RTL___near_mem___icache___rg_lower_word32_full  <=1'd0; 
                     RTL___near_mem___icache___rg_state  <=4'd0;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___icache___cfg_verbosity$EN ) 
                         RTL___near_mem___icache___cfg_verbosity  <= RTL___near_mem___icache___cfg_verbosity$D_IN ;
                     if ( RTL___near_mem___icache___ctr_wr_rsps_pending_crg$EN ) 
                         RTL___near_mem___icache___ctr_wr_rsps_pending_crg  <= RTL___near_mem___icache___ctr_wr_rsps_pending_crg$D_IN ;
                     if ( RTL___near_mem___icache___rg_cset_in_cache$EN ) 
                         RTL___near_mem___icache___rg_cset_in_cache  <= RTL___near_mem___icache___rg_cset_in_cache$D_IN ;
                     if ( RTL___near_mem___icache___rg_lower_word32_full$EN ) 
                         RTL___near_mem___icache___rg_lower_word32_full  <= RTL___near_mem___icache___rg_lower_word32_full$D_IN ;
                     if ( RTL___near_mem___icache___rg_state$EN ) 
                         RTL___near_mem___icache___rg_state  <= RTL___near_mem___icache___rg_state$D_IN ;
                 end 
             if ( RTL___near_mem___icache___rg_addr$EN ) 
                 RTL___near_mem___icache___rg_addr  <= RTL___near_mem___icache___rg_addr$D_IN ;
             if ( RTL___near_mem___icache___rg_error_during_refill$EN ) 
                 RTL___near_mem___icache___rg_error_during_refill  <= RTL___near_mem___icache___rg_error_during_refill$D_IN ;
             if ( RTL___near_mem___icache___rg_exc_code$EN ) 
                 RTL___near_mem___icache___rg_exc_code  <= RTL___near_mem___icache___rg_exc_code$D_IN ;
             if ( RTL___near_mem___icache___rg_f3$EN ) 
                 RTL___near_mem___icache___rg_f3  <= RTL___near_mem___icache___rg_f3$D_IN ;
             if ( RTL___near_mem___icache___rg_ld_val$EN ) 
                 RTL___near_mem___icache___rg_ld_val  <= RTL___near_mem___icache___rg_ld_val$D_IN ;
             if ( RTL___near_mem___icache___rg_lower_word32$EN ) 
                 RTL___near_mem___icache___rg_lower_word32  <= RTL___near_mem___icache___rg_lower_word32$D_IN ;
             if ( RTL___near_mem___icache___rg_op$EN ) 
                 RTL___near_mem___icache___rg_op  <= RTL___near_mem___icache___rg_op$D_IN ;
             if ( RTL___near_mem___icache___rg_pa$EN ) 
                 RTL___near_mem___icache___rg_pa  <= RTL___near_mem___icache___rg_pa$D_IN ;
             if ( RTL___near_mem___icache___rg_pte_pa$EN ) 
                 RTL___near_mem___icache___rg_pte_pa  <= RTL___near_mem___icache___rg_pte_pa$D_IN ;
             if ( RTL___near_mem___icache___rg_st_amo_val$EN ) 
                 RTL___near_mem___icache___rg_st_amo_val  <= RTL___near_mem___icache___rg_st_amo_val$D_IN ;
             if ( RTL___near_mem___icache___rg_word64_set_in_cache$EN ) 
                 RTL___near_mem___icache___rg_word64_set_in_cache  <= RTL___near_mem___icache___rg_word64_set_in_cache$D_IN ;
         end
  always @( negedge  RTL___near_mem___icache___CLK )
         begin #0;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___ctr_wr_rsps_pending_crg ==4'd15)
                     begin  
                         RTL___near_mem___icache___v__h2948  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h2942  = RTL___near_mem___icache___v__h2948 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___ctr_wr_rsps_pending_crg ==4'd15)$display("%0d: ERROR: CreditCounter: overflow", RTL___near_mem___icache___v__h2942 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___ctr_wr_rsps_pending_crg ==4'd15)$finish(32'd1);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Addr { ","awid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awaddr: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___mem_req_wr_addr_awaddr__h2473 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlen: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awsize: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___x__h2520 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awburst: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awlock: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awcache: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awprot: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awqos: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awregion: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","awuser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("                       ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Data { ","wdata: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___mem_req_wr_data_wdata__h2699 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wstrb: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___mem_req_wr_data_wstrb__h2700 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wlast: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("True");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","wuser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_fabric_send_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127&& RTL___near_mem___icache___cfg_verbosity !=4'd0&&! RTL___near_mem___icache___f_reset_reqs$D_OUT )
                     begin  
                         RTL___near_mem___icache___v__h3848  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h3842  = RTL___near_mem___icache___v__h3848 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127&& RTL___near_mem___icache___cfg_verbosity !=4'd0&&! RTL___near_mem___icache___f_reset_reqs$D_OUT )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL___near_mem___icache___v__h3842 ,"D_MMU_Cache",$signed(32'd128),$signed(32'd1));
                      else $display("%0d: %s.rl_reset: %0d sets x %0d ways: all tag states reset to CTAG_EMPTY", RTL___near_mem___icache___v__h3842 ,"I_MMU_Cache",$signed(32'd128),$signed(32'd1));
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___f_reset_reqs$D_OUT )
                     begin  
                         RTL___near_mem___icache___v__h3949  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h3943  = RTL___near_mem___icache___v__h3949 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_reset && RTL___near_mem___icache___rg_cset_in_cache ==7'd127&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___f_reset_reqs$D_OUT )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_reset: Flushed", RTL___near_mem___icache___v__h3943 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_reset: Flushed", RTL___near_mem___icache___v__h3943 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h4098  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h4092  = RTL___near_mem___icache___v__h4098 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL___near_mem___icache___v__h4092 ,"D_MMU_Cache", RTL___near_mem___icache___rg_addr );
                      else $display("%0d: %s: rl_probe_and_immed_rsp; eaddr %0h", RTL___near_mem___icache___v__h4092 ,"I_MMU_Cache", RTL___near_mem___icache___rg_addr );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        eaddr = {CTag 0x%0h  CSet 0x%0h  Word64 0x%0h  Byte 0x%0h}", RTL___near_mem___icache___pa_ctag__h4952 , RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_addr [4:3], RTL___near_mem___icache___rg_addr [2:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x: (state, tag):", RTL___near_mem___icache___rg_addr [11:5]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" (");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22])$write("CTAG_CLEAN");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22])$write("CTAG_EMPTY");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22])$write(", 0x%0x", RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [21:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22])$write(", --");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(")");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_addr [4:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" 0x%0x", RTL___near_mem___icache___ram_word64_set$DOB );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    TLB result: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_Xlate_Result { ","outcome: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("VM_XLATE_OK");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","pa: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___rg_addr );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","exc_code: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'hA," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp && RTL___near_mem___icache___dmem_not_imem &&! RTL___near_mem___icache___soc_map$m_is_mem_addr && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => IO_REQ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$display("        Write-Cache-Hit: pa 0x%0h word64 0x%0h", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_st_amo_val );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        New Word64_Set:");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_addr [4:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write(" 0x%0x", RTL___near_mem___icache___IF_rg_f3_16_EQ_0b0_17_THEN_IF_rg_addr_6_BITS_2_ETC___d178 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op_1_AND_ram_state_and_ctag_cset_b_read__5__ETC___d180 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op &&(! RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Miss: pa 0x%0h word64 0x%0h", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_st_amo_val );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Write-Cache-Hit/Miss: eaddr 0x%0h word64 0x%0h", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_st_amo_val );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___rg_op && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        => rl_write_response");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     begin  
                         RTL___near_mem___icache___v__h12540  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h12534  = RTL___near_mem___icache___v__h12540 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL___near_mem___icache___v__h12534 ,"D_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___word64__h5094 ,64'd0);
                      else $display("%0d: %s.drive_mem_rsp: addr 0x%0h ld_val 0x%0h st_amo_val 0x%0h", RTL___near_mem___icache___v__h12534 ,"I_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___word64__h5094 ,64'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&& RTL___near_mem___icache___NOT_rg_op_1_2_AND_ram_state_and_ctag_cset_b_re_ETC___d305 )$display("        Read-hit: addr 0x%0h word64 0x%0h", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___word64__h5094 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_probe_and_immed_rsp &&(! RTL___near_mem___icache___dmem_not_imem || RTL___near_mem___icache___soc_map$m_is_mem_addr )&&! RTL___near_mem___icache___rg_op &&(! RTL___near_mem___icache___ram_state_and_ctag_cset$DOB [22]||! RTL___near_mem___icache___ram_state_and_ctag_cset_b_read__5_BITS_21_TO_0_ETC___d102 )&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("        Read Miss: -> CACHE_START_REFILL.");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h14531  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h14525  = RTL___near_mem___icache___v__h14531 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_start_cache_refill: ", RTL___near_mem___icache___v__h14525 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_cache_refill: ", RTL___near_mem___icache___v__h14525 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    To fabric: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___cline_fabric_addr__h14584 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd3);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'b011);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_cache_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    Victim way %0d; => CACHE_REFILL",1'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     begin  
                         RTL___near_mem___icache___v__h15336  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h15330  = RTL___near_mem___icache___v__h15336 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop:", RTL___near_mem___icache___v__h15330 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_cache_refill_rsps_loop:", RTL___near_mem___icache___v__h15330 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rdata: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rresp: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","rlast: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 &&! RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(", ","ruser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h15578  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h15572  = RTL___near_mem___icache___v__h15578 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL___near_mem___icache___v__h15572 ,"D_MMU_Cache", RTL___near_mem___icache___access_exc_code__h2256 );
                      else $display("%0d: %s.rl_cache_refill_rsps_loop: FABRIC_RSP_ERR: raising access exception %0d", RTL___near_mem___icache___v__h15572 ,"I_MMU_Cache", RTL___near_mem___icache___access_exc_code__h2256 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]==2'd3&&( RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0|| RTL___near_mem___icache___rg_error_during_refill )&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => MODULE_EXCEPTION_RSP");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___rg_word64_set_in_cache [1:0]==2'd3&& RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&&! RTL___near_mem___icache___rg_error_during_refill && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => CACHE_REREQ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$display("        Updating Cache word64_set 0x%0h, word64_in_cline %0d) old => new", RTL___near_mem___icache___rg_word64_set_in_cache , RTL___near_mem___icache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL___near_mem___icache___ram_word64_set$DOB );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("        CSet 0x%0x, Word64 0x%0x: ", RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_word64_set_in_cache [1:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write(" 0x%0x", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_cache_refill_rsps_loop && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_2_30___d331 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_rereq && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL___near_mem___icache___rg_addr [11:5], RTL___near_mem___icache___rg_addr [11:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h17191  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h17185  = RTL___near_mem___icache___v__h17191 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL___near_mem___icache___v__h17185 ,"D_MMU_Cache", RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa );
                      else $display("%0d: %s.rl_io_read_req; f3 0x%0h vaddr %0h  paddr %0h", RTL___near_mem___icache___v__h17185 ,"I_MMU_Cache", RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("            To fabric: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Addr { ","arid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","araddr: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___fabric_addr__h17243 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlen: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",8'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arsize: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___value__h17372 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arburst: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",2'b01);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arlock: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arcache: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'b0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arprot: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",3'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arqos: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","arregion: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",4'd0);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","aruser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'h0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h17485  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h17479  = RTL___near_mem___icache___v__h17485 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL___near_mem___icache___v__h17479 ,"D_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa );
                      else $display("%0d: %s.rl_io_read_rsp: vaddr 0x%0h  paddr 0x%0h", RTL___near_mem___icache___v__h17479 ,"I_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Rd_Data { ","rid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [70:67]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rdata: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [66:3]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rresp: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","rlast: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [0])$write("True");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [0])$write("False");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","ruser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h18585  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h18579  = RTL___near_mem___icache___v__h18585 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___icache___v__h18579 ,"D_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___ld_val__h17594 );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___icache___v__h18579 ,"I_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___ld_val__h17594 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h18692  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h18686  = RTL___near_mem___icache___v__h18692 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_read_rsp && RTL___near_mem___icache___master_xactor_f_rd_data$D_OUT [2:1]!=2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL___near_mem___icache___v__h18686 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_io_read_rsp: FABRIC_RSP_ERR: raising trap LOAD_ACCESS_FAULT", RTL___near_mem___icache___v__h18686 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h18797  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h18791  = RTL___near_mem___icache___v__h18797 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_maintain_io_read_rsp && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___icache___v__h18791 ,"D_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_ld_val );
                      else $display("%0d: %s.drive_IO_read_rsp: addr 0x%0h ld_val 0x%0h", RTL___near_mem___icache___v__h18791 ,"I_MMU_Cache", RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_ld_val );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h18877  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h18871  = RTL___near_mem___icache___v__h18877 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL___near_mem___icache___v__h18871 ,"D_MMU_Cache", RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa , RTL___near_mem___icache___rg_st_amo_val );
                      else $display("%0d: %s: rl_io_write_req; f3 0x%0h  vaddr %0h  paddr %0h  word64 0x%0h", RTL___near_mem___icache___v__h18871 ,"I_MMU_Cache", RTL___near_mem___icache___rg_f3 , RTL___near_mem___icache___rg_addr , RTL___near_mem___icache___rg_pa , RTL___near_mem___icache___rg_st_amo_val );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_io_write_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    => rl_ST_AMO_response");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h19505  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h19499  = RTL___near_mem___icache___v__h19505 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL___near_mem___icache___v__h19499 ,"D_MMU_Cache",$unsigned( RTL___near_mem___icache___b__h14485 ));
                      else $write("%0d: %s.rl_discard_write_rsp: pending %0d ", RTL___near_mem___icache___v__h19499 ,"I_MMU_Cache",$unsigned( RTL___near_mem___icache___b__h14485 ));
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","bresp: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h", RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(", ","buser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("'h%h",1'd0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]==2'b0&& RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     begin  
                         RTL___near_mem___icache___v__h19466  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h19460  = RTL___near_mem___icache___v__h19466 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL___near_mem___icache___v__h19460 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_discard_write_rsp: fabric response error: exit", RTL___near_mem___icache___v__h19460 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("    ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("AXI4_Wr_Resp { ","bid: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [5:2]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","bresp: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h", RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]);
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write(", ","buser: ");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("'h%h",1'd0," }");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_discard_write_rsp && RTL___near_mem___icache___master_xactor_f_wr_resp$D_OUT [1:0]!=2'b0)$write("\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h3483  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h3477  = RTL___near_mem___icache___v__h3483 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___WILL_FIRE_RL_rl_start_reset && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     if ( RTL___near_mem___icache___dmem_not_imem )$display("%0d: %s.rl_start_reset", RTL___near_mem___icache___v__h3477 ,"D_MMU_Cache");
                      else $display("%0d: %s.rl_start_reset", RTL___near_mem___icache___v__h3477 ,"I_MMU_Cache");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )
                     begin  
                         RTL___near_mem___icache___v__h19852  =$stime;#0;
                     end  
             RTL___near_mem___icache___v__h19846  = RTL___near_mem___icache___v__h19852 /32'd10;
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("%0d: %m.req: op:", RTL___near_mem___icache___v__h19846 );
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___req_op )$write("CACHE_ST");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 &&! RTL___near_mem___icache___req_op )$write("CACHE_LD");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" f3:%0d addr:0x%0h st_value:0x%0h", RTL___near_mem___icache___req_f3 , RTL___near_mem___icache___req_addr , RTL___near_mem___icache___req_st_value ,"\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write("    priv:");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___req_priv ==2'b0)$write("U");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___req_priv ==2'b01)$write("S");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___req_priv ==2'b11)$write("M");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 && RTL___near_mem___icache___req_priv !=2'b0&& RTL___near_mem___icache___req_priv !=2'b01&& RTL___near_mem___icache___req_priv !=2'b11)$write("RESERVED");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$write(" sstatus_SUM:%0d mstatus_MXR:%0d satp:0x%0h", RTL___near_mem___icache___req_sstatus_SUM , RTL___near_mem___icache___req_mstatus_MXR , RTL___near_mem___icache___req_satp ,"\n");
             if ( RTL___near_mem___icache___RST_N !=1'b0)
                 if ( RTL___near_mem___icache___EN_req && RTL___near_mem___icache___req_f3_BITS_1_TO_0_18_EQ_0b0_19_OR_req_f3_BITS_ETC___d548 && RTL___near_mem___icache___NOT_cfg_verbosity_read__0_ULE_1_1___d42 )$display("    fa_req_ram_B tagCSet [0x%0x] word64_set [0x%0d]", RTL___near_mem___icache___req_addr [11:5], RTL___near_mem___icache___req_addr [11:3]);
         end
  assign  RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL___near_mem___icache___rg_addr ; 
  assign  RTL___near_mem___icache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL___near_mem___icache___rg_pa ;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL___near_mem___dcache___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL___near_mem___dcache___CLK = RTL___near_mem___CLK;
    assign RTL___near_mem___dcache___RST_N = RTL___near_mem___RST_N;
    assign RTL___near_mem___dcache___set_verbosity_verbosity = RTL___near_mem___dcache$set_verbosity_verbosity;
    assign RTL___near_mem___dcache___EN_set_verbosity = RTL___near_mem___dcache$EN_set_verbosity;
    assign RTL___near_mem___dcache___EN_server_reset_request_put = RTL___near_mem___dcache$EN_server_reset_request_put;
    assign RTL___near_mem___dcache$RDY_server_reset_request_put = RTL___near_mem___dcache___RDY_server_reset_request_put;
    assign RTL___near_mem___dcache___EN_server_reset_response_get = RTL___near_mem___dcache$EN_server_reset_response_get;
    assign RTL___near_mem___dcache$RDY_server_reset_response_get = RTL___near_mem___dcache___RDY_server_reset_response_get;
    assign RTL___near_mem___dcache___req_op = RTL___near_mem___dcache$req_op;
    assign RTL___near_mem___dcache___req_f3 = RTL___near_mem___dcache$req_f3;
    assign RTL___near_mem___dcache___req_addr = RTL___near_mem___dcache$req_addr;
    assign RTL___near_mem___dcache___req_st_value = RTL___near_mem___dcache$req_st_value;
    assign RTL___near_mem___dcache___req_priv = RTL___near_mem___dcache$req_priv;
    assign RTL___near_mem___dcache___req_sstatus_SUM = RTL___near_mem___dcache$req_sstatus_SUM;
    assign RTL___near_mem___dcache___req_mstatus_MXR = RTL___near_mem___dcache$req_mstatus_MXR;
    assign RTL___near_mem___dcache___req_satp = RTL___near_mem___dcache$req_satp;
    assign RTL___near_mem___dcache___EN_req = RTL___near_mem___dcache$EN_req;
    assign RTL___near_mem___dcache$valid = RTL___near_mem___dcache___valid;
    assign RTL___near_mem___dcache$word64 = RTL___near_mem___dcache___word64;
    assign RTL___near_mem___dcache$exc = RTL___near_mem___dcache___exc;
    assign RTL___near_mem___dcache$exc_code = RTL___near_mem___dcache___exc_code;
    assign RTL___near_mem___dcache___EN_server_flush_request_put = RTL___near_mem___dcache$EN_server_flush_request_put;
    assign RTL___near_mem___dcache$RDY_server_flush_request_put = RTL___near_mem___dcache___RDY_server_flush_request_put;
    assign RTL___near_mem___dcache___EN_server_flush_response_get = RTL___near_mem___dcache$EN_server_flush_response_get;
    assign RTL___near_mem___dcache$RDY_server_flush_response_get = RTL___near_mem___dcache___RDY_server_flush_response_get;
    assign RTL___near_mem___dcache___EN_tlb_flush = RTL___near_mem___dcache$EN_tlb_flush;
    assign RTL___near_mem___dcache$mem_master_awvalid = RTL___near_mem___dcache___mem_master_awvalid;
    assign RTL___near_mem___dcache$mem_master_awid = RTL___near_mem___dcache___mem_master_awid;
    assign RTL___near_mem___dcache$mem_master_awaddr = RTL___near_mem___dcache___mem_master_awaddr;
    assign RTL___near_mem___dcache$mem_master_awlen = RTL___near_mem___dcache___mem_master_awlen;
    assign RTL___near_mem___dcache$mem_master_awsize = RTL___near_mem___dcache___mem_master_awsize;
    assign RTL___near_mem___dcache$mem_master_awburst = RTL___near_mem___dcache___mem_master_awburst;
    assign RTL___near_mem___dcache$mem_master_awlock = RTL___near_mem___dcache___mem_master_awlock;
    assign RTL___near_mem___dcache$mem_master_awcache = RTL___near_mem___dcache___mem_master_awcache;
    assign RTL___near_mem___dcache$mem_master_awprot = RTL___near_mem___dcache___mem_master_awprot;
    assign RTL___near_mem___dcache$mem_master_awqos = RTL___near_mem___dcache___mem_master_awqos;
    assign RTL___near_mem___dcache$mem_master_awregion = RTL___near_mem___dcache___mem_master_awregion;
    assign RTL___near_mem___dcache___mem_master_awready = RTL___near_mem___dcache$mem_master_awready;
    assign RTL___near_mem___dcache$mem_master_wvalid = RTL___near_mem___dcache___mem_master_wvalid;
    assign RTL___near_mem___dcache$mem_master_wdata = RTL___near_mem___dcache___mem_master_wdata;
    assign RTL___near_mem___dcache$mem_master_wstrb = RTL___near_mem___dcache___mem_master_wstrb;
    assign RTL___near_mem___dcache$mem_master_wlast = RTL___near_mem___dcache___mem_master_wlast;
    assign RTL___near_mem___dcache___mem_master_wready = RTL___near_mem___dcache$mem_master_wready;
    assign RTL___near_mem___dcache___mem_master_bvalid = RTL___near_mem___dcache$mem_master_bvalid;
    assign RTL___near_mem___dcache___mem_master_bid = RTL___near_mem___dcache$mem_master_bid;
    assign RTL___near_mem___dcache___mem_master_bresp = RTL___near_mem___dcache$mem_master_bresp;
    assign RTL___near_mem___dcache$mem_master_bready = RTL___near_mem___dcache___mem_master_bready;
    assign RTL___near_mem___dcache$mem_master_arvalid = RTL___near_mem___dcache___mem_master_arvalid;
    assign RTL___near_mem___dcache$mem_master_arid = RTL___near_mem___dcache___mem_master_arid;
    assign RTL___near_mem___dcache$mem_master_araddr = RTL___near_mem___dcache___mem_master_araddr;
    assign RTL___near_mem___dcache$mem_master_arlen = RTL___near_mem___dcache___mem_master_arlen;
    assign RTL___near_mem___dcache$mem_master_arsize = RTL___near_mem___dcache___mem_master_arsize;
    assign RTL___near_mem___dcache$mem_master_arburst = RTL___near_mem___dcache___mem_master_arburst;
    assign RTL___near_mem___dcache$mem_master_arlock = RTL___near_mem___dcache___mem_master_arlock;
    assign RTL___near_mem___dcache$mem_master_arcache = RTL___near_mem___dcache___mem_master_arcache;
    assign RTL___near_mem___dcache$mem_master_arprot = RTL___near_mem___dcache___mem_master_arprot;
    assign RTL___near_mem___dcache$mem_master_arqos = RTL___near_mem___dcache___mem_master_arqos;
    assign RTL___near_mem___dcache$mem_master_arregion = RTL___near_mem___dcache___mem_master_arregion;
    assign RTL___near_mem___dcache___mem_master_arready = RTL___near_mem___dcache$mem_master_arready;
    assign RTL___near_mem___dcache___mem_master_rvalid = RTL___near_mem___dcache$mem_master_rvalid;
    assign RTL___near_mem___dcache___mem_master_rid = RTL___near_mem___dcache$mem_master_rid;
    assign RTL___near_mem___dcache___mem_master_rdata = RTL___near_mem___dcache$mem_master_rdata;
    assign RTL___near_mem___dcache___mem_master_rresp = RTL___near_mem___dcache$mem_master_rresp;
    assign RTL___near_mem___dcache___mem_master_rlast = RTL___near_mem___dcache$mem_master_rlast;
    assign RTL___near_mem___dcache$mem_master_rready = RTL___near_mem___dcache___mem_master_rready;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___icache___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___near_mem___icache___CLK = RTL___near_mem___CLK;
    assign RTL___near_mem___icache___RST_N = RTL___near_mem___RST_N;
    assign RTL___near_mem___icache___set_verbosity_verbosity = RTL___near_mem___icache$set_verbosity_verbosity;
    assign RTL___near_mem___icache___EN_set_verbosity = RTL___near_mem___icache$EN_set_verbosity;
    assign RTL___near_mem___icache___EN_server_reset_request_put = RTL___near_mem___icache$EN_server_reset_request_put;
    assign RTL___near_mem___icache$RDY_server_reset_request_put = RTL___near_mem___icache___RDY_server_reset_request_put;
    assign RTL___near_mem___icache___EN_server_reset_response_get = RTL___near_mem___icache$EN_server_reset_response_get;
    assign RTL___near_mem___icache$RDY_server_reset_response_get = RTL___near_mem___icache___RDY_server_reset_response_get;
    assign RTL___near_mem___icache___req_op = RTL___near_mem___icache$req_op;
    assign RTL___near_mem___icache___req_f3 = RTL___near_mem___icache$req_f3;
    assign RTL___near_mem___icache___req_addr = RTL___near_mem___icache$req_addr;
    assign RTL___near_mem___icache___req_st_value = RTL___near_mem___icache$req_st_value;
    assign RTL___near_mem___icache___req_priv = RTL___near_mem___icache$req_priv;
    assign RTL___near_mem___icache___req_sstatus_SUM = RTL___near_mem___icache$req_sstatus_SUM;
    assign RTL___near_mem___icache___req_mstatus_MXR = RTL___near_mem___icache$req_mstatus_MXR;
    assign RTL___near_mem___icache___req_satp = RTL___near_mem___icache$req_satp;
    assign RTL___near_mem___icache___EN_req = RTL___near_mem___icache$EN_req;
    assign RTL___near_mem___icache$valid = RTL___near_mem___icache___valid;
    assign RTL___near_mem___icache$addr = RTL___near_mem___icache___addr;
    assign RTL___near_mem___icache$word64 = RTL___near_mem___icache___word64;
    assign RTL___near_mem___icache$exc = RTL___near_mem___icache___exc;
    assign RTL___near_mem___icache$exc_code = RTL___near_mem___icache___exc_code;
    assign RTL___near_mem___icache___EN_server_flush_request_put = RTL___near_mem___icache$EN_server_flush_request_put;
    assign RTL___near_mem___icache$RDY_server_flush_request_put = RTL___near_mem___icache___RDY_server_flush_request_put;
    assign RTL___near_mem___icache___EN_server_flush_response_get = RTL___near_mem___icache$EN_server_flush_response_get;
    assign RTL___near_mem___icache$RDY_server_flush_response_get = RTL___near_mem___icache___RDY_server_flush_response_get;
    assign RTL___near_mem___icache___EN_tlb_flush = RTL___near_mem___icache$EN_tlb_flush;
    assign RTL___near_mem___icache$mem_master_awvalid = RTL___near_mem___icache___mem_master_awvalid;
    assign RTL___near_mem___icache$mem_master_awid = RTL___near_mem___icache___mem_master_awid;
    assign RTL___near_mem___icache$mem_master_awaddr = RTL___near_mem___icache___mem_master_awaddr;
    assign RTL___near_mem___icache$mem_master_awlen = RTL___near_mem___icache___mem_master_awlen;
    assign RTL___near_mem___icache$mem_master_awsize = RTL___near_mem___icache___mem_master_awsize;
    assign RTL___near_mem___icache$mem_master_awburst = RTL___near_mem___icache___mem_master_awburst;
    assign RTL___near_mem___icache$mem_master_awlock = RTL___near_mem___icache___mem_master_awlock;
    assign RTL___near_mem___icache$mem_master_awcache = RTL___near_mem___icache___mem_master_awcache;
    assign RTL___near_mem___icache$mem_master_awprot = RTL___near_mem___icache___mem_master_awprot;
    assign RTL___near_mem___icache$mem_master_awqos = RTL___near_mem___icache___mem_master_awqos;
    assign RTL___near_mem___icache$mem_master_awregion = RTL___near_mem___icache___mem_master_awregion;
    assign RTL___near_mem___icache___mem_master_awready = RTL___near_mem___icache$mem_master_awready;
    assign RTL___near_mem___icache$mem_master_wvalid = RTL___near_mem___icache___mem_master_wvalid;
    assign RTL___near_mem___icache$mem_master_wdata = RTL___near_mem___icache___mem_master_wdata;
    assign RTL___near_mem___icache$mem_master_wstrb = RTL___near_mem___icache___mem_master_wstrb;
    assign RTL___near_mem___icache$mem_master_wlast = RTL___near_mem___icache___mem_master_wlast;
    assign RTL___near_mem___icache___mem_master_wready = RTL___near_mem___icache$mem_master_wready;
    assign RTL___near_mem___icache___mem_master_bvalid = RTL___near_mem___icache$mem_master_bvalid;
    assign RTL___near_mem___icache___mem_master_bid = RTL___near_mem___icache$mem_master_bid;
    assign RTL___near_mem___icache___mem_master_bresp = RTL___near_mem___icache$mem_master_bresp;
    assign RTL___near_mem___icache$mem_master_bready = RTL___near_mem___icache___mem_master_bready;
    assign RTL___near_mem___icache$mem_master_arvalid = RTL___near_mem___icache___mem_master_arvalid;
    assign RTL___near_mem___icache$mem_master_arid = RTL___near_mem___icache___mem_master_arid;
    assign RTL___near_mem___icache$mem_master_araddr = RTL___near_mem___icache___mem_master_araddr;
    assign RTL___near_mem___icache$mem_master_arlen = RTL___near_mem___icache___mem_master_arlen;
    assign RTL___near_mem___icache$mem_master_arsize = RTL___near_mem___icache___mem_master_arsize;
    assign RTL___near_mem___icache$mem_master_arburst = RTL___near_mem___icache___mem_master_arburst;
    assign RTL___near_mem___icache$mem_master_arlock = RTL___near_mem___icache___mem_master_arlock;
    assign RTL___near_mem___icache$mem_master_arcache = RTL___near_mem___icache___mem_master_arcache;
    assign RTL___near_mem___icache$mem_master_arprot = RTL___near_mem___icache___mem_master_arprot;
    assign RTL___near_mem___icache$mem_master_arqos = RTL___near_mem___icache___mem_master_arqos;
    assign RTL___near_mem___icache$mem_master_arregion = RTL___near_mem___icache___mem_master_arregion;
    assign RTL___near_mem___icache___mem_master_arready = RTL___near_mem___icache$mem_master_arready;
    assign RTL___near_mem___icache___mem_master_rvalid = RTL___near_mem___icache$mem_master_rvalid;
    assign RTL___near_mem___icache___mem_master_rid = RTL___near_mem___icache$mem_master_rid;
    assign RTL___near_mem___icache___mem_master_rdata = RTL___near_mem___icache$mem_master_rdata;
    assign RTL___near_mem___icache___mem_master_rresp = RTL___near_mem___icache$mem_master_rresp;
    assign RTL___near_mem___icache___mem_master_rlast = RTL___near_mem___icache$mem_master_rlast;
    assign RTL___near_mem___icache$mem_master_rready = RTL___near_mem___icache___mem_master_rready;
      
    
    wire[63:0] RTL___near_mem___soc_map___m_boot_rom_addr_base , RTL___near_mem___soc_map___m_boot_rom_addr_lim , RTL___near_mem___soc_map___m_boot_rom_addr_size , RTL___near_mem___soc_map___m_mem0_controller_addr_base , RTL___near_mem___soc_map___m_mem0_controller_addr_lim , RTL___near_mem___soc_map___m_mem0_controller_addr_size , RTL___near_mem___soc_map___m_mtvec_reset_value , RTL___near_mem___soc_map___m_near_mem_io_addr_base , RTL___near_mem___soc_map___m_near_mem_io_addr_lim , RTL___near_mem___soc_map___m_near_mem_io_addr_size , RTL___near_mem___soc_map___m_nmivec_reset_value , RTL___near_mem___soc_map___m_pc_reset_value , RTL___near_mem___soc_map___m_plic_addr_base , RTL___near_mem___soc_map___m_plic_addr_lim , RTL___near_mem___soc_map___m_plic_addr_size , RTL___near_mem___soc_map___m_tcm_addr_base , RTL___near_mem___soc_map___m_tcm_addr_lim , RTL___near_mem___soc_map___m_tcm_addr_size , RTL___near_mem___soc_map___m_uart0_addr_base , RTL___near_mem___soc_map___m_uart0_addr_lim , RTL___near_mem___soc_map___m_uart0_addr_size ; 
    wire RTL___near_mem___soc_map___m_is_IO_addr , RTL___near_mem___soc_map___m_is_mem_addr , RTL___near_mem___soc_map___m_is_near_mem_IO_addr ; 
  assign  RTL___near_mem___soc_map___m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL___near_mem___soc_map___m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL___near_mem___soc_map___m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL___near_mem___soc_map___m_plic_addr_base =64'h000000000C000000; 
  assign  RTL___near_mem___soc_map___m_plic_addr_size =64'h0000000000400000; 
  assign  RTL___near_mem___soc_map___m_plic_addr_lim =64'd205520896; 
  assign  RTL___near_mem___soc_map___m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL___near_mem___soc_map___m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL___near_mem___soc_map___m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL___near_mem___soc_map___m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL___near_mem___soc_map___m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL___near_mem___soc_map___m_boot_rom_addr_lim =64'd8192; 
  assign  RTL___near_mem___soc_map___m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL___near_mem___soc_map___m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL___near_mem___soc_map___m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL___near_mem___soc_map___m_tcm_addr_base =64'h0; 
  assign  RTL___near_mem___soc_map___m_tcm_addr_size =64'd0; 
  assign  RTL___near_mem___soc_map___m_tcm_addr_lim =64'd0; 
  assign  RTL___near_mem___soc_map___m_is_mem_addr = RTL___near_mem___soc_map___m_is_mem_addr_addr >=64'h0000000000001000&& RTL___near_mem___soc_map___m_is_mem_addr_addr <64'd8192|| RTL___near_mem___soc_map___m_is_mem_addr_addr >=64'h0000000080000000&& RTL___near_mem___soc_map___m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL___near_mem___soc_map___m_is_IO_addr = RTL___near_mem___soc_map___m_is_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___soc_map___m_is_IO_addr_addr <64'd33603584|| RTL___near_mem___soc_map___m_is_IO_addr_addr >=64'h000000000C000000&& RTL___near_mem___soc_map___m_is_IO_addr_addr <64'd205520896|| RTL___near_mem___soc_map___m_is_IO_addr_addr >=64'h00000000C0000000&& RTL___near_mem___soc_map___m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL___near_mem___soc_map___m_is_near_mem_IO_addr = RTL___near_mem___soc_map___m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL___near_mem___soc_map___m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL___near_mem___soc_map___m_pc_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___soc_map___m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL___near_mem___soc_map___m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
    assign RTL___near_mem___dcache___soc_map___CLK = RTL___near_mem___dcache___CLK;
    assign RTL___near_mem___dcache___soc_map___RST_N = RTL___near_mem___dcache___RST_N;
    assign RTL___near_mem___dcache___soc_map___m_is_mem_addr_addr = RTL___near_mem___dcache___soc_map$m_is_mem_addr_addr;
    assign RTL___near_mem___dcache___soc_map$m_is_mem_addr = RTL___near_mem___dcache___soc_map___m_is_mem_addr;
    assign RTL___near_mem___dcache___soc_map___m_is_IO_addr_addr = RTL___near_mem___dcache___soc_map$m_is_IO_addr_addr;
    assign RTL___near_mem___dcache___soc_map___m_is_near_mem_IO_addr_addr = RTL___near_mem___dcache___soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL___near_mem___icache___soc_map___CLK = RTL___near_mem___icache___CLK;
    assign RTL___near_mem___icache___soc_map___RST_N = RTL___near_mem___icache___RST_N;
    assign RTL___near_mem___icache___soc_map___m_is_mem_addr_addr = RTL___near_mem___icache___soc_map$m_is_mem_addr_addr;
    assign RTL___near_mem___icache___soc_map$m_is_mem_addr = RTL___near_mem___icache___soc_map___m_is_mem_addr;
    assign RTL___near_mem___icache___soc_map___m_is_IO_addr_addr = RTL___near_mem___icache___soc_map$m_is_IO_addr_addr;
    assign RTL___near_mem___icache___soc_map___m_is_near_mem_IO_addr_addr = RTL___near_mem___icache___soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL___near_mem___soc_map___CLK = RTL___near_mem___CLK;
    assign RTL___near_mem___soc_map___RST_N = RTL___near_mem___RST_N;
    assign RTL___near_mem___soc_map___m_is_mem_addr_addr = RTL___near_mem___soc_map$m_is_mem_addr_addr;
    assign RTL___near_mem___soc_map___m_is_IO_addr_addr = RTL___near_mem___soc_map$m_is_IO_addr_addr;
    assign RTL___near_mem___soc_map___m_is_near_mem_IO_addr_addr = RTL___near_mem___soc_map$m_is_near_mem_IO_addr_addr;
     
  assign  RTL___near_mem___CAN_FIRE_RL_rl_reset = RTL___near_mem___dcache$RDY_server_reset_request_put && RTL___near_mem___icache$RDY_server_reset_request_put && RTL___near_mem___rg_state ==2'd0; 
  assign  RTL___near_mem___WILL_FIRE_RL_rl_reset = RTL___near_mem___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___CAN_FIRE_RL_rl_reset_complete = RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___WILL_FIRE_RL_rl_reset_complete = RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___MUX_rg_state$write_1__SEL_2 = RTL___near_mem___CAN_FIRE_RL_rl_reset &&! RTL___near_mem___EN_server_fence_request_put &&! RTL___near_mem___EN_server_fence_i_request_put ; 
  assign  RTL___near_mem___MUX_rg_state$write_1__SEL_3 = RTL___near_mem___dcache$RDY_server_reset_response_get && RTL___near_mem___icache$RDY_server_reset_response_get && RTL___near_mem___f_reset_rsps$FULL_N && RTL___near_mem___rg_state ==2'd1; 
  assign  RTL___near_mem___cfg_verbosity$D_IN =4'h0; 
  assign  RTL___near_mem___cfg_verbosity$EN =1'b0; 
  always @(    RTL___near_mem___EN_server_reset_request_put              or   RTL___near_mem___WILL_FIRE_RL_rl_reset           or   RTL___near_mem___WILL_FIRE_RL_rl_reset_complete  )
         begin 
             case (1'b1) 
              RTL___near_mem___EN_server_reset_request_put  : 
                  RTL___near_mem___rg_state$D_IN  =2'd0; 
              RTL___near_mem___WILL_FIRE_RL_rl_reset  : 
                  RTL___near_mem___rg_state$D_IN  =2'd1; 
              RTL___near_mem___WILL_FIRE_RL_rl_reset_complete  : 
                  RTL___near_mem___rg_state$D_IN  =2'd2;
              default : 
                  RTL___near_mem___rg_state$D_IN  =2'b10;endcase
         end
  assign  RTL___near_mem___rg_state$EN = RTL___near_mem___EN_server_reset_request_put || RTL___near_mem___WILL_FIRE_RL_rl_reset || RTL___near_mem___WILL_FIRE_RL_rl_reset_complete ; 
  assign  RTL___near_mem___dcache$mem_master_arready = RTL___near_mem___dmem_master_arready ; 
  assign  RTL___near_mem___dcache$mem_master_awready = RTL___near_mem___dmem_master_awready ; 
  assign  RTL___near_mem___dcache$mem_master_bid = RTL___near_mem___dmem_master_bid ; 
  assign  RTL___near_mem___dcache$mem_master_bresp = RTL___near_mem___dmem_master_bresp ; 
  assign  RTL___near_mem___dcache$mem_master_bvalid = RTL___near_mem___dmem_master_bvalid ; 
  assign  RTL___near_mem___dcache$mem_master_rdata = RTL___near_mem___dmem_master_rdata ; 
  assign  RTL___near_mem___dcache$mem_master_rid = RTL___near_mem___dmem_master_rid ; 
  assign  RTL___near_mem___dcache$mem_master_rlast = RTL___near_mem___dmem_master_rlast ; 
  assign  RTL___near_mem___dcache$mem_master_rresp = RTL___near_mem___dmem_master_rresp ; 
  assign  RTL___near_mem___dcache$mem_master_rvalid = RTL___near_mem___dmem_master_rvalid ; 
  assign  RTL___near_mem___dcache$mem_master_wready = RTL___near_mem___dmem_master_wready ; 
  assign  RTL___near_mem___dcache$req_addr = RTL___near_mem___dmem_req_addr ; 
  assign  RTL___near_mem___dcache$req_f3 = RTL___near_mem___dmem_req_f3 ; 
  assign  RTL___near_mem___dcache$req_mstatus_MXR = RTL___near_mem___dmem_req_mstatus_MXR ; 
  assign  RTL___near_mem___dcache$req_op = RTL___near_mem___dmem_req_op ; 
  assign  RTL___near_mem___dcache$req_priv = RTL___near_mem___dmem_req_priv ; 
  assign  RTL___near_mem___dcache$req_satp = RTL___near_mem___dmem_req_satp ; 
  assign  RTL___near_mem___dcache$req_sstatus_SUM = RTL___near_mem___dmem_req_sstatus_SUM ; 
  assign  RTL___near_mem___dcache$req_st_value = RTL___near_mem___dmem_req_store_value ; 
  assign  RTL___near_mem___dcache$set_verbosity_verbosity =4'h0; 
  assign  RTL___near_mem___dcache$EN_set_verbosity =1'b0; 
  assign  RTL___near_mem___dcache$EN_server_reset_request_put = RTL___near_mem___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___dcache$EN_server_reset_response_get = RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___dcache$EN_req = RTL___near_mem___EN_dmem_req ; 
  assign  RTL___near_mem___dcache$EN_server_flush_request_put = RTL___near_mem___EN_server_fence_i_request_put || RTL___near_mem___EN_server_fence_request_put ; 
  assign  RTL___near_mem___dcache$EN_server_flush_response_get = RTL___near_mem___EN_server_fence_i_response_get || RTL___near_mem___EN_server_fence_response_get ; 
  assign  RTL___near_mem___dcache$EN_tlb_flush = RTL___near_mem___EN_sfence_vma ; 
  assign  RTL___near_mem___f_reset_rsps$ENQ = RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___f_reset_rsps$DEQ = RTL___near_mem___EN_server_reset_response_get ; 
  assign  RTL___near_mem___f_reset_rsps$CLR =1'b0; 
  assign  RTL___near_mem___icache$mem_master_arready = RTL___near_mem___imem_master_arready ; 
  assign  RTL___near_mem___icache$mem_master_awready = RTL___near_mem___imem_master_awready ; 
  assign  RTL___near_mem___icache$mem_master_bid = RTL___near_mem___imem_master_bid ; 
  assign  RTL___near_mem___icache$mem_master_bresp = RTL___near_mem___imem_master_bresp ; 
  assign  RTL___near_mem___icache$mem_master_bvalid = RTL___near_mem___imem_master_bvalid ; 
  assign  RTL___near_mem___icache$mem_master_rdata = RTL___near_mem___imem_master_rdata ; 
  assign  RTL___near_mem___icache$mem_master_rid = RTL___near_mem___imem_master_rid ; 
  assign  RTL___near_mem___icache$mem_master_rlast = RTL___near_mem___imem_master_rlast ; 
  assign  RTL___near_mem___icache$mem_master_rresp = RTL___near_mem___imem_master_rresp ; 
  assign  RTL___near_mem___icache$mem_master_rvalid = RTL___near_mem___imem_master_rvalid ; 
  assign  RTL___near_mem___icache$mem_master_wready = RTL___near_mem___imem_master_wready ; 
  assign  RTL___near_mem___icache$req_addr = RTL___near_mem___imem_req_addr ; 
  assign  RTL___near_mem___icache$req_f3 = RTL___near_mem___imem_req_f3 ; 
  assign  RTL___near_mem___icache$req_mstatus_MXR = RTL___near_mem___imem_req_mstatus_MXR ; 
  assign  RTL___near_mem___icache$req_op =1'd0; 
  assign  RTL___near_mem___icache$req_priv = RTL___near_mem___imem_req_priv ; 
  assign  RTL___near_mem___icache$req_satp = RTL___near_mem___imem_req_satp ; 
  assign  RTL___near_mem___icache$req_sstatus_SUM = RTL___near_mem___imem_req_sstatus_SUM ; 
  assign  RTL___near_mem___icache$req_st_value =64'hAAAAAAAAAAAAAAAA; 
  assign  RTL___near_mem___icache$set_verbosity_verbosity =4'h0; 
  assign  RTL___near_mem___icache$EN_set_verbosity =1'b0; 
  assign  RTL___near_mem___icache$EN_server_reset_request_put = RTL___near_mem___MUX_rg_state$write_1__SEL_2 ; 
  assign  RTL___near_mem___icache$EN_server_reset_response_get = RTL___near_mem___MUX_rg_state$write_1__SEL_3 ; 
  assign  RTL___near_mem___icache$EN_req = RTL___near_mem___EN_imem_req ; 
  assign  RTL___near_mem___icache$EN_server_flush_request_put = RTL___near_mem___EN_server_fence_i_request_put ; 
  assign  RTL___near_mem___icache$EN_server_flush_response_get = RTL___near_mem___EN_server_fence_i_response_get ; 
  assign  RTL___near_mem___icache$EN_tlb_flush = RTL___near_mem___EN_sfence_vma ; 
  assign  RTL___near_mem___soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL___near_mem___soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 = RTL___near_mem___cfg_verbosity >4'd1; 
  always @( posedge  RTL___near_mem___CLK )
         begin 
             if ( RTL___near_mem___RST_N ==1'b0)
                 begin  
                     RTL___near_mem___cfg_verbosity  <=4'd0; 
                     RTL___near_mem___rg_state  <=2'd2;
                 end 
              else 
                 begin 
                     if ( RTL___near_mem___cfg_verbosity$EN ) 
                         RTL___near_mem___cfg_verbosity  <= RTL___near_mem___cfg_verbosity$D_IN ;
                     if ( RTL___near_mem___rg_state$EN ) 
                         RTL___near_mem___rg_state  <= RTL___near_mem___rg_state$D_IN ;
                 end 
         end
  always @( negedge  RTL___near_mem___CLK )
         begin #0;
             if ( RTL___near_mem___RST_N !=1'b0)
                 if ( RTL___near_mem___WILL_FIRE_RL_rl_reset && RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 )
                     begin  
                         RTL___near_mem___v__h1643  =$stime;#0;
                     end  
             RTL___near_mem___v__h1637  = RTL___near_mem___v__h1643 /32'd10;
             if ( RTL___near_mem___RST_N !=1'b0)
                 if ( RTL___near_mem___WILL_FIRE_RL_rl_reset && RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 )$display("%0d: Near_Mem.rl_reset", RTL___near_mem___v__h1637 );
             if ( RTL___near_mem___RST_N !=1'b0)
                 if ( RTL___near_mem___WILL_FIRE_RL_rl_reset_complete && RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 )
                     begin  
                         RTL___near_mem___v__h1794  =$stime;#0;
                     end  
             RTL___near_mem___v__h1788  = RTL___near_mem___v__h1794 /32'd10;
             if ( RTL___near_mem___RST_N !=1'b0)
                 if ( RTL___near_mem___WILL_FIRE_RL_rl_reset_complete && RTL___near_mem___NOT_cfg_verbosity_read_ULE_1___d9 )$display("%0d: Near_Mem.rl_reset_complete", RTL___near_mem___v__h1788 );
         end
 
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL___near_mem___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___near_mem___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL___near_mem___CLK = RTL___CLK;
    assign RTL___near_mem___RST_N = RTL___RST_N;
    assign RTL___near_mem___EN_server_reset_request_put = RTL___near_mem$EN_server_reset_request_put;
    assign RTL___near_mem$RDY_server_reset_request_put = RTL___near_mem___RDY_server_reset_request_put;
    assign RTL___near_mem___EN_server_reset_response_get = RTL___near_mem$EN_server_reset_response_get;
    assign RTL___near_mem$RDY_server_reset_response_get = RTL___near_mem___RDY_server_reset_response_get;
    assign RTL___near_mem___imem_req_f3 = RTL___near_mem$imem_req_f3;
    assign RTL___near_mem___imem_req_addr = RTL___near_mem$imem_req_addr;
    assign RTL___near_mem___imem_req_priv = RTL___near_mem$imem_req_priv;
    assign RTL___near_mem___imem_req_sstatus_SUM = RTL___near_mem$imem_req_sstatus_SUM;
    assign RTL___near_mem___imem_req_mstatus_MXR = RTL___near_mem$imem_req_mstatus_MXR;
    assign RTL___near_mem___imem_req_satp = RTL___near_mem$imem_req_satp;
    assign RTL___near_mem___EN_imem_req = RTL___near_mem$EN_imem_req;
    assign RTL___near_mem$imem_valid = RTL___near_mem___imem_valid;
    assign RTL___near_mem$imem_is_i32_not_i16 = RTL___near_mem___imem_is_i32_not_i16;
    assign RTL___near_mem$imem_pc = RTL___near_mem___imem_pc;
    assign RTL___near_mem$imem_instr = RTL___near_mem___imem_instr;
    assign RTL___near_mem$imem_exc = RTL___near_mem___imem_exc;
    assign RTL___near_mem$imem_exc_code = RTL___near_mem___imem_exc_code;
    assign RTL___near_mem$imem_tval = RTL___near_mem___imem_tval;
    assign RTL___near_mem$imem_master_awvalid = RTL___near_mem___imem_master_awvalid;
    assign RTL___near_mem$imem_master_awid = RTL___near_mem___imem_master_awid;
    assign RTL___near_mem$imem_master_awaddr = RTL___near_mem___imem_master_awaddr;
    assign RTL___near_mem$imem_master_awlen = RTL___near_mem___imem_master_awlen;
    assign RTL___near_mem$imem_master_awsize = RTL___near_mem___imem_master_awsize;
    assign RTL___near_mem$imem_master_awburst = RTL___near_mem___imem_master_awburst;
    assign RTL___near_mem$imem_master_awlock = RTL___near_mem___imem_master_awlock;
    assign RTL___near_mem$imem_master_awcache = RTL___near_mem___imem_master_awcache;
    assign RTL___near_mem$imem_master_awprot = RTL___near_mem___imem_master_awprot;
    assign RTL___near_mem$imem_master_awqos = RTL___near_mem___imem_master_awqos;
    assign RTL___near_mem$imem_master_awregion = RTL___near_mem___imem_master_awregion;
    assign RTL___near_mem___imem_master_awready = RTL___near_mem$imem_master_awready;
    assign RTL___near_mem$imem_master_wvalid = RTL___near_mem___imem_master_wvalid;
    assign RTL___near_mem$imem_master_wdata = RTL___near_mem___imem_master_wdata;
    assign RTL___near_mem$imem_master_wstrb = RTL___near_mem___imem_master_wstrb;
    assign RTL___near_mem$imem_master_wlast = RTL___near_mem___imem_master_wlast;
    assign RTL___near_mem___imem_master_wready = RTL___near_mem$imem_master_wready;
    assign RTL___near_mem___imem_master_bvalid = RTL___near_mem$imem_master_bvalid;
    assign RTL___near_mem___imem_master_bid = RTL___near_mem$imem_master_bid;
    assign RTL___near_mem___imem_master_bresp = RTL___near_mem$imem_master_bresp;
    assign RTL___near_mem$imem_master_bready = RTL___near_mem___imem_master_bready;
    assign RTL___near_mem$imem_master_arvalid = RTL___near_mem___imem_master_arvalid;
    assign RTL___near_mem$imem_master_arid = RTL___near_mem___imem_master_arid;
    assign RTL___near_mem$imem_master_araddr = RTL___near_mem___imem_master_araddr;
    assign RTL___near_mem$imem_master_arlen = RTL___near_mem___imem_master_arlen;
    assign RTL___near_mem$imem_master_arsize = RTL___near_mem___imem_master_arsize;
    assign RTL___near_mem$imem_master_arburst = RTL___near_mem___imem_master_arburst;
    assign RTL___near_mem$imem_master_arlock = RTL___near_mem___imem_master_arlock;
    assign RTL___near_mem$imem_master_arcache = RTL___near_mem___imem_master_arcache;
    assign RTL___near_mem$imem_master_arprot = RTL___near_mem___imem_master_arprot;
    assign RTL___near_mem$imem_master_arqos = RTL___near_mem___imem_master_arqos;
    assign RTL___near_mem$imem_master_arregion = RTL___near_mem___imem_master_arregion;
    assign RTL___near_mem___imem_master_arready = RTL___near_mem$imem_master_arready;
    assign RTL___near_mem___imem_master_rvalid = RTL___near_mem$imem_master_rvalid;
    assign RTL___near_mem___imem_master_rid = RTL___near_mem$imem_master_rid;
    assign RTL___near_mem___imem_master_rdata = RTL___near_mem$imem_master_rdata;
    assign RTL___near_mem___imem_master_rresp = RTL___near_mem$imem_master_rresp;
    assign RTL___near_mem___imem_master_rlast = RTL___near_mem$imem_master_rlast;
    assign RTL___near_mem$imem_master_rready = RTL___near_mem___imem_master_rready;
    assign RTL___near_mem___dmem_req_op = RTL___near_mem$dmem_req_op;
    assign RTL___near_mem___dmem_req_f3 = RTL___near_mem$dmem_req_f3;
    assign RTL___near_mem___dmem_req_addr = RTL___near_mem$dmem_req_addr;
    assign RTL___near_mem___dmem_req_store_value = RTL___near_mem$dmem_req_store_value;
    assign RTL___near_mem___dmem_req_priv = RTL___near_mem$dmem_req_priv;
    assign RTL___near_mem___dmem_req_sstatus_SUM = RTL___near_mem$dmem_req_sstatus_SUM;
    assign RTL___near_mem___dmem_req_mstatus_MXR = RTL___near_mem$dmem_req_mstatus_MXR;
    assign RTL___near_mem___dmem_req_satp = RTL___near_mem$dmem_req_satp;
    assign RTL___near_mem___EN_dmem_req = RTL___near_mem$EN_dmem_req;
    assign RTL___near_mem$dmem_valid = RTL___near_mem___dmem_valid;
    assign RTL___near_mem$dmem_word64 = RTL___near_mem___dmem_word64;
    assign RTL___near_mem$dmem_exc = RTL___near_mem___dmem_exc;
    assign RTL___near_mem$dmem_exc_code = RTL___near_mem___dmem_exc_code;
    assign RTL___near_mem$dmem_master_awvalid = RTL___near_mem___dmem_master_awvalid;
    assign RTL___near_mem$dmem_master_awid = RTL___near_mem___dmem_master_awid;
    assign RTL___near_mem$dmem_master_awaddr = RTL___near_mem___dmem_master_awaddr;
    assign RTL___near_mem$dmem_master_awlen = RTL___near_mem___dmem_master_awlen;
    assign RTL___near_mem$dmem_master_awsize = RTL___near_mem___dmem_master_awsize;
    assign RTL___near_mem$dmem_master_awburst = RTL___near_mem___dmem_master_awburst;
    assign RTL___near_mem$dmem_master_awlock = RTL___near_mem___dmem_master_awlock;
    assign RTL___near_mem$dmem_master_awcache = RTL___near_mem___dmem_master_awcache;
    assign RTL___near_mem$dmem_master_awprot = RTL___near_mem___dmem_master_awprot;
    assign RTL___near_mem$dmem_master_awqos = RTL___near_mem___dmem_master_awqos;
    assign RTL___near_mem$dmem_master_awregion = RTL___near_mem___dmem_master_awregion;
    assign RTL___near_mem___dmem_master_awready = RTL___near_mem$dmem_master_awready;
    assign RTL___near_mem$dmem_master_wvalid = RTL___near_mem___dmem_master_wvalid;
    assign RTL___near_mem$dmem_master_wdata = RTL___near_mem___dmem_master_wdata;
    assign RTL___near_mem$dmem_master_wstrb = RTL___near_mem___dmem_master_wstrb;
    assign RTL___near_mem$dmem_master_wlast = RTL___near_mem___dmem_master_wlast;
    assign RTL___near_mem___dmem_master_wready = RTL___near_mem$dmem_master_wready;
    assign RTL___near_mem___dmem_master_bvalid = RTL___near_mem$dmem_master_bvalid;
    assign RTL___near_mem___dmem_master_bid = RTL___near_mem$dmem_master_bid;
    assign RTL___near_mem___dmem_master_bresp = RTL___near_mem$dmem_master_bresp;
    assign RTL___near_mem$dmem_master_bready = RTL___near_mem___dmem_master_bready;
    assign RTL___near_mem$dmem_master_arvalid = RTL___near_mem___dmem_master_arvalid;
    assign RTL___near_mem$dmem_master_arid = RTL___near_mem___dmem_master_arid;
    assign RTL___near_mem$dmem_master_araddr = RTL___near_mem___dmem_master_araddr;
    assign RTL___near_mem$dmem_master_arlen = RTL___near_mem___dmem_master_arlen;
    assign RTL___near_mem$dmem_master_arsize = RTL___near_mem___dmem_master_arsize;
    assign RTL___near_mem$dmem_master_arburst = RTL___near_mem___dmem_master_arburst;
    assign RTL___near_mem$dmem_master_arlock = RTL___near_mem___dmem_master_arlock;
    assign RTL___near_mem$dmem_master_arcache = RTL___near_mem___dmem_master_arcache;
    assign RTL___near_mem$dmem_master_arprot = RTL___near_mem___dmem_master_arprot;
    assign RTL___near_mem$dmem_master_arqos = RTL___near_mem___dmem_master_arqos;
    assign RTL___near_mem$dmem_master_arregion = RTL___near_mem___dmem_master_arregion;
    assign RTL___near_mem___dmem_master_arready = RTL___near_mem$dmem_master_arready;
    assign RTL___near_mem___dmem_master_rvalid = RTL___near_mem$dmem_master_rvalid;
    assign RTL___near_mem___dmem_master_rid = RTL___near_mem$dmem_master_rid;
    assign RTL___near_mem___dmem_master_rdata = RTL___near_mem$dmem_master_rdata;
    assign RTL___near_mem___dmem_master_rresp = RTL___near_mem$dmem_master_rresp;
    assign RTL___near_mem___dmem_master_rlast = RTL___near_mem$dmem_master_rlast;
    assign RTL___near_mem$dmem_master_rready = RTL___near_mem___dmem_master_rready;
    assign RTL___near_mem___EN_server_fence_i_request_put = RTL___near_mem$EN_server_fence_i_request_put;
    assign RTL___near_mem$RDY_server_fence_i_request_put = RTL___near_mem___RDY_server_fence_i_request_put;
    assign RTL___near_mem___EN_server_fence_i_response_get = RTL___near_mem$EN_server_fence_i_response_get;
    assign RTL___near_mem$RDY_server_fence_i_response_get = RTL___near_mem___RDY_server_fence_i_response_get;
    assign RTL___near_mem___server_fence_request_put = RTL___near_mem$server_fence_request_put;
    assign RTL___near_mem___EN_server_fence_request_put = RTL___near_mem$EN_server_fence_request_put;
    assign RTL___near_mem$RDY_server_fence_request_put = RTL___near_mem___RDY_server_fence_request_put;
    assign RTL___near_mem___EN_server_fence_response_get = RTL___near_mem$EN_server_fence_response_get;
    assign RTL___near_mem$RDY_server_fence_response_get = RTL___near_mem___RDY_server_fence_response_get;
    assign RTL___near_mem___EN_sfence_vma = RTL___near_mem$EN_sfence_vma;
      
    
    wire[63:0] RTL___soc_map___m_boot_rom_addr_base , RTL___soc_map___m_boot_rom_addr_lim , RTL___soc_map___m_boot_rom_addr_size , RTL___soc_map___m_mem0_controller_addr_base , RTL___soc_map___m_mem0_controller_addr_lim , RTL___soc_map___m_mem0_controller_addr_size , RTL___soc_map___m_mtvec_reset_value , RTL___soc_map___m_near_mem_io_addr_base , RTL___soc_map___m_near_mem_io_addr_lim , RTL___soc_map___m_near_mem_io_addr_size , RTL___soc_map___m_nmivec_reset_value , RTL___soc_map___m_pc_reset_value , RTL___soc_map___m_plic_addr_base , RTL___soc_map___m_plic_addr_lim , RTL___soc_map___m_plic_addr_size , RTL___soc_map___m_tcm_addr_base , RTL___soc_map___m_tcm_addr_lim , RTL___soc_map___m_tcm_addr_size , RTL___soc_map___m_uart0_addr_base , RTL___soc_map___m_uart0_addr_lim , RTL___soc_map___m_uart0_addr_size ; 
    wire RTL___soc_map___m_is_IO_addr , RTL___soc_map___m_is_mem_addr , RTL___soc_map___m_is_near_mem_IO_addr ; 
  assign  RTL___soc_map___m_near_mem_io_addr_base =64'h0000000002000000; 
  assign  RTL___soc_map___m_near_mem_io_addr_size =64'h000000000000C000; 
  assign  RTL___soc_map___m_near_mem_io_addr_lim =64'd33603584; 
  assign  RTL___soc_map___m_plic_addr_base =64'h000000000C000000; 
  assign  RTL___soc_map___m_plic_addr_size =64'h0000000000400000; 
  assign  RTL___soc_map___m_plic_addr_lim =64'd205520896; 
  assign  RTL___soc_map___m_uart0_addr_base =64'h00000000C0000000; 
  assign  RTL___soc_map___m_uart0_addr_size =64'h0000000000000080; 
  assign  RTL___soc_map___m_uart0_addr_lim =64'h00000000C0000080; 
  assign  RTL___soc_map___m_boot_rom_addr_base =64'h0000000000001000; 
  assign  RTL___soc_map___m_boot_rom_addr_size =64'h0000000000001000; 
  assign  RTL___soc_map___m_boot_rom_addr_lim =64'd8192; 
  assign  RTL___soc_map___m_mem0_controller_addr_base =64'h0000000080000000; 
  assign  RTL___soc_map___m_mem0_controller_addr_size =64'h0000000010000000; 
  assign  RTL___soc_map___m_mem0_controller_addr_lim =64'h0000000090000000; 
  assign  RTL___soc_map___m_tcm_addr_base =64'h0; 
  assign  RTL___soc_map___m_tcm_addr_size =64'd0; 
  assign  RTL___soc_map___m_tcm_addr_lim =64'd0; 
  assign  RTL___soc_map___m_is_mem_addr = RTL___soc_map___m_is_mem_addr_addr >=64'h0000000000001000&& RTL___soc_map___m_is_mem_addr_addr <64'd8192|| RTL___soc_map___m_is_mem_addr_addr >=64'h0000000080000000&& RTL___soc_map___m_is_mem_addr_addr <64'h0000000090000000; 
  assign  RTL___soc_map___m_is_IO_addr = RTL___soc_map___m_is_IO_addr_addr >=64'h0000000002000000&& RTL___soc_map___m_is_IO_addr_addr <64'd33603584|| RTL___soc_map___m_is_IO_addr_addr >=64'h000000000C000000&& RTL___soc_map___m_is_IO_addr_addr <64'd205520896|| RTL___soc_map___m_is_IO_addr_addr >=64'h00000000C0000000&& RTL___soc_map___m_is_IO_addr_addr <64'h00000000C0000080; 
  assign  RTL___soc_map___m_is_near_mem_IO_addr = RTL___soc_map___m_is_near_mem_IO_addr_addr >=64'h0000000002000000&& RTL___soc_map___m_is_near_mem_IO_addr_addr <64'd33603584; 
  assign  RTL___soc_map___m_pc_reset_value =64'h0000000000001000; 
  assign  RTL___soc_map___m_mtvec_reset_value =64'h0000000000001000; 
  assign  RTL___soc_map___m_nmivec_reset_value =64'hAAAAAAAAAAAAAAAA;
    assign RTL___csr_regfile___soc_map___CLK = RTL___csr_regfile___CLK;
    assign RTL___csr_regfile___soc_map___RST_N = RTL___csr_regfile___RST_N;
    assign RTL___csr_regfile___soc_map___m_is_mem_addr_addr = RTL___csr_regfile___soc_map$m_is_mem_addr_addr;
    assign RTL___csr_regfile___soc_map___m_is_IO_addr_addr = RTL___csr_regfile___soc_map$m_is_IO_addr_addr;
    assign RTL___csr_regfile___soc_map___m_is_near_mem_IO_addr_addr = RTL___csr_regfile___soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL___csr_regfile___soc_map$m_mtvec_reset_value = RTL___csr_regfile___soc_map___m_mtvec_reset_value;
    assign RTL___csr_regfile___soc_map$m_nmivec_reset_value = RTL___csr_regfile___soc_map___m_nmivec_reset_value;
    assign RTL___soc_map___CLK = RTL___CLK;
    assign RTL___soc_map___RST_N = RTL___RST_N;
    assign RTL___soc_map___m_is_mem_addr_addr = RTL___soc_map$m_is_mem_addr_addr;
    assign RTL___soc_map___m_is_IO_addr_addr = RTL___soc_map$m_is_IO_addr_addr;
    assign RTL___soc_map___m_is_near_mem_IO_addr_addr = RTL___soc_map$m_is_near_mem_IO_addr_addr;
    assign RTL___soc_map$m_pc_reset_value = RTL___soc_map___m_pc_reset_value;
      
    
    reg RTL___stage1_f_reset_reqs___empty_reg ; 
    reg RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___FULL_N = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___EMPTY_N = RTL___stage1_f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___stage1_f_reset_reqs___CLK )
         begin 
             if ( RTL___stage1_f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___stage1_f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___stage1_f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage1_f_reset_reqs___CLR )
                         begin  
                             RTL___stage1_f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___stage1_f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage1_f_reset_reqs___ENQ &&! RTL___stage1_f_reset_reqs___DEQ )
                             begin  
                                 RTL___stage1_f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___stage1_f_reset_reqs___full_reg  <=! RTL___stage1_f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage1_f_reset_reqs___ENQ && RTL___stage1_f_reset_reqs___DEQ )
                                 begin  
                                     RTL___stage1_f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___stage1_f_reset_reqs___empty_reg  <=! RTL___stage1_f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage1_f_reset_reqs___CLK )
         begin : RTL___stage1_f_reset_reqs___error_checks 
           reg RTL___stage1_f_reset_reqs___deqerror , RTL___stage1_f_reset_reqs___enqerror ; 
             RTL___stage1_f_reset_reqs___deqerror  =0; 
             RTL___stage1_f_reset_reqs___enqerror  =0;
             if ( RTL___stage1_f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___stage1_f_reset_reqs___empty_reg && RTL___stage1_f_reset_reqs___DEQ )
                         begin  
                             RTL___stage1_f_reset_reqs___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage1_f_reset_reqs___full_reg && RTL___stage1_f_reset_reqs___ENQ &&(! RTL___stage1_f_reset_reqs___DEQ || RTL___stage1_f_reset_reqs___guarded ))
                         begin  
                             RTL___stage1_f_reset_reqs___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_reqs___full_reg ; 
  assign  RTL___stage1_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_reqs___empty_reg ;
    reg RTL___stage1_f_reset_rsps___empty_reg ; 
    reg RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___FULL_N = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___EMPTY_N = RTL___stage1_f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___stage1_f_reset_rsps___CLK )
         begin 
             if ( RTL___stage1_f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___stage1_f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___stage1_f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage1_f_reset_rsps___CLR )
                         begin  
                             RTL___stage1_f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___stage1_f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage1_f_reset_rsps___ENQ &&! RTL___stage1_f_reset_rsps___DEQ )
                             begin  
                                 RTL___stage1_f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___stage1_f_reset_rsps___full_reg  <=! RTL___stage1_f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage1_f_reset_rsps___ENQ && RTL___stage1_f_reset_rsps___DEQ )
                                 begin  
                                     RTL___stage1_f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___stage1_f_reset_rsps___empty_reg  <=! RTL___stage1_f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage1_f_reset_rsps___CLK )
         begin : RTL___stage1_f_reset_rsps___error_checks 
           reg RTL___stage1_f_reset_rsps___deqerror , RTL___stage1_f_reset_rsps___enqerror ; 
             RTL___stage1_f_reset_rsps___deqerror  =0; 
             RTL___stage1_f_reset_rsps___enqerror  =0;
             if ( RTL___stage1_f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___stage1_f_reset_rsps___empty_reg && RTL___stage1_f_reset_rsps___DEQ )
                         begin  
                             RTL___stage1_f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage1_f_reset_rsps___full_reg && RTL___stage1_f_reset_rsps___ENQ &&(! RTL___stage1_f_reset_rsps___DEQ || RTL___stage1_f_reset_rsps___guarded ))
                         begin  
                             RTL___stage1_f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___full_reg ; 
  assign  RTL___stage1_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___empty_reg ;
    reg RTL___stage2_f_reset_reqs___empty_reg ; 
    reg RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___FULL_N = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___EMPTY_N = RTL___stage2_f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___stage2_f_reset_reqs___CLK )
         begin 
             if ( RTL___stage2_f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___stage2_f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___stage2_f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage2_f_reset_reqs___CLR )
                         begin  
                             RTL___stage2_f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___stage2_f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage2_f_reset_reqs___ENQ &&! RTL___stage2_f_reset_reqs___DEQ )
                             begin  
                                 RTL___stage2_f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___stage2_f_reset_reqs___full_reg  <=! RTL___stage2_f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage2_f_reset_reqs___ENQ && RTL___stage2_f_reset_reqs___DEQ )
                                 begin  
                                     RTL___stage2_f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___stage2_f_reset_reqs___empty_reg  <=! RTL___stage2_f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage2_f_reset_reqs___CLK )
         begin : RTL___stage2_f_reset_reqs___error_checks 
           reg RTL___stage2_f_reset_reqs___deqerror , RTL___stage2_f_reset_reqs___enqerror ; 
             RTL___stage2_f_reset_reqs___deqerror  =0; 
             RTL___stage2_f_reset_reqs___enqerror  =0;
             if ( RTL___stage2_f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___stage2_f_reset_reqs___empty_reg && RTL___stage2_f_reset_reqs___DEQ )
                         begin  
                             RTL___stage2_f_reset_reqs___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage2_f_reset_reqs___full_reg && RTL___stage2_f_reset_reqs___ENQ &&(! RTL___stage2_f_reset_reqs___DEQ || RTL___stage2_f_reset_reqs___guarded ))
                         begin  
                             RTL___stage2_f_reset_reqs___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_reqs___full_reg ; 
  assign  RTL___stage2_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_reqs___empty_reg ;
    reg RTL___stage2_f_reset_rsps___empty_reg ; 
    reg RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___FULL_N = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___EMPTY_N = RTL___stage2_f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___stage2_f_reset_rsps___CLK )
         begin 
             if ( RTL___stage2_f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___stage2_f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___stage2_f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage2_f_reset_rsps___CLR )
                         begin  
                             RTL___stage2_f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___stage2_f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage2_f_reset_rsps___ENQ &&! RTL___stage2_f_reset_rsps___DEQ )
                             begin  
                                 RTL___stage2_f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___stage2_f_reset_rsps___full_reg  <=! RTL___stage2_f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage2_f_reset_rsps___ENQ && RTL___stage2_f_reset_rsps___DEQ )
                                 begin  
                                     RTL___stage2_f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___stage2_f_reset_rsps___empty_reg  <=! RTL___stage2_f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage2_f_reset_rsps___CLK )
         begin : RTL___stage2_f_reset_rsps___error_checks 
           reg RTL___stage2_f_reset_rsps___deqerror , RTL___stage2_f_reset_rsps___enqerror ; 
             RTL___stage2_f_reset_rsps___deqerror  =0; 
             RTL___stage2_f_reset_rsps___enqerror  =0;
             if ( RTL___stage2_f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___stage2_f_reset_rsps___empty_reg && RTL___stage2_f_reset_rsps___DEQ )
                         begin  
                             RTL___stage2_f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage2_f_reset_rsps___full_reg && RTL___stage2_f_reset_rsps___ENQ &&(! RTL___stage2_f_reset_rsps___DEQ || RTL___stage2_f_reset_rsps___guarded ))
                         begin  
                             RTL___stage2_f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___full_reg ; 
  assign  RTL___stage2_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___empty_reg ;
    reg RTL___stage3_f_reset_reqs___empty_reg ; 
    reg RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___FULL_N = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___EMPTY_N = RTL___stage3_f_reset_reqs___empty_reg ; 
  always @( posedge  RTL___stage3_f_reset_reqs___CLK )
         begin 
             if ( RTL___stage3_f_reset_reqs___RST ==1'b0)
                 begin  
                     RTL___stage3_f_reset_reqs___empty_reg  <=1'b0; 
                     RTL___stage3_f_reset_reqs___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage3_f_reset_reqs___CLR )
                         begin  
                             RTL___stage3_f_reset_reqs___empty_reg  <=1'b0; 
                             RTL___stage3_f_reset_reqs___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage3_f_reset_reqs___ENQ &&! RTL___stage3_f_reset_reqs___DEQ )
                             begin  
                                 RTL___stage3_f_reset_reqs___empty_reg  <=1'b1; 
                                 RTL___stage3_f_reset_reqs___full_reg  <=! RTL___stage3_f_reset_reqs___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage3_f_reset_reqs___ENQ && RTL___stage3_f_reset_reqs___DEQ )
                                 begin  
                                     RTL___stage3_f_reset_reqs___full_reg  <=1'b1; 
                                     RTL___stage3_f_reset_reqs___empty_reg  <=! RTL___stage3_f_reset_reqs___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage3_f_reset_reqs___CLK )
         begin : RTL___stage3_f_reset_reqs___error_checks 
           reg RTL___stage3_f_reset_reqs___deqerror , RTL___stage3_f_reset_reqs___enqerror ; 
             RTL___stage3_f_reset_reqs___deqerror  =0; 
             RTL___stage3_f_reset_reqs___enqerror  =0;
             if ( RTL___stage3_f_reset_reqs___RST ==!1'b0)
                 begin 
                     if (! RTL___stage3_f_reset_reqs___empty_reg && RTL___stage3_f_reset_reqs___DEQ )
                         begin  
                             RTL___stage3_f_reset_reqs___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage3_f_reset_reqs___full_reg && RTL___stage3_f_reset_reqs___ENQ &&(! RTL___stage3_f_reset_reqs___DEQ || RTL___stage3_f_reset_reqs___guarded ))
                         begin  
                             RTL___stage3_f_reset_reqs___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_reqs___full_reg ; 
  assign  RTL___stage3_f_reset_reqs___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_reqs___empty_reg ;
    reg RTL___stage3_f_reset_rsps___empty_reg ; 
    reg RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___FULL_N = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___EMPTY_N = RTL___stage3_f_reset_rsps___empty_reg ; 
  always @( posedge  RTL___stage3_f_reset_rsps___CLK )
         begin 
             if ( RTL___stage3_f_reset_rsps___RST ==1'b0)
                 begin  
                     RTL___stage3_f_reset_rsps___empty_reg  <=1'b0; 
                     RTL___stage3_f_reset_rsps___full_reg  <=1'b1;
                 end 
              else 
                 begin 
                     if ( RTL___stage3_f_reset_rsps___CLR )
                         begin  
                             RTL___stage3_f_reset_rsps___empty_reg  <=1'b0; 
                             RTL___stage3_f_reset_rsps___full_reg  <=1'b1;
                         end 
                      else 
                         if ( RTL___stage3_f_reset_rsps___ENQ &&! RTL___stage3_f_reset_rsps___DEQ )
                             begin  
                                 RTL___stage3_f_reset_rsps___empty_reg  <=1'b1; 
                                 RTL___stage3_f_reset_rsps___full_reg  <=! RTL___stage3_f_reset_rsps___empty_reg ;
                             end 
                          else 
                             if (! RTL___stage3_f_reset_rsps___ENQ && RTL___stage3_f_reset_rsps___DEQ )
                                 begin  
                                     RTL___stage3_f_reset_rsps___full_reg  <=1'b1; 
                                     RTL___stage3_f_reset_rsps___empty_reg  <=! RTL___stage3_f_reset_rsps___full_reg ;
                                 end 
                 end 
         end
  always @( posedge  RTL___stage3_f_reset_rsps___CLK )
         begin : RTL___stage3_f_reset_rsps___error_checks 
           reg RTL___stage3_f_reset_rsps___deqerror , RTL___stage3_f_reset_rsps___enqerror ; 
             RTL___stage3_f_reset_rsps___deqerror  =0; 
             RTL___stage3_f_reset_rsps___enqerror  =0;
             if ( RTL___stage3_f_reset_rsps___RST ==!1'b0)
                 begin 
                     if (! RTL___stage3_f_reset_rsps___empty_reg && RTL___stage3_f_reset_rsps___DEQ )
                         begin  
                             RTL___stage3_f_reset_rsps___deqerror  =1;$display("Warning: FIFO20: %m -- Dequeuing from empty fifo");
                         end 
                     if (! RTL___stage3_f_reset_rsps___full_reg && RTL___stage3_f_reset_rsps___ENQ &&(! RTL___stage3_f_reset_rsps___DEQ || RTL___stage3_f_reset_rsps___guarded ))
                         begin  
                             RTL___stage3_f_reset_rsps___enqerror  =1;$display("Warning: FIFO20: %m -- Enqueuing to a full fifo");
                         end 
                 end 
         end
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___full_reg ; 
  assign  RTL___stage3_f_reset_rsps___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___empty_reg ;
    assign RTL___csr_regfile___f_reset_rsps___RST = RTL___csr_regfile___RST_N;
    assign RTL___csr_regfile___f_reset_rsps___CLK = RTL___csr_regfile___CLK;
    assign RTL___csr_regfile___f_reset_rsps___ENQ = RTL___csr_regfile___f_reset_rsps$ENQ;
    assign RTL___csr_regfile___f_reset_rsps___CLR = RTL___csr_regfile___f_reset_rsps$CLR;
    assign RTL___csr_regfile___f_reset_rsps___DEQ = RTL___csr_regfile___f_reset_rsps$DEQ;
    assign RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL___csr_regfile___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___csr_regfile___f_reset_rsps___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL___csr_regfile___f_reset_rsps$FULL_N = RTL___csr_regfile___f_reset_rsps___FULL_N;
    assign RTL___csr_regfile___f_reset_rsps$EMPTY_N = RTL___csr_regfile___f_reset_rsps___EMPTY_N;
    assign RTL___stage1_f_reset_reqs___RST = RTL___RST_N;
    assign RTL___stage1_f_reset_reqs___CLK = RTL___CLK;
    assign RTL___stage1_f_reset_reqs___ENQ = RTL___stage1_f_reset_reqs$ENQ;
    assign RTL___stage1_f_reset_reqs___CLR = RTL___stage1_f_reset_reqs$CLR;
    assign RTL___stage1_f_reset_reqs___DEQ = RTL___stage1_f_reset_reqs$DEQ;
    assign RTL___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___stage1_f_reset_reqs___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL___stage1_f_reset_reqs$FULL_N = RTL___stage1_f_reset_reqs___FULL_N;
    assign RTL___stage1_f_reset_reqs$EMPTY_N = RTL___stage1_f_reset_reqs___EMPTY_N;
    assign RTL___stage1_f_reset_rsps___RST = RTL___RST_N;
    assign RTL___stage1_f_reset_rsps___CLK = RTL___CLK;
    assign RTL___stage1_f_reset_rsps___ENQ = RTL___stage1_f_reset_rsps$ENQ;
    assign RTL___stage1_f_reset_rsps___CLR = RTL___stage1_f_reset_rsps$CLR;
    assign RTL___stage1_f_reset_rsps___DEQ = RTL___stage1_f_reset_rsps$DEQ;
    assign RTL___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___stage1_f_reset_rsps___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL___stage1_f_reset_rsps$FULL_N = RTL___stage1_f_reset_rsps___FULL_N;
    assign RTL___stage1_f_reset_rsps$EMPTY_N = RTL___stage1_f_reset_rsps___EMPTY_N;
    assign RTL___stage2_f_reset_reqs___RST = RTL___RST_N;
    assign RTL___stage2_f_reset_reqs___CLK = RTL___CLK;
    assign RTL___stage2_f_reset_reqs___ENQ = RTL___stage2_f_reset_reqs$ENQ;
    assign RTL___stage2_f_reset_reqs___CLR = RTL___stage2_f_reset_reqs$CLR;
    assign RTL___stage2_f_reset_reqs___DEQ = RTL___stage2_f_reset_reqs$DEQ;
    assign RTL___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    assign RTL___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___stage2_f_reset_reqs___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    assign RTL___stage2_f_reset_reqs$FULL_N = RTL___stage2_f_reset_reqs___FULL_N;
    assign RTL___stage2_f_reset_reqs$EMPTY_N = RTL___stage2_f_reset_reqs___EMPTY_N;
    assign RTL___stage2_f_reset_rsps___RST = RTL___RST_N;
    assign RTL___stage2_f_reset_rsps___CLK = RTL___CLK;
    assign RTL___stage2_f_reset_rsps___ENQ = RTL___stage2_f_reset_rsps$ENQ;
    assign RTL___stage2_f_reset_rsps___CLR = RTL___stage2_f_reset_rsps$CLR;
    assign RTL___stage2_f_reset_rsps___DEQ = RTL___stage2_f_reset_rsps$DEQ;
    assign RTL___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    assign RTL___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___stage2_f_reset_rsps___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    assign RTL___stage2_f_reset_rsps$FULL_N = RTL___stage2_f_reset_rsps___FULL_N;
    assign RTL___stage2_f_reset_rsps$EMPTY_N = RTL___stage2_f_reset_rsps___EMPTY_N;
    assign RTL___stage3_f_reset_reqs___RST = RTL___RST_N;
    assign RTL___stage3_f_reset_reqs___CLK = RTL___CLK;
    assign RTL___stage3_f_reset_reqs___ENQ = RTL___stage3_f_reset_reqs$ENQ;
    assign RTL___stage3_f_reset_reqs___CLR = RTL___stage3_f_reset_reqs$CLR;
    assign RTL___stage3_f_reset_reqs___DEQ = RTL___stage3_f_reset_reqs$DEQ;
    assign RTL___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___stage3_f_reset_reqs___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    assign RTL___stage3_f_reset_reqs$FULL_N = RTL___stage3_f_reset_reqs___FULL_N;
    assign RTL___stage3_f_reset_reqs$EMPTY_N = RTL___stage3_f_reset_reqs___EMPTY_N;
    assign RTL___stage3_f_reset_rsps___RST = RTL___RST_N;
    assign RTL___stage3_f_reset_rsps___CLK = RTL___CLK;
    assign RTL___stage3_f_reset_rsps___ENQ = RTL___stage3_f_reset_rsps$ENQ;
    assign RTL___stage3_f_reset_rsps___CLR = RTL___stage3_f_reset_rsps$CLR;
    assign RTL___stage3_f_reset_rsps___DEQ = RTL___stage3_f_reset_rsps$DEQ;
    assign RTL___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    assign RTL___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___stage3_f_reset_rsps___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    assign RTL___stage3_f_reset_rsps$FULL_N = RTL___stage3_f_reset_rsps___FULL_N;
    assign RTL___stage3_f_reset_rsps$EMPTY_N = RTL___stage3_f_reset_rsps___EMPTY_N;
     
  assign  RTL___CAN_FIRE_RL_rl_show_pipe = RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL___rg_state !=4'd0&& RTL___rg_state !=4'd1&& RTL___rg_state !=4'd12; 
  assign  RTL___WILL_FIRE_RL_rl_show_pipe = RTL___CAN_FIRE_RL_rl_show_pipe ; 
  assign  RTL___CAN_FIRE_RL_rl_reset_complete = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___WILL_FIRE_RL_rl_reset_complete = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___CAN_FIRE_RL_rl_pipe = RTL___rg_state ==4'd3&&( RTL___stage3_rg_full || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0|| RTL___stage1_rg_full )&&( RTL___stage3_rg_full || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)&&( RTL___stage3_rg_full || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0||! RTL___stage1_rg_full || RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 )&&( RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0|| RTL___stage3_rg_full ); 
  assign  RTL___WILL_FIRE_RL_rl_pipe = RTL___CAN_FIRE_RL_rl_pipe ; 
  assign  RTL___CAN_FIRE_RL_rl_stage2_nonpipe = RTL___rg_state ==4'd3&&! RTL___stage3_rg_full && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3; 
  assign  RTL___WILL_FIRE_RL_rl_stage2_nonpipe = RTL___CAN_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_trap = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd11; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_trap = RTL___CAN_FIRE_RL_rl_stage1_trap ; 
  assign  RTL___CAN_FIRE_RL_rl_trap = RTL___rg_state ==4'd4&&(! RTL___stage1_rg_full || RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 ); 
  assign  RTL___WILL_FIRE_RL_rl_trap = RTL___CAN_FIRE_RL_rl_trap ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_CSRR_W = RTL___MUX_rg_state$write_1__SEL_9 ; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_CSRR_W = RTL___MUX_rg_state$write_1__SEL_9 ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_CSRR_W_2 = RTL___rg_state ==4'd6; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 = RTL___rg_state ==4'd6; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_CSRR_S_or_C = RTL___MUX_rg_state$write_1__SEL_10 ; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C = RTL___MUX_rg_state$write_1__SEL_10 ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_CSRR_S_or_C_2 = RTL___rg_state ==4'd7; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 = RTL___rg_state ==4'd7; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_restart_after_csrrx = RTL___rg_state ==4'd8; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx = RTL___CAN_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_xRET = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 &&( RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7|| RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8|| RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9); 
  assign  RTL___WILL_FIRE_RL_rl_stage1_xRET = RTL___CAN_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_FENCE_I = RTL___near_mem$RDY_server_fence_i_request_put && RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_FENCE_I = RTL___CAN_FIRE_RL_rl_stage1_FENCE_I ; 
  assign  RTL___CAN_FIRE_RL_rl_finish_FENCE_I = RTL___near_mem$RDY_server_fence_i_response_get && RTL___rg_state ==4'd9; 
  assign  RTL___WILL_FIRE_RL_rl_finish_FENCE_I = RTL___CAN_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_FENCE = RTL___near_mem$RDY_server_fence_request_put && RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_FENCE = RTL___CAN_FIRE_RL_rl_stage1_FENCE ; 
  assign  RTL___CAN_FIRE_RL_rl_finish_FENCE = RTL___near_mem$RDY_server_fence_response_get && RTL___rg_state ==4'd10; 
  assign  RTL___WILL_FIRE_RL_rl_finish_FENCE = RTL___CAN_FIRE_RL_rl_finish_FENCE ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_SFENCE_VMA = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA = RTL___CAN_FIRE_RL_rl_stage1_SFENCE_VMA ; 
  assign  RTL___CAN_FIRE_RL_rl_finish_SFENCE_VMA = RTL___rg_state ==4'd11; 
  assign  RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA = RTL___CAN_FIRE_RL_rl_finish_SFENCE_VMA ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_WFI = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_WFI = RTL___CAN_FIRE_RL_rl_stage1_WFI ; 
  assign  RTL___CAN_FIRE_RL_rl_WFI_resume = RTL___rg_state ==4'd12&& RTL___csr_regfile$wfi_resume ; 
  assign  RTL___WILL_FIRE_RL_rl_WFI_resume = RTL___CAN_FIRE_RL_rl_WFI_resume ; 
  assign  RTL___CAN_FIRE_RL_rl_reset_from_WFI = RTL___rg_state ==4'd12&& RTL___f_reset_reqs$EMPTY_N ; 
  assign  RTL___WILL_FIRE_RL_rl_reset_from_WFI = RTL___MUX_rg_state$write_1__SEL_4 ; 
  assign  RTL___CAN_FIRE_RL_rl_trap_fetch = RTL___rg_state ==4'd5; 
  assign  RTL___WILL_FIRE_RL_rl_trap_fetch = RTL___CAN_FIRE_RL_rl_trap_fetch ; 
  assign  RTL___CAN_FIRE_RL_rl_stage1_interrupt =( RTL___csr_regfile$interrupt_pending [4]|| RTL___csr_regfile$nmi_pending )&& RTL___rg_state ==4'd3&& RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0&&! RTL___stage3_rg_full ; 
  assign  RTL___WILL_FIRE_RL_rl_stage1_interrupt = RTL___CAN_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL___CAN_FIRE_RL_rl_reset_start = RTL___gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 && RTL___rg_state ==4'd0; 
  assign  RTL___WILL_FIRE_RL_rl_reset_start = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___CAN_FIRE_RL_stage3_rl_reset = RTL___stage3_f_reset_reqs$EMPTY_N && RTL___stage3_f_reset_rsps$FULL_N ; 
  assign  RTL___WILL_FIRE_RL_stage3_rl_reset = RTL___CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL___CAN_FIRE_RL_stage2_rl_reset_end = RTL___stage2_f_reset_rsps$FULL_N && RTL___stage2_rg_resetting ; 
  assign  RTL___WILL_FIRE_RL_stage2_rl_reset_end = RTL___CAN_FIRE_RL_stage2_rl_reset_end ; 
  assign  RTL___CAN_FIRE_RL_stage2_rl_reset_begin = RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___WILL_FIRE_RL_stage2_rl_reset_begin = RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___CAN_FIRE_RL_stage1_rl_reset = RTL___stage1_f_reset_reqs$EMPTY_N && RTL___stage1_f_reset_rsps$FULL_N ; 
  assign  RTL___WILL_FIRE_RL_stage1_rl_reset = RTL___CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL___MUX_csr_regfile$mav_csr_write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 ; 
  assign  RTL___MUX_gpr_regfile$write_rd_1__SEL_3 = RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 ; 
  assign  RTL___MUX_near_mem$imem_req_1__SEL_1 = RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset ; 
  assign  RTL___MUX_near_mem$imem_req_1__SEL_2 = RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 ; 
  assign  RTL___MUX_near_mem$imem_req_1__SEL_5 = RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL___MUX_rg_next_pc$write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_stage1_WFI || RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_stage1_FENCE || RTL___WILL_FIRE_RL_rl_stage1_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W ; 
  assign  RTL___MUX_rg_retiring$write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2; 
  assign  RTL___MUX_rg_state$write_1__SEL_1 = RTL___gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 && RTL___rg_state ==4'd1; 
  assign  RTL___MUX_rg_state$write_1__SEL_4 = RTL___CAN_FIRE_RL_rl_reset_from_WFI &&! RTL___WILL_FIRE_RL_rl_WFI_resume ; 
  assign  RTL___MUX_rg_state$write_1__SEL_6 = RTL___WILL_FIRE_RL_rl_trap_fetch || RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  assign  RTL___MUX_rg_state$write_1__SEL_7 = RTL___WILL_FIRE_RL_rl_stage1_interrupt || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL___MUX_rg_state$write_1__SEL_8 = RTL___WILL_FIRE_RL_rl_stage1_xRET || RTL___WILL_FIRE_RL_rl_trap ; 
  assign  RTL___MUX_rg_state$write_1__SEL_9 = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2; 
  assign  RTL___MUX_rg_state$write_1__SEL_10 = RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3; 
  assign  RTL___MUX_rg_trap_info$write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W ; 
  assign  RTL___MUX_rg_trap_instr$write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_stage1_interrupt || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage1_trap ; 
  assign  RTL___MUX_rg_trap_interrupt$write_1__SEL_1 = RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage2_nonpipe ; 
  always @(     RTL___rg_trap_instr                or   RTL___csr_regfile$read_csr            or   RTL___y__h12191           or   RTL___IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868  )
         begin 
             case ( RTL___rg_trap_instr [14:12])
              3 'b010,3'b110: 
                  RTL___MUX_csr_regfile$mav_csr_write_2__VAL_2  = RTL___IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 ;
              default : 
                  RTL___MUX_csr_regfile$mav_csr_write_2__VAL_2  = RTL___csr_regfile$read_csr [31:0]& RTL___y__h12191 ;endcase
         end
  assign  RTL___MUX_rg_state$write_1__VAL_1 = RTL___rg_run_on_reset  ? 4'd3:4'd2; 
  assign  RTL___MUX_rg_state$write_1__VAL_2 = RTL___csr_regfile$access_permitted_1  ? 4'd8:4'd4; 
  assign  RTL___MUX_rg_state$write_1__VAL_3 = RTL___csr_regfile$access_permitted_2  ? 4'd8:4'd4; 
  assign  RTL___MUX_rg_trap_info$write_1__VAL_1 ={ RTL___near_mem$imem_pc ,4'd2, RTL___value__h6967 }; 
  assign  RTL___MUX_rg_trap_info$write_1__VAL_2 ={ RTL___stage2_rg_stage2 [166:135], RTL___near_mem$dmem_exc_code , RTL___stage2_rg_stage2 [95:64]}; 
  assign  RTL___MUX_rg_trap_info$write_1__VAL_3 ={ RTL___near_mem$imem_pc , RTL___IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 }; 
  assign  RTL___MUX_rg_trap_info$write_1__VAL_4 ={ RTL___near_mem$imem_pc , RTL___x_exc_code__h15410 ,32'd0}; 
  assign  RTL___MUX_s1_to_s2$write_1__VAL_1 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL___MUX_stage1_rg_full$write_1__VAL_10 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 ||( RTL___csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 || RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 )&& RTL___stage1_rg_full ; 
  assign  RTL___MUX_stage2_rg_full$write_1__VAL_3 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd2&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0; 
  assign  RTL___cfg_logdelay$D_IN = RTL___set_verbosity_logdelay ; 
  assign  RTL___cfg_logdelay$EN = RTL___EN_set_verbosity ; 
  assign  RTL___cfg_verbosity$D_IN = RTL___set_verbosity_verbosity ; 
  assign  RTL___cfg_verbosity$EN = RTL___EN_set_verbosity ; 
  assign  RTL___rg_csr_pc$D_IN = RTL___near_mem$imem_pc ; 
  assign  RTL___rg_csr_pc$EN = RTL___MUX_rg_trap_info$write_1__SEL_1 ; 
  assign  RTL___rg_csr_val1$D_IN = RTL___x_out_data_to_stage2_val1__h5224 ; 
  assign  RTL___rg_csr_val1$EN = RTL___MUX_rg_trap_info$write_1__SEL_1 ; 
  always @(      RTL___WILL_FIRE_RL_rl_trap                  or   RTL___csr_regfile$csr_trap_actions             or   RTL___WILL_FIRE_RL_rl_stage1_xRET            or   RTL___csr_regfile$csr_ret_actions           or   RTL___WILL_FIRE_RL_rl_reset_start  )
         begin 
             case (1'b1) 
              RTL___WILL_FIRE_RL_rl_trap  : 
                  RTL___rg_cur_priv$D_IN  = RTL___csr_regfile$csr_trap_actions [1:0]; 
              RTL___WILL_FIRE_RL_rl_stage1_xRET  : 
                  RTL___rg_cur_priv$D_IN  = RTL___csr_regfile$csr_ret_actions [33:32]; 
              RTL___WILL_FIRE_RL_rl_reset_start  : 
                  RTL___rg_cur_priv$D_IN  =2'b11;
              default : 
                  RTL___rg_cur_priv$D_IN  =2'b10;endcase
         end
  assign  RTL___rg_cur_priv$EN = RTL___WILL_FIRE_RL_rl_trap || RTL___WILL_FIRE_RL_rl_stage1_xRET || RTL___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___rg_mstatus_MXR$D_IN = RTL___csr_regfile$read_mstatus [19]; 
  assign  RTL___rg_mstatus_MXR$EN = RTL___MUX_rg_state$write_1__SEL_8 ; 
  always @(       RTL___MUX_rg_next_pc$write_1__SEL_1                    or   RTL___x_out_next_pc__h5189              or   RTL___WILL_FIRE_RL_rl_trap             or   RTL___csr_regfile$csr_trap_actions            or   RTL___WILL_FIRE_RL_rl_stage1_xRET           or   RTL___csr_regfile$csr_ret_actions  )
         begin 
             case (1'b1) 
              RTL___MUX_rg_next_pc$write_1__SEL_1  : 
                  RTL___rg_next_pc$D_IN  = RTL___x_out_next_pc__h5189 ; 
              RTL___WILL_FIRE_RL_rl_trap  : 
                  RTL___rg_next_pc$D_IN  = RTL___csr_regfile$csr_trap_actions [97:66]; 
              RTL___WILL_FIRE_RL_rl_stage1_xRET  : 
                  RTL___rg_next_pc$D_IN  = RTL___csr_regfile$csr_ret_actions [65:34];
              default : 
                  RTL___rg_next_pc$D_IN  =32'hAAAAAAAA;endcase
         end
  assign  RTL___rg_next_pc$EN = RTL___WILL_FIRE_RL_rl_stage1_WFI || RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_stage1_FENCE || RTL___WILL_FIRE_RL_rl_stage1_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_trap || RTL___WILL_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL___rg_retiring$D_IN =1'd1; 
  assign  RTL___rg_retiring$EN = RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 || RTL___WILL_FIRE_RL_rl_stage1_WFI || RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_stage1_FENCE || RTL___WILL_FIRE_RL_rl_stage1_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_xRET || RTL___WILL_FIRE_RL_rl_trap || RTL___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___rg_run_on_reset$D_IN = RTL___f_reset_reqs$D_OUT ; 
  assign  RTL___rg_run_on_reset$EN = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___rg_sstatus_SUM$D_IN =1'd0; 
  assign  RTL___rg_sstatus_SUM$EN = RTL___MUX_rg_state$write_1__SEL_8 ; 
  assign  RTL___rg_start_CPI_cycles$D_IN = RTL___csr_regfile$read_csr_mcycle ; 
  assign  RTL___rg_start_CPI_cycles$EN = RTL___MUX_near_mem$imem_req_1__SEL_1 ; 
  assign  RTL___rg_start_CPI_instrs$D_IN = RTL___csr_regfile$read_csr_minstret ; 
  assign  RTL___rg_start_CPI_instrs$EN = RTL___MUX_near_mem$imem_req_1__SEL_1 ; 
  always @(                  RTL___WILL_FIRE_RL_rl_reset_complete                                          or   RTL___MUX_rg_state$write_1__VAL_1                         or   RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2                        or   RTL___MUX_rg_state$write_1__VAL_2                       or   RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2                      or   RTL___MUX_rg_state$write_1__VAL_3                     or   RTL___WILL_FIRE_RL_rl_reset_from_WFI                    or   RTL___WILL_FIRE_RL_rl_reset_start                   or   RTL___MUX_rg_state$write_1__SEL_6                  or   RTL___MUX_rg_state$write_1__SEL_7                 or   RTL___MUX_rg_state$write_1__SEL_8                or   RTL___WILL_FIRE_RL_rl_stage1_CSRR_W               or   RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C              or   RTL___WILL_FIRE_RL_rl_stage1_FENCE_I             or   RTL___WILL_FIRE_RL_rl_stage1_FENCE            or   RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA           or   RTL___WILL_FIRE_RL_rl_stage1_WFI  )
         begin 
             case (1'b1) 
              RTL___WILL_FIRE_RL_rl_reset_complete  : 
                  RTL___rg_state$D_IN  = RTL___MUX_rg_state$write_1__VAL_1 ; 
              RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2  : 
                  RTL___rg_state$D_IN  = RTL___MUX_rg_state$write_1__VAL_2 ; 
              RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2  : 
                  RTL___rg_state$D_IN  = RTL___MUX_rg_state$write_1__VAL_3 ; 
              RTL___WILL_FIRE_RL_rl_reset_from_WFI  : 
                  RTL___rg_state$D_IN  =4'd0; 
              RTL___WILL_FIRE_RL_rl_reset_start  : 
                  RTL___rg_state$D_IN  =4'd1; 
              RTL___MUX_rg_state$write_1__SEL_6  : 
                  RTL___rg_state$D_IN  =4'd3; 
              RTL___MUX_rg_state$write_1__SEL_7  : 
                  RTL___rg_state$D_IN  =4'd4; 
              RTL___MUX_rg_state$write_1__SEL_8  : 
                  RTL___rg_state$D_IN  =4'd5; 
              RTL___WILL_FIRE_RL_rl_stage1_CSRR_W  : 
                  RTL___rg_state$D_IN  =4'd6; 
              RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C  : 
                  RTL___rg_state$D_IN  =4'd7; 
              RTL___WILL_FIRE_RL_rl_stage1_FENCE_I  : 
                  RTL___rg_state$D_IN  =4'd9; 
              RTL___WILL_FIRE_RL_rl_stage1_FENCE  : 
                  RTL___rg_state$D_IN  =4'd10; 
              RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA  : 
                  RTL___rg_state$D_IN  =4'd11; 
              RTL___WILL_FIRE_RL_rl_stage1_WFI  : 
                  RTL___rg_state$D_IN  =4'd12;
              default : 
                  RTL___rg_state$D_IN  =4'b1010;endcase
         end
  assign  RTL___rg_state$EN = RTL___WILL_FIRE_RL_rl_reset_complete || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 || RTL___WILL_FIRE_RL_rl_reset_from_WFI || RTL___WILL_FIRE_RL_rl_reset_start || RTL___WILL_FIRE_RL_rl_trap_fetch || RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL___WILL_FIRE_RL_rl_stage1_interrupt || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage2_nonpipe || RTL___WILL_FIRE_RL_rl_stage1_xRET || RTL___WILL_FIRE_RL_rl_trap || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_FENCE || RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_stage1_WFI ; 
  always @(         RTL___MUX_rg_trap_info$write_1__SEL_1                        or   RTL___MUX_rg_trap_info$write_1__VAL_1                or   RTL___WILL_FIRE_RL_rl_stage2_nonpipe               or   RTL___MUX_rg_trap_info$write_1__VAL_2              or   RTL___WILL_FIRE_RL_rl_stage1_trap             or   RTL___MUX_rg_trap_info$write_1__VAL_3            or   RTL___WILL_FIRE_RL_rl_stage1_interrupt           or   RTL___MUX_rg_trap_info$write_1__VAL_4  )
         begin 
             case (1'b1) 
              RTL___MUX_rg_trap_info$write_1__SEL_1  : 
                  RTL___rg_trap_info$D_IN  = RTL___MUX_rg_trap_info$write_1__VAL_1 ; 
              RTL___WILL_FIRE_RL_rl_stage2_nonpipe  : 
                  RTL___rg_trap_info$D_IN  = RTL___MUX_rg_trap_info$write_1__VAL_2 ; 
              RTL___WILL_FIRE_RL_rl_stage1_trap  : 
                  RTL___rg_trap_info$D_IN  = RTL___MUX_rg_trap_info$write_1__VAL_3 ; 
              RTL___WILL_FIRE_RL_rl_stage1_interrupt  : 
                  RTL___rg_trap_info$D_IN  = RTL___MUX_rg_trap_info$write_1__VAL_4 ;
              default : 
                  RTL___rg_trap_info$D_IN  =68'hAAAAAAAAAAAAAAAAA;endcase
         end
  assign  RTL___rg_trap_info$EN = RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage2_nonpipe || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL___rg_trap_instr$D_IN = RTL___MUX_rg_trap_instr$write_1__SEL_1  ?  RTL___near_mem$imem_instr : RTL___stage2_rg_stage2 [134:103]; 
  assign  RTL___rg_trap_instr$EN = RTL___WILL_FIRE_RL_rl_stage1_interrupt || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage2_nonpipe ; 
  assign  RTL___rg_trap_interrupt$D_IN =! RTL___MUX_rg_trap_interrupt$write_1__SEL_1 ; 
  assign  RTL___rg_trap_interrupt$EN = RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C || RTL___WILL_FIRE_RL_rl_stage1_CSRR_W || RTL___WILL_FIRE_RL_rl_stage1_trap || RTL___WILL_FIRE_RL_rl_stage2_nonpipe || RTL___WILL_FIRE_RL_rl_stage1_interrupt ; 
  assign  RTL___s1_to_s2$D_IN = RTL___WILL_FIRE_RL_rl_pipe && RTL___MUX_s1_to_s2$write_1__VAL_1 ; 
  assign  RTL___s1_to_s2$EN = RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___s2_to_s3$D_IN = RTL___MUX_rg_retiring$write_1__SEL_1 ; 
  assign  RTL___s2_to_s3$EN = RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_rl_reset_start ; 
  assign  RTL___s3_deq$D_IN = RTL___WILL_FIRE_RL_rl_pipe && RTL___stage3_rg_full ; 
  assign  RTL___s3_deq$EN = RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_rl_reset_start ; 
  always @(             RTL___WILL_FIRE_RL_stage1_rl_reset                                or   RTL___WILL_FIRE_RL_rl_trap_fetch                    or   RTL___WILL_FIRE_RL_rl_WFI_resume                   or   RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA                  or   RTL___WILL_FIRE_RL_rl_finish_FENCE                 or   RTL___WILL_FIRE_RL_rl_finish_FENCE_I                or   RTL___WILL_FIRE_RL_rl_stage1_xRET               or   RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx              or   RTL___WILL_FIRE_RL_rl_trap             or   RTL___WILL_FIRE_RL_rl_pipe            or   RTL___MUX_stage1_rg_full$write_1__VAL_10           or   RTL___MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL___WILL_FIRE_RL_stage1_rl_reset  : 
              RTL___stage1_rg_full$D_IN  =1'd0; 
          RTL___WILL_FIRE_RL_rl_trap_fetch  || RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I : 
              RTL___stage1_rg_full$D_IN  =1'd1; 
          RTL___WILL_FIRE_RL_rl_stage1_xRET  : 
              RTL___stage1_rg_full$D_IN  =1'd0; 
          RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx  : 
              RTL___stage1_rg_full$D_IN  =1'd1; 
          RTL___WILL_FIRE_RL_rl_trap  : 
              RTL___stage1_rg_full$D_IN  =1'd0; 
          RTL___WILL_FIRE_RL_rl_pipe  : 
              RTL___stage1_rg_full$D_IN  = RTL___MUX_stage1_rg_full$write_1__VAL_10 ; 
          RTL___MUX_near_mem$imem_req_1__SEL_1  : 
              RTL___stage1_rg_full$D_IN  =1'd1;
          default : 
              RTL___stage1_rg_full$D_IN  =1'b0;endcase
  assign  RTL___stage1_rg_full$EN = RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset || RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_rl_stage1_xRET || RTL___WILL_FIRE_RL_rl_trap || RTL___WILL_FIRE_RL_stage1_rl_reset || RTL___WILL_FIRE_RL_rl_trap_fetch || RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx ; 
  always @(      RTL___stage2_f_reset_reqs$EMPTY_N                  or   RTL___WILL_FIRE_RL_rl_trap             or   RTL___WILL_FIRE_RL_rl_pipe            or   RTL___MUX_stage2_rg_full$write_1__VAL_3           or   RTL___MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL___stage2_f_reset_reqs$EMPTY_N  || RTL___WILL_FIRE_RL_rl_trap : 
              RTL___stage2_rg_full$D_IN  =1'd0; 
          RTL___WILL_FIRE_RL_rl_pipe  : 
              RTL___stage2_rg_full$D_IN  = RTL___MUX_stage2_rg_full$write_1__VAL_3 ; 
          RTL___MUX_near_mem$imem_req_1__SEL_1  : 
              RTL___stage2_rg_full$D_IN  =1'd0;
          default : 
              RTL___stage2_rg_full$D_IN  =1'b0;endcase
  assign  RTL___stage2_rg_full$EN = RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset || RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_rl_trap || RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___stage2_rg_resetting$D_IN = RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___stage2_rg_resetting$EN = RTL___WILL_FIRE_RL_stage2_rl_reset_end || RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___stage2_rg_stage2$D_IN ={ RTL___rg_cur_priv , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 , RTL___x_out_data_to_stage2_rd__h5222 , RTL___x_out_data_to_stage2_addr__h5223 , RTL___x_out_data_to_stage2_val1__h5224 , RTL___x_out_data_to_stage2_val2__h5225 }; 
  assign  RTL___stage2_rg_stage2$EN = RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 ; 
  always @(     RTL___WILL_FIRE_RL_stage3_rl_reset                or   RTL___WILL_FIRE_RL_rl_pipe            or   RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86           or   RTL___MUX_near_mem$imem_req_1__SEL_1  )
         case (1'b1) 
          RTL___WILL_FIRE_RL_stage3_rl_reset  : 
              RTL___stage3_rg_full$D_IN  =1'd0; 
          RTL___WILL_FIRE_RL_rl_pipe  : 
              RTL___stage3_rg_full$D_IN  = RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2; 
          RTL___MUX_near_mem$imem_req_1__SEL_1  : 
              RTL___stage3_rg_full$D_IN  =1'd0;
          default : 
              RTL___stage3_rg_full$D_IN  =1'b0;endcase
  assign  RTL___stage3_rg_full$EN = RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset || RTL___WILL_FIRE_RL_rl_pipe || RTL___WILL_FIRE_RL_stage3_rl_reset ; 
  assign  RTL___stage3_rg_stage3$D_IN ={ RTL___stage2_rg_stage2 [166:103], RTL___stage2_rg_stage2 [168:167], RTL___stage2_rg_stage2 [102:101]==2'd0|| RTL___near_mem$dmem_valid &&! RTL___near_mem$dmem_exc , RTL___x_out_data_to_stage3_rd__h4667 , RTL___x_out_data_to_stage3_rd_val__h4668 }; 
  assign  RTL___stage3_rg_stage3$EN = RTL___MUX_rg_retiring$write_1__SEL_1 ; 
  assign  RTL___csr_regfile$access_permitted_1_csr_addr = RTL___rg_trap_instr [31:20]; 
  assign  RTL___csr_regfile$access_permitted_1_priv = RTL___rg_cur_priv ; 
  assign  RTL___csr_regfile$access_permitted_1_read_not_write =1'd0; 
  assign  RTL___csr_regfile$access_permitted_2_csr_addr = RTL___rg_trap_instr [31:20]; 
  assign  RTL___csr_regfile$access_permitted_2_priv = RTL___rg_cur_priv ; 
  assign  RTL___csr_regfile$access_permitted_2_read_not_write = RTL___rs1_val__h11920 ==32'd0; 
  assign  RTL___csr_regfile$csr_counter_read_fault_csr_addr =12'h0; 
  assign  RTL___csr_regfile$csr_counter_read_fault_priv =2'h0; 
  always @(  RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415  )
         begin 
             case ( RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 )
              4 'd7: 
                  RTL___csr_regfile$csr_ret_actions_from_priv  =2'b11;
              4 'd8: 
                  RTL___csr_regfile$csr_ret_actions_from_priv  =2'b01;
              default : 
                  RTL___csr_regfile$csr_ret_actions_from_priv  =2'b0;endcase
         end
  assign  RTL___csr_regfile$csr_trap_actions_exc_code = RTL___rg_trap_info [35:32]; 
  assign  RTL___csr_regfile$csr_trap_actions_from_priv = RTL___rg_cur_priv ; 
  assign  RTL___csr_regfile$csr_trap_actions_interrupt = RTL___rg_trap_interrupt &&! RTL___csr_regfile$nmi_pending ; 
  assign  RTL___csr_regfile$csr_trap_actions_nmi = RTL___rg_trap_interrupt && RTL___csr_regfile$nmi_pending ; 
  assign  RTL___csr_regfile$csr_trap_actions_pc = RTL___rg_trap_info [67:36]; 
  assign  RTL___csr_regfile$csr_trap_actions_xtval = RTL___rg_trap_info [31:0]; 
  assign  RTL___csr_regfile$interrupt_pending_cur_priv = RTL___rg_cur_priv ; 
  assign  RTL___csr_regfile$m_external_interrupt_req_set_not_clear = RTL___m_external_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile$mav_csr_write_csr_addr = RTL___rg_trap_instr [31:20]; 
  assign  RTL___csr_regfile$mav_csr_write_word = RTL___MUX_csr_regfile$mav_csr_write_1__SEL_1  ?  RTL___rs1_val__h11213 : RTL___MUX_csr_regfile$mav_csr_write_2__VAL_2 ; 
  assign  RTL___csr_regfile$mav_read_csr_csr_addr =12'h0; 
  assign  RTL___csr_regfile$nmi_req_set_not_clear = RTL___nmi_req_set_not_clear ; 
  assign  RTL___csr_regfile$read_csr_csr_addr = RTL___rg_trap_instr [31:20]; 
  assign  RTL___csr_regfile$read_csr_port2_csr_addr =12'h0; 
  assign  RTL___csr_regfile$s_external_interrupt_req_set_not_clear = RTL___s_external_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile$software_interrupt_req_set_not_clear = RTL___software_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile$timer_interrupt_req_set_not_clear = RTL___timer_interrupt_req_set_not_clear ; 
  assign  RTL___csr_regfile$EN_server_reset_request_put = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___csr_regfile$EN_server_reset_response_get = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___csr_regfile$EN_mav_read_csr =1'b0; 
  assign  RTL___csr_regfile$EN_mav_csr_write = RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 && RTL___rg_trap_instr [19:15]!=5'd0; 
  assign  RTL___csr_regfile$EN_csr_trap_actions = RTL___CAN_FIRE_RL_rl_trap ; 
  assign  RTL___csr_regfile$EN_csr_ret_actions = RTL___CAN_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL___csr_regfile$EN_csr_minstret_incr = RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 || RTL___WILL_FIRE_RL_rl_stage1_WFI || RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_stage1_FENCE || RTL___WILL_FIRE_RL_rl_stage1_FENCE_I || RTL___WILL_FIRE_RL_rl_stage1_xRET ; 
  assign  RTL___csr_regfile$EN_debug =1'b0; 
  assign  RTL___f_reset_reqs$D_IN = RTL___hart0_server_reset_request_put ; 
  assign  RTL___f_reset_reqs$ENQ = RTL___EN_hart0_server_reset_request_put ; 
  assign  RTL___f_reset_reqs$DEQ = RTL___gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 && RTL___rg_state ==4'd0; 
  assign  RTL___f_reset_reqs$CLR =1'b0; 
  assign  RTL___f_reset_rsps$D_IN = RTL___rg_run_on_reset ; 
  assign  RTL___f_reset_rsps$ENQ = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___f_reset_rsps$DEQ = RTL___EN_hart0_server_reset_response_get ; 
  assign  RTL___f_reset_rsps$CLR =1'b0; 
  assign  RTL___gpr_regfile$read_rs1_port2_rs1 =5'h0; 
  assign  RTL___gpr_regfile$read_rs1_rs1 = RTL___near_mem$imem_instr [19:15]; 
  assign  RTL___gpr_regfile$read_rs2_rs2 = RTL___near_mem$imem_instr [24:20]; 
  assign  RTL___gpr_regfile$write_rd_rd =( RTL___MUX_csr_regfile$mav_csr_write_1__SEL_1 || RTL___MUX_gpr_regfile$write_rd_1__SEL_3 ) ?  RTL___rg_trap_instr [11:7]: RTL___stage3_rg_stage3 [36:32]; 
  assign  RTL___gpr_regfile$write_rd_rd_val =( RTL___MUX_csr_regfile$mav_csr_write_1__SEL_1 || RTL___MUX_gpr_regfile$write_rd_1__SEL_3 ) ?  RTL___csr_regfile$read_csr [31:0]: RTL___stage3_rg_stage3 [31:0]; 
  assign  RTL___gpr_regfile$EN_server_reset_request_put = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___gpr_regfile$EN_server_reset_response_get = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___gpr_regfile$EN_write_rd = RTL___WILL_FIRE_RL_rl_pipe && RTL___stage3_rg_full && RTL___stage3_rg_stage3 [37]|| RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 || RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 ; 
  assign  RTL___near_mem$dmem_master_arready = RTL___dmem_master_arready ; 
  assign  RTL___near_mem$dmem_master_awready = RTL___dmem_master_awready ; 
  assign  RTL___near_mem$dmem_master_bid = RTL___dmem_master_bid ; 
  assign  RTL___near_mem$dmem_master_bresp = RTL___dmem_master_bresp ; 
  assign  RTL___near_mem$dmem_master_bvalid = RTL___dmem_master_bvalid ; 
  assign  RTL___near_mem$dmem_master_rdata = RTL___dmem_master_rdata ; 
  assign  RTL___near_mem$dmem_master_rid = RTL___dmem_master_rid ; 
  assign  RTL___near_mem$dmem_master_rlast = RTL___dmem_master_rlast ; 
  assign  RTL___near_mem$dmem_master_rresp = RTL___dmem_master_rresp ; 
  assign  RTL___near_mem$dmem_master_rvalid = RTL___dmem_master_rvalid ; 
  assign  RTL___near_mem$dmem_master_wready = RTL___dmem_master_wready ; 
  assign  RTL___near_mem$dmem_req_addr = RTL___x_out_data_to_stage2_addr__h5223 ; 
  assign  RTL___near_mem$dmem_req_f3 = RTL___near_mem$imem_instr [14:12]; 
  assign  RTL___near_mem$dmem_req_mstatus_MXR = RTL___csr_regfile$read_mstatus [19]; 
  assign  RTL___near_mem$dmem_req_op = RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1; 
  assign  RTL___near_mem$dmem_req_priv = RTL___csr_regfile$read_mstatus [17] ?  RTL___csr_regfile$read_mstatus [12:11]: RTL___rg_cur_priv ; 
  assign  RTL___near_mem$dmem_req_satp = RTL___csr_regfile$read_satp ; 
  assign  RTL___near_mem$dmem_req_sstatus_SUM =1'd0; 
  assign  RTL___near_mem$dmem_req_store_value ={32'd0, RTL___x_out_data_to_stage2_val2__h5225 }; 
  assign  RTL___near_mem$imem_master_arready = RTL___imem_master_arready ; 
  assign  RTL___near_mem$imem_master_awready = RTL___imem_master_awready ; 
  assign  RTL___near_mem$imem_master_bid = RTL___imem_master_bid ; 
  assign  RTL___near_mem$imem_master_bresp = RTL___imem_master_bresp ; 
  assign  RTL___near_mem$imem_master_bvalid = RTL___imem_master_bvalid ; 
  assign  RTL___near_mem$imem_master_rdata = RTL___imem_master_rdata ; 
  assign  RTL___near_mem$imem_master_rid = RTL___imem_master_rid ; 
  assign  RTL___near_mem$imem_master_rlast = RTL___imem_master_rlast ; 
  assign  RTL___near_mem$imem_master_rresp = RTL___imem_master_rresp ; 
  assign  RTL___near_mem$imem_master_rvalid = RTL___imem_master_rvalid ; 
  assign  RTL___near_mem$imem_master_wready = RTL___imem_master_wready ; 
  always @(         RTL___MUX_near_mem$imem_req_1__SEL_1                        or   RTL___soc_map$m_pc_reset_value                or   RTL___WILL_FIRE_RL_rl_trap_fetch               or   RTL___MUX_near_mem$imem_req_1__SEL_5              or   RTL___rg_next_pc             or   RTL___MUX_near_mem$imem_req_1__SEL_2            or   RTL___x_out_next_pc__h5189           or   RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx  )
         begin 
             case (1'b1) 
              RTL___MUX_near_mem$imem_req_1__SEL_1  : 
                  RTL___near_mem$imem_req_addr  = RTL___soc_map$m_pc_reset_value [31:0]; 
              RTL___WILL_FIRE_RL_rl_trap_fetch  || RTL___MUX_near_mem$imem_req_1__SEL_5 : 
                  RTL___near_mem$imem_req_addr  = RTL___rg_next_pc ; 
              RTL___MUX_near_mem$imem_req_1__SEL_2  : 
                  RTL___near_mem$imem_req_addr  = RTL___x_out_next_pc__h5189 ; 
              RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx  : 
                  RTL___near_mem$imem_req_addr  = RTL___x_out_next_pc__h5189 ;
              default : 
                  RTL___near_mem$imem_req_addr  =32'hAAAAAAAA;endcase
         end
  assign  RTL___near_mem$imem_req_f3 =3'b010; 
  assign  RTL___near_mem$imem_req_mstatus_MXR =( RTL___MUX_near_mem$imem_req_1__SEL_1 || RTL___MUX_near_mem$imem_req_1__SEL_2 || RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL___MUX_near_mem$imem_req_1__SEL_5 ) ?  RTL___csr_regfile$read_mstatus [19]: RTL___rg_mstatus_MXR ; 
  assign  RTL___near_mem$imem_req_priv = RTL___rg_cur_priv ; 
  assign  RTL___near_mem$imem_req_satp = RTL___csr_regfile$read_satp ; 
  assign  RTL___near_mem$imem_req_sstatus_SUM = RTL___WILL_FIRE_RL_rl_trap_fetch && RTL___rg_sstatus_SUM ; 
  assign  RTL___near_mem$server_fence_request_put =8'b10101010; 
  assign  RTL___near_mem$EN_server_reset_request_put = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___near_mem$EN_server_reset_response_get = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___near_mem$EN_imem_req = RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset || RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 || RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx || RTL___WILL_FIRE_RL_rl_trap_fetch || RTL___WILL_FIRE_RL_rl_WFI_resume || RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA || RTL___WILL_FIRE_RL_rl_finish_FENCE || RTL___WILL_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL___near_mem$EN_dmem_req = RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 &&( RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1|| RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd2); 
  assign  RTL___near_mem$EN_server_fence_i_request_put = RTL___CAN_FIRE_RL_rl_stage1_FENCE_I ; 
  assign  RTL___near_mem$EN_server_fence_i_response_get = RTL___CAN_FIRE_RL_rl_finish_FENCE_I ; 
  assign  RTL___near_mem$EN_server_fence_request_put = RTL___CAN_FIRE_RL_rl_stage1_FENCE ; 
  assign  RTL___near_mem$EN_server_fence_response_get = RTL___CAN_FIRE_RL_rl_finish_FENCE ; 
  assign  RTL___near_mem$EN_sfence_vma = RTL___CAN_FIRE_RL_rl_stage1_SFENCE_VMA ; 
  assign  RTL___soc_map$m_is_IO_addr_addr =64'h0; 
  assign  RTL___soc_map$m_is_mem_addr_addr =64'h0; 
  assign  RTL___soc_map$m_is_near_mem_IO_addr_addr =64'h0; 
  assign  RTL___stage1_f_reset_reqs$ENQ = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___stage1_f_reset_reqs$DEQ = RTL___CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL___stage1_f_reset_reqs$CLR =1'b0; 
  assign  RTL___stage1_f_reset_rsps$ENQ = RTL___CAN_FIRE_RL_stage1_rl_reset ; 
  assign  RTL___stage1_f_reset_rsps$DEQ = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___stage1_f_reset_rsps$CLR =1'b0; 
  assign  RTL___stage2_f_reset_reqs$ENQ = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___stage2_f_reset_reqs$DEQ = RTL___stage2_f_reset_reqs$EMPTY_N ; 
  assign  RTL___stage2_f_reset_reqs$CLR =1'b0; 
  assign  RTL___stage2_f_reset_rsps$ENQ = RTL___CAN_FIRE_RL_stage2_rl_reset_end ; 
  assign  RTL___stage2_f_reset_rsps$DEQ = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___stage2_f_reset_rsps$CLR =1'b0; 
  assign  RTL___stage3_f_reset_reqs$ENQ = RTL___CAN_FIRE_RL_rl_reset_start ; 
  assign  RTL___stage3_f_reset_reqs$DEQ = RTL___CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL___stage3_f_reset_reqs$CLR =1'b0; 
  assign  RTL___stage3_f_reset_rsps$ENQ = RTL___CAN_FIRE_RL_stage3_rl_reset ; 
  assign  RTL___stage3_f_reset_rsps$DEQ = RTL___MUX_rg_state$write_1__SEL_1 ; 
  assign  RTL___stage3_f_reset_rsps$CLR =1'b0; 
  assign  RTL___IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 =(( RTL___near_mem$imem_instr [6:0]==7'b1100011) ?  RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 : RTL___near_mem$imem_instr [6:0]==7'b1101111|| RTL___near_mem$imem_instr [6:0]==7'b1100111) ?  RTL___data_to_stage2_addr__h5215 :(( RTL___near_mem$imem_instr [6:0]==7'b1110011&& RTL___near_mem$imem_instr [14:12]==3'b0&& RTL___near_mem$imem_instr [11:7]==5'd0&& RTL___near_mem$imem_instr [19:15]==5'd0&& RTL___near_mem$imem_instr [31:20]==12'b000000000001) ?  RTL___near_mem$imem_pc :32'd0); 
  assign  RTL___IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 = RTL___NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252  ? 4'd11:4'd0; 
  assign  RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 = RTL___near_mem$imem_exc  ? 4'd11: RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413 ; 
  assign  RTL___IF_csr_regfile_read_csr_rg_trap_instr_15_BITS__ETC___d868 = RTL___csr_regfile$read_csr [31:0]| RTL___rs1_val__h11920 ; 
  assign  RTL___IF_near_mem_imem_exc__78_THEN_near_mem_imem_ex_ETC___d799 = RTL___near_mem$imem_exc  ? { RTL___near_mem$imem_exc_code , RTL___near_mem$imem_tval }:{ RTL___alu_outputs_exc_code__h5862 , RTL___trap_info_tval__h6925 }; 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 = RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 && RTL___alu_outputs___1_val2__h5367 [1]|| RTL___near_mem$imem_instr [14:12]!=3'b0&& RTL___near_mem$imem_instr [14:12]!=3'b001&& RTL___near_mem$imem_instr [14:12]!=3'b100&& RTL___near_mem$imem_instr [14:12]!=3'b101&& RTL___near_mem$imem_instr [14:12]!=3'b110&& RTL___near_mem$imem_instr [14:12]!=3'b111; 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 = RTL___rs1_val_bypassed__h3337 == RTL___rs2_val__h5339 ; 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 =( RTL___rs1_val_bypassed__h3337 ^32'h80000000)<( RTL___rs2_val__h5339 ^32'h80000000); 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 = RTL___rs1_val_bypassed__h3337 < RTL___rs2_val__h5339 ; 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 =( RTL___near_mem$imem_instr [6:0]==7'b1100011) ?  RTL___near_mem$imem_instr [14:12]!=3'b0&& RTL___near_mem$imem_instr [14:12]!=3'b001&& RTL___near_mem$imem_instr [14:12]!=3'b100&& RTL___near_mem$imem_instr [14:12]!=3'b101&& RTL___near_mem$imem_instr [14:12]!=3'b110&& RTL___near_mem$imem_instr [14:12]!=3'b111|| RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 :((( RTL___near_mem$imem_instr [6:0]==7'b0010011|| RTL___near_mem$imem_instr [6:0]==7'b0110011)&&( RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b101)) ?  RTL___near_mem$imem_instr [25]: RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8 ); 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 =( RTL___near_mem$imem_instr [6:0]==7'b1100011) ? ( RTL___near_mem$imem_instr [14:12]==3'b0|| RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b100|| RTL___near_mem$imem_instr [14:12]==3'b101|| RTL___near_mem$imem_instr [14:12]==3'b110|| RTL___near_mem$imem_instr [14:12]==3'b111)&& RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 :((( RTL___near_mem$imem_instr [6:0]==7'b0010011|| RTL___near_mem$imem_instr [6:0]==7'b0110011)&&( RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b101)) ? ! RTL___near_mem$imem_instr [25]: RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9 ); 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 =(( RTL___near_mem$imem_instr [6:0]==7'b0010011|| RTL___near_mem$imem_instr [6:0]==7'b0110011)&&( RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b101)) ?  RTL___alu_outputs___1_val1__h5480 : RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570 ; 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649 =( RTL___near_mem$imem_instr [6:0]==7'b1100011) ?  RTL___near_mem$imem_instr [14:12]!=3'b0&& RTL___near_mem$imem_instr [14:12]!=3'b001&& RTL___near_mem$imem_instr [14:12]!=3'b100&& RTL___near_mem$imem_instr [14:12]!=3'b101&& RTL___near_mem$imem_instr [14:12]!=3'b110&& RTL___near_mem$imem_instr [14:12]!=3'b111|| RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ||! RTL___alu_outputs___1_val2__h5367 [1]: RTL___near_mem$imem_instr [6:0]!=7'b1101111&& RTL___near_mem$imem_instr [6:0]!=7'b1100111&&( RTL___near_mem$imem_instr [6:0]!=7'b1110011|| RTL___near_mem$imem_instr [14:12]!=3'b0|| RTL___near_mem$imem_instr [11:7]!=5'd0|| RTL___near_mem$imem_instr [19:15]!=5'd0|| RTL___near_mem$imem_instr [31:20]!=12'b0&& RTL___near_mem$imem_instr [31:20]!=12'b000000000001); 
  assign  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d910 = RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 || RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL___IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 =(( RTL___rg_cur_priv ==2'b11|| RTL___rg_cur_priv ==2'b01&&! RTL___csr_regfile$read_mstatus [22])&& RTL___near_mem$imem_instr [31:20]==12'b000100000010) ? 4'd8:( RTL___rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392  ? 4'd10:4'd11); 
  assign  RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 = RTL___stage2_rg_full  ?  RTL___CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5 :2'd0; 
  assign  RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 = RTL___stage2_rg_stage2 [100:96]== RTL___near_mem$imem_instr [19:15]; 
  assign  RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 = RTL___stage2_rg_stage2 [100:96]== RTL___near_mem$imem_instr [24:20]; 
  assign  RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 = RTL___stage2_rg_full  ?  RTL___IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 :2'd0; 
  assign  RTL___IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 =( RTL___stage2_rg_stage2 [100:96]==5'd0) ? 2'd0:(( RTL___near_mem$dmem_valid &&! RTL___near_mem$dmem_exc ) ? 2'd2:2'd1); 
  assign  RTL___IF_stage2_rg_stage2_4_BITS_102_TO_101_5_EQ_0_6_ETC___d85 =( RTL___stage2_rg_stage2 [102:101]==2'd0) ? 2'd2:( RTL___near_mem$dmem_valid  ? ( RTL___near_mem$dmem_exc  ? 2'd3:2'd2):2'd1); 
  assign  RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 = RTL___cur_verbosity__h1827 >4'd1; 
  assign  RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 = RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 &&( RTL___stage2_rg_stage2 [102:101]==2'd0|| RTL___near_mem$dmem_valid &&! RTL___near_mem$dmem_exc ); 
  assign  RTL___NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 = RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3&&( RTL___stage2_rg_stage2 [102:101]==2'd0|| RTL___near_mem$dmem_valid &&! RTL___near_mem$dmem_exc ); 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 =! RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending ||(! RTL___stage1_rg_full || RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 )&&(! RTL___stage1_rg_full || RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 ); 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 =! RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending || RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 &&( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)&& RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d734 &&( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)&& RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ||! RTL___stage1_rg_full ; 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d769 =(! RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending || RTL____0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 )&& RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ; 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 =(! RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending || RTL____0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 )&&( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2|| RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0); 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d776 = RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 &&( RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d773 && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 ||! RTL___stage1_rg_full ); 
  assign  RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 =! RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending ||! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL___NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 =! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd0&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd1&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd2&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd3&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd4&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd5&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd6&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd7&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd8&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd9&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd10; 
  assign  RTL___NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 =( RTL___near_mem$imem_instr [14:12]!=3'b0|| RTL___near_mem$imem_instr [6:0]==7'b0110011&& RTL___near_mem$imem_instr [30])&&( RTL___near_mem$imem_instr [14:12]!=3'b0|| RTL___near_mem$imem_instr [6:0]!=7'b0110011||! RTL___near_mem$imem_instr [30])&& RTL___near_mem$imem_instr [14:12]!=3'b010&& RTL___near_mem$imem_instr [14:12]!=3'b011&& RTL___near_mem$imem_instr [14:12]!=3'b100&& RTL___near_mem$imem_instr [14:12]!=3'b110&& RTL___near_mem$imem_instr [14:12]!=3'b111; 
  assign  RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 =! RTL___near_mem$imem_valid || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd1&&( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 || RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ); 
  assign  RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d702 = RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 ||! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d713 = RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 || RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL___SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 ={{20{ RTL___near_memimem_instr_BITS_31_TO_20__q7 [11]}}, RTL___near_memimem_instr_BITS_31_TO_20__q7 }; 
  assign  RTL____0_OR_0_OR_near_mem_imem_exc__78_OR_IF_near_mem_ETC___d767 = RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ; 
  assign  RTL____theResult_____1_fst__h6562 =( RTL___near_mem$imem_instr [14:12]==3'b0&& RTL___near_mem$imem_instr [6:0]==7'b0110011&& RTL___near_mem$imem_instr [30]) ?  RTL___rd_val___1__h6558 : RTL____theResult_____1_fst__h6569 ; 
  assign  RTL____theResult_____1_fst__h6597 = RTL___rs1_val_bypassed__h3337 & RTL____theResult___snd__h7382 ; 
  assign  RTL____theResult____h10743 =( RTL___delta_CPI_instrs__h10742 ==64'd0) ?  RTL___delta_CPI_instrs___1__h10778 : RTL___delta_CPI_instrs__h10742 ; 
  assign  RTL____theResult___snd__h7382 =( RTL___near_mem$imem_instr [6:0]==7'b0010011) ?  RTL___SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 : RTL___rs2_val__h5339 ; 
  assign  RTL___alu_outputs___1_addr__h5365 = RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  ?  RTL___alu_outputs___1_val2__h5367 : RTL___alu_outputs___1_val1__h5386 ; 
  assign  RTL___alu_outputs___1_addr__h5385 = RTL___near_mem$imem_pc +{{11{ RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 [20]}}, RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 }; 
  assign  RTL___alu_outputs___1_addr__h5410 ={ RTL___eaddr__h5553 [31:1],1'd0}; 
  assign  RTL___alu_outputs___1_addr__h5583 = RTL___rs1_val_bypassed__h3337 +{{20{ RTL___near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 [11]}}, RTL___near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 }; 
  assign  RTL___alu_outputs___1_exc_code__h5362 = RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616  ? 4'd0:4'd2; 
  assign  RTL___alu_outputs___1_exc_code__h5843 =( RTL___near_mem$imem_instr [14:12]==3'b0) ? (( RTL___near_mem$imem_instr [11:7]==5'd0&& RTL___near_mem$imem_instr [19:15]==5'd0) ?  RTL___CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4 :4'd2):4'd2; 
  assign  RTL___alu_outputs___1_val1__h5386 = RTL___near_mem$imem_pc +32'd4; 
  assign  RTL___alu_outputs___1_val1__h5480 =( RTL___near_mem$imem_instr [14:12]==3'b001) ?  RTL___rd_val__h7278 :( RTL___near_mem$imem_instr [30] ?  RTL___rd_val__h7352 : RTL___rd_val__h7330 ); 
  assign  RTL___alu_outputs___1_val1__h5516 =( RTL___near_mem$imem_instr [14:12]==3'b0&&( RTL___near_mem$imem_instr [6:0]!=7'b0110011||! RTL___near_mem$imem_instr [30])) ?  RTL___rd_val___1__h6550 : RTL____theResult_____1_fst__h6562 ; 
  assign  RTL___alu_outputs___1_val1__h5847 = RTL___near_mem$imem_instr [14] ? {27'd0, RTL___near_mem$imem_instr [19:15]}: RTL___rs1_val_bypassed__h3337 ; 
  assign  RTL___alu_outputs___1_val2__h5367 = RTL___near_mem$imem_pc +{{19{ RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 [12]}}, RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 }; 
  assign  RTL___cpi__h10745 = RTL___x__h10744 /64'd10; 
  assign  RTL___cpifrac__h10746 = RTL___x__h10744 %64'd10; 
  assign  RTL___csr_regfile_interrupt_pending_rg_cur_priv_9_07_ETC___d779 =( RTL___csr_regfile$interrupt_pending [4]|| RTL___csr_regfile$nmi_pending )&&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )|| RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd2&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0; 
  assign  RTL___csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 = RTL___delta_CPI_cycles__h10741 *64'd10; 
  assign  RTL___cur_verbosity__h1827 =( RTL___csr_regfile$read_csr_minstret < RTL___cfg_logdelay ) ? 4'd0: RTL___cfg_verbosity ; 
  assign  RTL___data_to_stage2_addr__h5215 = RTL___x_out_data_to_stage2_addr__h5223 ; 
  assign  RTL___delta_CPI_cycles__h10741 = RTL___csr_regfile$read_csr_mcycle - RTL___rg_start_CPI_cycles ; 
  assign  RTL___delta_CPI_instrs___1__h10778 = RTL___delta_CPI_instrs__h10742 +64'd1; 
  assign  RTL___delta_CPI_instrs__h10742 = RTL___csr_regfile$read_csr_minstret - RTL___rg_start_CPI_instrs ; 
  assign  RTL___eaddr__h5553 = RTL___rs1_val_bypassed__h3337 + RTL___SEXT_near_mem_imem_instr__59_BITS_31_TO_20_02___d303 ; 
  assign  RTL___fall_through_pc__h5175 = RTL___near_mem$imem_pc +( RTL___near_mem$imem_is_i32_not_i16  ? 32'd4:32'd2); 
  assign  RTL___gpr_regfile_RDY_server_reset_request_put__59_A_ETC___d671 = RTL___gpr_regfile$RDY_server_reset_request_put && RTL___near_mem$RDY_server_reset_request_put && RTL___csr_regfile$RDY_server_reset_request_put && RTL___f_reset_reqs$EMPTY_N && RTL___stage1_f_reset_reqs$FULL_N && RTL___stage2_f_reset_reqs$FULL_N && RTL___stage3_f_reset_reqs$FULL_N ; 
  assign  RTL___gpr_regfile_RDY_server_reset_response_get__76__ETC___d688 = RTL___gpr_regfile$RDY_server_reset_response_get && RTL___near_mem$RDY_server_reset_response_get && RTL___csr_regfile$RDY_server_reset_response_get && RTL___stage1_f_reset_rsps$EMPTY_N && RTL___stage2_f_reset_rsps$EMPTY_N && RTL___stage3_f_reset_rsps$EMPTY_N && RTL___f_reset_rsps$FULL_N ; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd0; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd1; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10; 
  assign  RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 =( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd0&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd1&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd2&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd3&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd4&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd5&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd6&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd7&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd8&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd9&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 !=4'd10; 
  assign  RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 = RTL___near_mem$imem_instr [14:12]==3'b0&&( RTL___near_mem$imem_instr [6:0]!=7'b0110011||! RTL___near_mem$imem_instr [30])|| RTL___near_mem$imem_instr [14:12]==3'b0&& RTL___near_mem$imem_instr [6:0]==7'b0110011&& RTL___near_mem$imem_instr [30]|| RTL___near_mem$imem_instr [14:12]==3'b010|| RTL___near_mem$imem_instr [14:12]==3'b011|| RTL___near_mem$imem_instr [14:12]==3'b100|| RTL___near_mem$imem_instr [14:12]==3'b110|| RTL___near_mem$imem_instr [14:12]==3'b111; 
  assign  RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d616 =( RTL___near_mem$imem_instr [14:12]==3'b0|| RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b100|| RTL___near_mem$imem_instr [14:12]==3'b101|| RTL___near_mem$imem_instr [14:12]==3'b110|| RTL___near_mem$imem_instr [14:12]==3'b111)&& RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 && RTL___alu_outputs___1_val2__h5367 [1]; 
  assign  RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 = RTL___near_mem$imem_valid &&( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd1||! RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 &&! RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ); 
  assign  RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 = RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&( RTL___near_mem$imem_exc || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d274 && RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308 ); 
  assign  RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 = RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 ); 
  assign  RTL___near_memimem_instr_BITS_31_TO_20__q7 = RTL___near_mem$imem_instr [31:20]; 
  assign  RTL___near_memimem_instr_BITS_31_TO_25_CONCAT_near__ETC__q6 ={ RTL___near_mem$imem_instr [31:25], RTL___near_mem$imem_instr [11:7]}; 
  assign  RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q1 ={ RTL___near_mem$imem_instr [31], RTL___near_mem$imem_instr [7], RTL___near_mem$imem_instr [30:25], RTL___near_mem$imem_instr [11:8],1'b0}; 
  assign  RTL___near_memimem_instr_BIT_31_CONCAT_near_memime_ETC__q2 ={ RTL___near_mem$imem_instr [31], RTL___near_mem$imem_instr [19:12], RTL___near_mem$imem_instr [20], RTL___near_mem$imem_instr [30:21],1'b0}; 
  assign  RTL___output_stage2___1_bypass_rd_val__h4960 =(! RTL___near_mem$dmem_valid ||! RTL___near_mem$dmem_exc ) ? (( RTL___stage2_rg_stage2 [100:96]==5'd0) ?  RTL___stage2_rg_stage2 [63:32]: RTL___near_mem$dmem_word64 [31:0]): RTL___stage2_rg_stage2 [63:32]; 
  assign  RTL___rd_val___1__h6550 = RTL___rs1_val_bypassed__h3337 + RTL____theResult___snd__h7382 ; 
  assign  RTL___rd_val___1__h6558 = RTL___rs1_val_bypassed__h3337 - RTL____theResult___snd__h7382 ; 
  assign  RTL___rd_val___1__h6565 =(( RTL___rs1_val_bypassed__h3337 ^32'h80000000)<( RTL____theResult___snd__h7382 ^32'h80000000)) ? 32'd1:32'd0; 
  assign  RTL___rd_val___1__h6572 =( RTL___rs1_val_bypassed__h3337 < RTL____theResult___snd__h7382 ) ? 32'd1:32'd0; 
  assign  RTL___rd_val___1__h6579 = RTL___rs1_val_bypassed__h3337 ^ RTL____theResult___snd__h7382 ; 
  assign  RTL___rd_val___1__h6586 = RTL___rs1_val_bypassed__h3337 | RTL____theResult___snd__h7382 ; 
  assign  RTL___rd_val__h5072 =( RTL___stage3_rg_full && RTL___stage3_rg_stage3 [37]&& RTL___stage3_rg_stage3 [36:32]== RTL___near_mem$imem_instr [19:15]) ?  RTL___stage3_rg_stage3 [31:0]: RTL___gpr_regfile$read_rs1 ; 
  assign  RTL___rd_val__h5132 =( RTL___stage3_rg_full && RTL___stage3_rg_stage3 [37]&& RTL___stage3_rg_stage3 [36:32]== RTL___near_mem$imem_instr [24:20]) ?  RTL___stage3_rg_stage3 [31:0]: RTL___gpr_regfile$read_rs2 ; 
  assign  RTL___rd_val__h5523 ={ RTL___near_mem$imem_instr [31:12],12'h0}; 
  assign  RTL___rd_val__h5537 = RTL___near_mem$imem_pc + RTL___rd_val__h5523 ; 
  assign  RTL___rd_val__h7278 = RTL___rs1_val_bypassed__h3337 << RTL___shamt__h5467 ; 
  assign  RTL___rd_val__h7330 = RTL___rs1_val_bypassed__h3337 >> RTL___shamt__h5467 ; 
  assign  RTL___rd_val__h7352 = RTL___rs1_val_bypassed__h3337 >> RTL___shamt__h5467 |~(32'hFFFFFFFF>> RTL___shamt__h5467 )&{32{ RTL___rs1_val_bypassed__h3337 [31]}}; 
  assign  RTL___rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_EQ_0_ETC___d392 =( RTL___rg_cur_priv ==2'b11|| RTL___rg_cur_priv ==2'b01&&! RTL___csr_regfile$read_mstatus [21]|| RTL___rg_cur_priv ==2'b0&& RTL___csr_regfile$read_misa [13])&& RTL___near_mem$imem_instr [31:20]==12'b000100000101; 
  assign  RTL___rg_state_8_EQ_3_97_AND_NOT_csr_regfile_interru_ETC___d793 = RTL___rg_state ==4'd3&& RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d790 &&! RTL___stage3_rg_full && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0; 
  assign  RTL___rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 = RTL___rg_trap_info [67:36]== RTL___csr_regfile$csr_trap_actions [97:66]; 
  assign  RTL___rs1_val__h11213 =( RTL___rg_trap_instr [14:12]==3'b001) ?  RTL___rg_csr_val1 :{27'd0, RTL___rg_trap_instr [19:15]}; 
  assign  RTL___rs1_val_bypassed__h3337 =( RTL___near_mem$imem_instr [19:15]==5'd0) ? 32'd0: RTL___val__h5074 ; 
  assign  RTL___rs2_val__h5339 =( RTL___near_mem$imem_instr [24:20]==5'd0) ? 32'd0: RTL___val__h5134 ; 
  assign  RTL___shamt__h5467 =( RTL___near_mem$imem_instr [6:0]==7'b0010011) ?  RTL___near_mem$imem_instr [24:20]: RTL___rs2_val__h5339 [4:0]; 
  assign  RTL___trap_info_tval__h6925 = RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d649  ?  RTL___near_mem$imem_instr : RTL___IF_IF_near_mem_imem_instr__59_BITS_6_TO_0_79_E_ETC___d655 ; 
  assign  RTL___val__h5074 =( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd2&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d161 ) ?  RTL___x_out_bypass_rd_val__h4969 : RTL___rd_val__h5072 ; 
  assign  RTL___val__h5134 =( RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd2&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d163 ) ?  RTL___x_out_bypass_rd_val__h4969 : RTL___rd_val__h5132 ; 
  assign  RTL___value__h6967 = RTL___near_mem$imem_exc  ?  RTL___near_mem$imem_tval : RTL___trap_info_tval__h6925 ; 
  assign  RTL___x__h10744 = RTL___csr_regfile_read_csr_mcycle__8_MINUS_rg_start__ETC___d818 [63:0]/ RTL____theResult____h10743 ; 
  assign  RTL___x_exc_code__h15410 =( RTL___csr_regfile$interrupt_pending [4]&&! RTL___csr_regfile$nmi_pending ) ?  RTL___csr_regfile$interrupt_pending [3:0]:4'd0; 
  assign  RTL___x_out_bypass_rd_val__h4969 =( RTL___stage2_rg_stage2 [102:101]==2'd0) ?  RTL___stage2_rg_stage2 [63:32]: RTL___output_stage2___1_bypass_rd_val__h4960 ; 
  assign  RTL___x_out_data_to_stage2_rd__h5222 =( RTL___near_mem$imem_instr [6:0]==7'b1100011) ? 5'd0: RTL___near_mem$imem_instr [11:7]; 
  assign  RTL___x_out_data_to_stage2_val2__h5225 =( RTL___near_mem$imem_instr [6:0]==7'b1100011) ?  RTL___alu_outputs___1_val2__h5367 : RTL___rs2_val__h5339 ; 
  assign  RTL___x_out_next_pc__h5189 = RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  ?  RTL___data_to_stage2_addr__h5215 : RTL___fall_through_pc__h5175 ; 
  assign  RTL___x_out_trap_info_exc_code__h6928 = RTL___near_mem$imem_exc  ?  RTL___near_mem$imem_exc_code : RTL___alu_outputs_exc_code__h5862 ; 
  assign  RTL___y__h12191 =~ RTL___rs1_val__h11920 ; 
  always @(  RTL___stage2_rg_stage2  )
         begin 
             case ( RTL___stage2_rg_stage2 [102:101])
              2 'd0,2'd1: 
                  RTL___x_out_data_to_stage3_rd__h4667  = RTL___stage2_rg_stage2 [100:96];
              default : 
                  RTL___x_out_data_to_stage3_rd__h4667  =5'd0;endcase
         end
  always @(   RTL___stage2_rg_stage2            or   RTL___near_mem$dmem_word64  )
         begin 
             case ( RTL___stage2_rg_stage2 [102:101])
              2 'd0: 
                  RTL___x_out_data_to_stage3_rd_val__h4668  = RTL___stage2_rg_stage2 [63:32];
              2 'd1: 
                  RTL___x_out_data_to_stage3_rd_val__h4668  = RTL___near_mem$dmem_word64 [31:0];
              default : 
                  RTL___x_out_data_to_stage3_rd_val__h4668  = RTL___stage2_rg_stage2 [63:32];endcase
         end
  always @(   RTL___rg_trap_instr            or   RTL___rg_csr_val1  )
         begin 
             case ( RTL___rg_trap_instr [14:12])
              3 'b010,3'b011: 
                  RTL___rs1_val__h11920  = RTL___rg_csr_val1 ;
              default : 
                  RTL___rs1_val__h11920  ={27'd0, RTL___rg_trap_instr [19:15]};endcase
         end
  always @(  RTL___rg_cur_priv  )
         begin 
             case ( RTL___rg_cur_priv )
              2 'b0: 
                  RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd8;
              2 'b01: 
                  RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd9;
              default : 
                  RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  =4'd11;endcase
         end
  always @(   RTL___near_mem$imem_instr            or   RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3  )
         begin 
             case ( RTL___near_mem$imem_instr [31:20])
              12 'b0: 
                  RTL___CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  = RTL___CASE_rg_cur_priv_0b0_8_0b1_9_11__q3 ;
              12 'b000000000001: 
                  RTL___CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  =4'd3;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_31_TO_20_0b0_CAS_ETC__q4  =4'd2;endcase
         end
  always @(     RTL___stage2_rg_stage2                or   RTL___near_mem$dmem_valid            or   RTL___near_mem$dmem_exc           or   RTL___IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137  )
         begin 
             case ( RTL___stage2_rg_stage2 [102:101])
              2 'd0: 
                  RTL___CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =2'd2;
              2 'd1: 
                  RTL___CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =(! RTL___near_mem$dmem_valid ||! RTL___near_mem$dmem_exc ) ?  RTL___IF_stage2_rg_stage2_4_BITS_100_TO_96_13_EQ_0_3_ETC___d137 :2'd0;
              default : 
                  RTL___CASE_stage2_rg_stage2_BITS_102_TO_101_0_2_1_IF_ETC__q5  =2'd0;endcase
         end
  always @(     RTL___near_mem$imem_instr                or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220            or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216           or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b001: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  =! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b100: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b101: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  =! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b110: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  = RTL___near_mem$imem_instr [14:12]==3'b111&&! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;endcase
         end
  always @(       RTL___near_mem$imem_instr                    or   RTL___alu_outputs___1_addr__h5583              or   RTL___eaddr__h5553             or   RTL___alu_outputs___1_addr__h5365            or   RTL___alu_outputs___1_addr__h5410           or   RTL___alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL___x_out_data_to_stage2_addr__h5223  = RTL___eaddr__h5553 ;
              7 'b1100011: 
                  RTL___x_out_data_to_stage2_addr__h5223  = RTL___alu_outputs___1_addr__h5365 ;
              7 'b1100111: 
                  RTL___x_out_data_to_stage2_addr__h5223  = RTL___alu_outputs___1_addr__h5410 ;
              7 'b1101111: 
                  RTL___x_out_data_to_stage2_addr__h5223  = RTL___alu_outputs___1_addr__h5385 ;
              default : 
                  RTL___x_out_data_to_stage2_addr__h5223  = RTL___alu_outputs___1_addr__h5583 ;endcase
         end
  always @(       RTL___near_mem$imem_instr                    or   RTL____theResult_____1_fst__h6597              or   RTL___rd_val___1__h6565             or   RTL___rd_val___1__h6572            or   RTL___rd_val___1__h6579           or   RTL___rd_val___1__h6586  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b010: 
                  RTL____theResult_____1_fst__h6569  = RTL___rd_val___1__h6565 ;
              3 'b011: 
                  RTL____theResult_____1_fst__h6569  = RTL___rd_val___1__h6572 ;
              3 'b100: 
                  RTL____theResult_____1_fst__h6569  = RTL___rd_val___1__h6579 ;
              3 'b110: 
                  RTL____theResult_____1_fst__h6569  = RTL___rd_val___1__h6586 ;
              default : 
                  RTL____theResult_____1_fst__h6569  = RTL____theResult_____1_fst__h6597 ;endcase
         end
  always @(     RTL___near_mem$imem_instr                or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220            or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216           or   RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b001: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d216 ;
              3 'b100: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b101: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d218 ;
              3 'b110: 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  =! RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291  = RTL___near_mem$imem_instr [14:12]!=3'b111|| RTL___IF_near_mem_imem_instr__59_BITS_19_TO_15_60_EQ_ETC___d220 ;endcase
         end
  always @(   RTL___near_mem$imem_instr            or   RTL___NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8  = RTL___NOT_near_mem_imem_instr__59_BITS_14_TO_12_81_E_ETC___d252 ;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_N_ETC__q8  = RTL___near_mem$imem_instr [6:0]!=7'b0110111&& RTL___near_mem$imem_instr [6:0]!=7'b0010111&&(( RTL___near_mem$imem_instr [6:0]==7'b0000011) ?  RTL___near_mem$imem_instr [14:12]!=3'b0&& RTL___near_mem$imem_instr [14:12]!=3'b100&& RTL___near_mem$imem_instr [14:12]!=3'b001&& RTL___near_mem$imem_instr [14:12]!=3'b101&& RTL___near_mem$imem_instr [14:12]!=3'b010: RTL___near_mem$imem_instr [6:0]!=7'b0100011|| RTL___near_mem$imem_instr [14:12]!=3'b0&& RTL___near_mem$imem_instr [14:12]!=3'b001&& RTL___near_mem$imem_instr [14:12]!=3'b010);endcase
         end
  always @(      RTL___near_mem$imem_instr                  or   RTL___eaddr__h5553             or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285            or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291           or   RTL___alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285 || RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ;
              7 'b1101111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL___alu_outputs___1_addr__h5385 [1];
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d308  = RTL___near_mem$imem_instr [6:0]!=7'b1100111|| RTL___eaddr__h5553 [1];endcase
         end
  always @(   RTL___near_mem$imem_instr            or   RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9  = RTL___near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_0b_ETC___d328 ;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_6_TO_0_0b10011_n_ETC__q9  = RTL___near_mem$imem_instr [6:0]==7'b0110111|| RTL___near_mem$imem_instr [6:0]==7'b0010111||(( RTL___near_mem$imem_instr [6:0]==7'b0000011) ?  RTL___near_mem$imem_instr [14:12]==3'b0|| RTL___near_mem$imem_instr [14:12]==3'b100|| RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b101|| RTL___near_mem$imem_instr [14:12]==3'b010: RTL___near_mem$imem_instr [6:0]==7'b0100011&&( RTL___near_mem$imem_instr [14:12]==3'b0|| RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b010));endcase
         end
  always @(       RTL___near_mem$imem_instr                    or   RTL___eaddr__h5553              or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291             or   RTL___alu_outputs___1_val2__h5367            or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227           or   RTL___alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  =( RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d291 ||! RTL___alu_outputs___1_val2__h5367 [1])&&( RTL___near_mem$imem_instr [14:12]==3'b0|| RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b100|| RTL___near_mem$imem_instr [14:12]==3'b101|| RTL___near_mem$imem_instr [14:12]==3'b110|| RTL___near_mem$imem_instr [14:12]==3'b111)&& RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227 ;
              7 'b1101111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  =! RTL___alu_outputs___1_addr__h5385 [1];
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352  = RTL___near_mem$imem_instr [6:0]==7'b1100111&&! RTL___eaddr__h5553 [1];endcase
         end
  always @(    RTL___near_mem$imem_instr              or   RTL___rg_cur_priv           or   RTL___IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394  )
         begin 
             case ( RTL___near_mem$imem_instr [31:20])
              12 'b0,12'b000000000001: 
                  RTL___IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  =4'd11;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  =( RTL___rg_cur_priv ==2'b11&& RTL___near_mem$imem_instr [31:20]==12'b001100000010) ? 4'd7: RTL___IF_rg_cur_priv_9_EQ_0b11_75_OR_rg_cur_priv_9_E_ETC___d394 ;endcase
         end
  always @(  RTL___near_mem$imem_instr  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0,3'b001,3'b010,3'b100,3'b101: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10  =4'd0;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10  =4'd11;endcase
         end
  always @(  RTL___near_mem$imem_instr  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd4;
              3 'b001: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd5;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11  =4'd11;endcase
         end
  always @(  RTL___near_mem$imem_instr  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0,3'b001,3'b010: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12  =4'd0;
              default : 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12  =4'd11;endcase
         end
  always @(   RTL___near_mem$imem_instr            or   RTL___IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396  )
         begin 
             case ( RTL___near_mem$imem_instr [14:12])
              3 'b0: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =( RTL___near_mem$imem_instr [11:7]==5'd0&& RTL___near_mem$imem_instr [19:15]==5'd0) ?  RTL___IF_near_mem_imem_instr__59_BITS_31_TO_20_02_EQ_ETC___d396 :4'd11;
              3 'b001,3'b101: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd2;
              3 'b010,3'b011,3'b110,3'b111: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd3;
              3 'd4: 
                  RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  =4'd11;endcase
         end
  always @(       RTL___near_mem$imem_instr                    or   RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10              or   RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11             or   RTL___IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362            or   RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12           or   RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q10 ;
              7 'b0001111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_4_0_ETC__q11 ;
              7 'b0010011,7'b0110011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL___IF_NOT_near_mem_imem_instr__59_BITS_14_TO_12_8_ETC___d362 ;
              7 'b0010111,7'b0110111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  =4'd0;
              7 'b0100011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_0_0_ETC__q12 ;
              7 'b1110011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  = RTL___CASE_near_memimem_instr_BITS_14_TO_12_0b0_IF__ETC__q13 ;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409  =4'd11;endcase
         end
  always @(       RTL___near_mem$imem_instr                    or   RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409              or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285             or   RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227            or   RTL___eaddr__h5553           or   RTL___alu_outputs___1_addr__h5385  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b1100011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d285  ? 4'd11:( RTL___IF_near_mem_imem_instr__59_BITS_14_TO_12_81_EQ_ETC___d227  ? 4'd1:4'd0);
              7 'b1100111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL___eaddr__h5553 [1] ? 4'd11:4'd1;
              7 'b1101111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  = RTL___alu_outputs___1_addr__h5385 [1] ? 4'd11:4'd1;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d413  =(( RTL___near_mem$imem_instr [6:0]==7'b0010011|| RTL___near_mem$imem_instr [6:0]==7'b0110011)&&( RTL___near_mem$imem_instr [14:12]==3'b001|| RTL___near_mem$imem_instr [14:12]==3'b101)) ? ( RTL___near_mem$imem_instr [25] ? 4'd11:4'd0): RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d409 ;endcase
         end
  always @(  RTL___near_mem$imem_instr  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0000011: 
                  RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd1;
              7 'b0010011,7'b0010111,7'b0110011,7'b0110111,7'b1100011,7'b1100111,7'b1101111: 
                  RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd0;
              default : 
                  RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491  =2'd2;endcase
         end
  always @(    RTL___near_mem$imem_instr              or   RTL___alu_outputs___1_exc_code__h5362           or   RTL___alu_outputs___1_exc_code__h5843  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0000011,7'b0001111,7'b0010011,7'b0010111,7'b0100011,7'b0110011,7'b0110111: 
                  RTL___alu_outputs_exc_code__h5862  =4'd2;
              7 'b1100011: 
                  RTL___alu_outputs_exc_code__h5862  = RTL___alu_outputs___1_exc_code__h5362 ;
              7 'b1100111,7'b1101111: 
                  RTL___alu_outputs_exc_code__h5862  =4'd0;
              7 'b1110011: 
                  RTL___alu_outputs_exc_code__h5862  = RTL___alu_outputs___1_exc_code__h5843 ;
              default : 
                  RTL___alu_outputs_exc_code__h5862  =4'd2;endcase
         end
  always @(      RTL___near_mem$imem_instr                  or   RTL___alu_outputs___1_val1__h5847             or   RTL___alu_outputs___1_val1__h5516            or   RTL___rd_val__h5537           or   RTL___rd_val__h5523  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b0010011,7'b0110011: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL___alu_outputs___1_val1__h5516 ;
              7 'b0010111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL___rd_val__h5537 ;
              7 'b0110111: 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL___rd_val__h5523 ;
              default : 
                  RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d570  = RTL___alu_outputs___1_val1__h5847 ;endcase
         end
  always @(    RTL___near_mem$imem_instr              or   RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571           or   RTL___alu_outputs___1_val1__h5386  )
         begin 
             case ( RTL___near_mem$imem_instr [6:0])
              7 'b1100111,7'b1101111: 
                  RTL___x_out_data_to_stage2_val1__h5224  = RTL___alu_outputs___1_val1__h5386 ;
              default : 
                  RTL___x_out_data_to_stage2_val1__h5224  = RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d571 ;endcase
         end
  always @( posedge  RTL___CLK )
         begin 
             if ( RTL___RST_N ==1'b0)
                 begin  
                     RTL___cfg_logdelay  <=64'd0; 
                     RTL___cfg_verbosity  <=4'd0; 
                     RTL___rg_cur_priv  <=2'b11; 
                     RTL___rg_retiring  <=1'd0; 
                     RTL___rg_run_on_reset  <=1'd0; 
                     RTL___rg_state  <=4'd0; 
                     RTL___s1_to_s2  <=1'd0; 
                     RTL___s2_to_s3  <=1'd0; 
                     RTL___s3_deq  <=1'd0; 
                     RTL___stage1_rg_full  <=1'd0; 
                     RTL___stage2_rg_full  <=1'd0; 
                     RTL___stage2_rg_resetting  <=1'd0; 
                     RTL___stage3_rg_full  <=1'd0;
                 end 
              else 
                 begin 
                     if ( RTL___cfg_logdelay$EN ) 
                         RTL___cfg_logdelay  <= RTL___cfg_logdelay$D_IN ;
                     if ( RTL___cfg_verbosity$EN ) 
                         RTL___cfg_verbosity  <= RTL___cfg_verbosity$D_IN ;
                     if ( RTL___rg_cur_priv$EN ) 
                         RTL___rg_cur_priv  <= RTL___rg_cur_priv$D_IN ;
                     if ( RTL___rg_retiring$EN ) 
                         RTL___rg_retiring  <= RTL___rg_retiring$D_IN ;
                     if ( RTL___rg_run_on_reset$EN ) 
                         RTL___rg_run_on_reset  <= RTL___rg_run_on_reset$D_IN ;
                     if ( RTL___rg_state$EN ) 
                         RTL___rg_state  <= RTL___rg_state$D_IN ;
                     if ( RTL___s1_to_s2$EN ) 
                         RTL___s1_to_s2  <= RTL___s1_to_s2$D_IN ;
                     if ( RTL___s2_to_s3$EN ) 
                         RTL___s2_to_s3  <= RTL___s2_to_s3$D_IN ;
                     if ( RTL___s3_deq$EN ) 
                         RTL___s3_deq  <= RTL___s3_deq$D_IN ;
                     if ( RTL___stage1_rg_full$EN ) 
                         RTL___stage1_rg_full  <= RTL___stage1_rg_full$D_IN ;
                     if ( RTL___stage2_rg_full$EN ) 
                         RTL___stage2_rg_full  <= RTL___stage2_rg_full$D_IN ;
                     if ( RTL___stage2_rg_resetting$EN ) 
                         RTL___stage2_rg_resetting  <= RTL___stage2_rg_resetting$D_IN ;
                     if ( RTL___stage3_rg_full$EN ) 
                         RTL___stage3_rg_full  <= RTL___stage3_rg_full$D_IN ;
                 end 
             if ( RTL___rg_csr_pc$EN ) 
                 RTL___rg_csr_pc  <= RTL___rg_csr_pc$D_IN ;
             if ( RTL___rg_csr_val1$EN ) 
                 RTL___rg_csr_val1  <= RTL___rg_csr_val1$D_IN ;
             if ( RTL___rg_mstatus_MXR$EN ) 
                 RTL___rg_mstatus_MXR  <= RTL___rg_mstatus_MXR$D_IN ;
             if ( RTL___rg_next_pc$EN ) 
                 RTL___rg_next_pc  <= RTL___rg_next_pc$D_IN ;
             if ( RTL___rg_sstatus_SUM$EN ) 
                 RTL___rg_sstatus_SUM  <= RTL___rg_sstatus_SUM$D_IN ;
             if ( RTL___rg_start_CPI_cycles$EN ) 
                 RTL___rg_start_CPI_cycles  <= RTL___rg_start_CPI_cycles$D_IN ;
             if ( RTL___rg_start_CPI_instrs$EN ) 
                 RTL___rg_start_CPI_instrs  <= RTL___rg_start_CPI_instrs$D_IN ;
             if ( RTL___rg_trap_info$EN ) 
                 RTL___rg_trap_info  <= RTL___rg_trap_info$D_IN ;
             if ( RTL___rg_trap_instr$EN ) 
                 RTL___rg_trap_instr  <= RTL___rg_trap_instr$D_IN ;
             if ( RTL___rg_trap_interrupt$EN ) 
                 RTL___rg_trap_interrupt  <= RTL___rg_trap_interrupt$D_IN ;
             if ( RTL___stage2_rg_stage2$EN ) 
                 RTL___stage2_rg_stage2  <= RTL___stage2_rg_stage2$D_IN ;
             if ( RTL___stage3_rg_stage3$EN ) 
                 RTL___stage3_rg_stage3  <= RTL___stage3_rg_stage3$D_IN ;
         end
  always @( negedge  RTL___CLK )
         begin #0;
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$display("================================================================");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$display("%0d: Pipeline State:  minstret:%0d  cur_priv:%0d  mstatus:%0x", RTL___csr_regfile$read_csr_mcycle , RTL___csr_regfile$read_csr_minstret , RTL___rg_cur_priv , RTL___csr_regfile$read_mstatus );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("    ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("MStatus{","sd:%0d", RTL___csr_regfile$read_mstatus [14:13]==2'h3|| RTL___csr_regfile$read_mstatus [16:15]==2'h3);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___csr_regfile$read_misa [27:26]==2'd2)$write(" sxl:%0d uxl:%0d",2'd0,2'd0);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___csr_regfile$read_misa [27:26]!=2'd2)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" tsr:%0d", RTL___csr_regfile$read_mstatus [22]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" tw:%0d", RTL___csr_regfile$read_mstatus [21]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" tvm:%0d", RTL___csr_regfile$read_mstatus [20]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" mxr:%0d", RTL___csr_regfile$read_mstatus [19]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" sum:%0d", RTL___csr_regfile$read_mstatus [18]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" mprv:%0d", RTL___csr_regfile$read_mstatus [17]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" xs:%0d", RTL___csr_regfile$read_mstatus [16:15]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" fs:%0d", RTL___csr_regfile$read_mstatus [14:13]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" mpp:%0d", RTL___csr_regfile$read_mstatus [12:11]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" spp:%0d", RTL___csr_regfile$read_mstatus [8]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" pies:%0d_%0d%0d", RTL___csr_regfile$read_mstatus [7], RTL___csr_regfile$read_mstatus [5], RTL___csr_regfile$read_mstatus [4]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write(" ies:%0d_%0d%0d", RTL___csr_regfile$read_mstatus [3], RTL___csr_regfile$read_mstatus [1], RTL___csr_regfile$read_mstatus [0]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("    Stage3: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("Output_Stage3");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage3_rg_full )$write(" PIPE");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage3_rg_full )$write(" EMPTY");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("        Bypass  to Stage1: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("Bypass {");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&(! RTL___stage3_rg_full ||! RTL___stage3_rg_stage3 [37]))$write("Rd -");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage3_rg_full && RTL___stage3_rg_stage3 [37])$write("Rd %0d ", RTL___stage3_rg_stage3 [36:32],"rd_val:%h", RTL___stage3_rg_stage3 [31:0]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$display("    Stage2: pc 0x%08h instr 0x%08h priv %0d", RTL___stage2_rg_stage2 [166:135], RTL___stage2_rg_stage2 [134:103], RTL___stage2_rg_stage2 [168:167]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("        ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("Output_Stage2"," EMPTY");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("Output_Stage2"," BUSY: pc:%0h", RTL___stage2_rg_stage2 [166:135]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Output_Stage2"," NONPIPE: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("Output_Stage2"," PIPE: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("data_to_Stage3 {pc:%h  instr:%h  priv:%0d\n", RTL___stage2_rg_stage2 [166:135], RTL___stage2_rg_stage2 [134:103], RTL___stage2_rg_stage2 [168:167]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("        rd_valid:");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3&& RTL___stage2_rg_stage2 [102:101]!=2'd0&&(! RTL___near_mem$dmem_valid || RTL___near_mem$dmem_exc ))$write("False");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___NOT_IF_stage2_rg_full_3_THEN_IF_stage2_rg_stag_ETC___d109 )$write("True");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("  grd:%0d  rd_val:%h\n", RTL___x_out_data_to_stage3_rd__h4667 , RTL___x_out_data_to_stage3_rd_val__h4668 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Trap_Info { ","epc: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___stage2_rg_stage2 [166:135]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","exc_code: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___near_mem$dmem_exc_code );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","tval: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___stage2_rg_stage2 [95:64]," }");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(" ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("Trap_Info { ","epc: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___stage2_rg_stage2 [166:135]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","exc_code: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___near_mem$dmem_exc_code );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write(", ","tval: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd1)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd3)$write("'h%h", RTL___stage2_rg_stage2 [95:64]," }");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd1&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 !=2'd3)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("        Bypass  to Stage1: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("Bypass {");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd0)$write("Rd -");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd0)$write("Rd %0d ", RTL___stage2_rg_stage2 [100:96]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd0)$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 ==2'd1)$write("-");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd0&& RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d142 !=2'd1)$write("rd_val:%h", RTL___x_out_bypass_rd_val__h4969 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("}");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$display("    Stage1: pc 0x%08h instr 0x%08h priv %0d", RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("        ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("Output_Stage1"," BUSY pc:%h", RTL___near_mem$imem_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("Output_Stage1"," NONPIPE: pc:%h", RTL___near_mem$imem_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("Output_Stage1");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("Output_Stage1"," EMPTY");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write(" PIPE: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd0)$write("CONTROL_STRAIGHT");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd1)$write("CONTROL_BRANCH");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd2)$write("CONTROL_CSRR_W");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd3)$write("CONTROL_CSRR_S_or_C");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd4)$write("CONTROL_FENCE");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd5)$write("CONTROL_FENCE_I");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd6)$write("CONTROL_SFENCE_VMA");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd7)$write("CONTROL_MRET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd8)$write("CONTROL_SRET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd9)$write("CONTROL_URET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d415 ==4'd10)$write("CONTROL_WFI");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___NOT_near_mem_imem_exc__78_13_AND_IF_near_mem_i_ETC___d481 )$write("CONTROL_TRAP");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write(" ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("}");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("data_to_Stage 2 {pc:%h  instr:%h  priv:%0d\n", RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("            op_stage2:");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd0)$write("OP_Stage2_ALU");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1)$write("OP_Stage2_LD");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 &&! RTL___near_mem$imem_exc &&( RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d343 || RTL___IF_near_mem_imem_instr__59_BITS_6_TO_0_79_EQ_0_ETC___d352 )&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd0&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1)$write("OP_Stage2_ST");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("  rd:%0d\n", RTL___x_out_data_to_stage2_rd__h5222 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("            addr:%h  val1:%h  val2:%h}", RTL___x_out_data_to_stage2_addr__h5223 , RTL___x_out_data_to_stage2_val1__h5224 , RTL___x_out_data_to_stage2_val2__h5225 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(" ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d578 )$write("CONTROL_STRAIGHT");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d581 )$write("CONTROL_BRANCH");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d584 )$write("CONTROL_CSRR_W");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d587 )$write("CONTROL_CSRR_S_or_C");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d590 )$write("CONTROL_FENCE");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d593 )$write("CONTROL_FENCE_I");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d596 )$write("CONTROL_SFENCE_VMA");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d599 )$write("CONTROL_MRET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d602 )$write("CONTROL_SRET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d605 )$write("CONTROL_URET");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d608 )$write("CONTROL_WFI");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d177 && RTL___near_mem_imem_exc__78_OR_IF_near_mem_imem_inst_ETC___d611 )$write("CONTROL_TRAP");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(" ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("Trap_Info { ","epc: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL___near_mem$imem_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(", ","exc_code: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL___x_out_trap_info_exc_code__h6928 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write(", ","tval: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d311 )$write("'h%h", RTL___value__h6967 ," }");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___near_mem_imem_valid__57_AND_NOT_IF_stage2_rg_f_ETC___d355 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe && RTL___stage1_rg_full && RTL___NOT_near_mem_imem_valid__57_58_OR_IF_stage2_rg_ETC___d166 )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe &&! RTL___stage1_rg_full )$write("");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_show_pipe )$display("----------------");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___soc_map$m_pc_reset_value [31:0]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_complete && RTL___rg_run_on_reset )$display("%0d: %m.rl_reset_complete: restart at PC = 0x%0h", RTL___csr_regfile$read_csr_mcycle , RTL___soc_map$m_pc_reset_value [31:0]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_complete &&! RTL___rg_run_on_reset )$display("%0d: %m.rl_reset_complete: entering DEBUG_MODE", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_pipe", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___stage3_rg_full && RTL___stage3_rg_stage3 [37]&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S3.fa_deq: write GRd 0x%0h, rd_val 0x%0h", RTL___stage3_rg_stage3 [36:32], RTL___stage3_rg_stage3 [31:0]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("    S3.enq: ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("data_to_Stage3 {pc:%h  instr:%h  priv:%0d\n", RTL___stage2_rg_stage2 [166:135], RTL___stage2_rg_stage2 [134:103], RTL___stage2_rg_stage2 [168:167]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("        rd_valid:");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL___stage2_rg_stage2 [102:101]!=2'd0&&(! RTL___near_mem$dmem_valid || RTL___near_mem$dmem_exc ))$write("False");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d730 )$write("True");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("  grd:%0d  rd_val:%h\n", RTL___x_out_data_to_stage3_rd__h4667 , RTL___x_out_data_to_stage3_rd_val__h4668 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___IF_stage2_rg_full_3_THEN_IF_stage2_rg_stage2_4_ETC___d86 ==2'd2&& RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___stage2_rg_stage2 [166:135], RTL___stage2_rg_stage2 [134:103], RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("    CPU_Stage2.enq (Data_Stage1_to_Stage2) ");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("data_to_Stage 2 {pc:%h  instr:%h  priv:%0d\n", RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("            op_stage2:");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd0)$write("OP_Stage2_ALU");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 ==2'd1)$write("OP_Stage2_LD");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 && RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd0&& RTL___IF_NOT_stage1_rg_full_55_56_OR_NOT_near_mem_im_ETC___d491 !=2'd1)$write("OP_Stage2_ST");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("  rd:%0d\n", RTL___x_out_data_to_stage2_rd__h5222 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("            addr:%h  val1:%h  val2:%h}", RTL___x_out_data_to_stage2_addr__h5223 , RTL___x_out_data_to_stage2_val1__h5224 , RTL___x_out_data_to_stage2_val2__h5225 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d737 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$write("\n");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_pipe && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d716 && RTL___NOT_csr_regfile_interrupt_pending_rg_cur_priv__ETC___d756 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___x_out_next_pc__h5189 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage2_nonpipe && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage2_nonpipe", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_trap && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_trap", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap && RTL___rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$display("%0d: %m.rl_stage1_trap: Tight infinite trap loop: pc 0x%0x instr 0x%08x", RTL___csr_regfile$read_csr_mcycle , RTL___csr_regfile$csr_trap_actions [97:66], RTL___rg_trap_instr );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap && RTL___rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$display("CPI: %0d.%0d = (%0d/%0d) since last 'continue'", RTL___cpi__h10745 , RTL___cpifrac__h10746 , RTL___delta_CPI_cycles__h10741 , RTL____theResult____h10743 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap && RTL___rg_trap_info_04_BITS_67_TO_36_05_EQ_csr_regfil_ETC___d814 )$finish(32'd0);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___rg_trap_info [67:36], RTL___rg_trap_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap && RTL___cur_verbosity__h1827 !=4'd0)$display("    mcause:0x%0h  epc 0x%0h  tval:0x%0h  next_pc 0x%0h, new_priv %0d new_mstatus 0x%0h", RTL___csr_regfile$csr_trap_actions [33:2], RTL___rg_trap_info [67:36], RTL___rg_trap_info [31:0], RTL___csr_regfile$csr_trap_actions [97:66], RTL___csr_regfile$csr_trap_actions [1:0], RTL___csr_regfile$csr_trap_actions [65:34]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_W && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_W", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_W_2", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___rg_csr_pc , RTL___rg_trap_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 && RTL___csr_regfile$access_permitted_1 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S1: write CSRRW/CSRRWI Rs1 %0d Rs1_val 0x%0h csr 0x%0h csr_val 0x%0h Rd %0d", RTL___rg_trap_instr [19:15], RTL___rs1_val__h11213 , RTL___rg_trap_instr [31:20], RTL___csr_regfile$read_csr [31:0], RTL___rg_trap_instr [11:7]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_W_2 &&! RTL___csr_regfile$access_permitted_1 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    rl_stage1_CSRR_W: Trap on CSR permissions: Rs1 %0d Rs1_val 0x%0h csr 0x%0h Rd %0d", RTL___rg_trap_instr [19:15], RTL___rs1_val__h11213 , RTL___rg_trap_instr [31:20], RTL___rg_trap_instr [11:7]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_S_or_C", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_CSRR_S_or_C_2", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___rg_csr_pc , RTL___rg_trap_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 && RTL___csr_regfile$access_permitted_2 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    S1: write CSRR_S_or_C: Rs1 %0d Rs1_val 0x%0h csr 0x%0h csr_val 0x%0h Rd %0d", RTL___rg_trap_instr [19:15], RTL___rs1_val__h11920 , RTL___rg_trap_instr [31:20], RTL___csr_regfile$read_csr [31:0], RTL___rg_trap_instr [11:7]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_CSRR_S_or_C_2 &&! RTL___csr_regfile$access_permitted_2 && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    rl_stage1_CSRR_S_or_C: Trap on CSR permissions: Rs1 %0d Rs1_val 0x%0h csr 0x%0h Rd %0d", RTL___rg_trap_instr [19:15], RTL___rs1_val__h11920 , RTL___rg_trap_instr [31:20], RTL___rg_trap_instr [11:7]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___x_out_next_pc__h5189 );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_restart_after_csrrx && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: rl_stage1_restart_after_csrrx: minstret:%0d  pc:%0x  cur_priv:%0d", RTL___csr_regfile$read_csr_mcycle , RTL___csr_regfile$read_csr_minstret , RTL___x_out_next_pc__h5189 , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_xRET && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_xRET", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_xRET && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_xRET && RTL___cur_verbosity__h1827 !=4'd0)$display("    xRET: next_pc:0x%0h  new mstatus:0x%0h  new priv:%0d", RTL___csr_regfile$csr_ret_actions [65:34], RTL___csr_regfile$csr_ret_actions [31:0], RTL___csr_regfile$csr_ret_actions [33:32]);
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE_I && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE_I", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE_I && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE_I && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE_I", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE_I && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_FENCE_I", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE_I && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___rg_next_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE_I && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_FENCE_I");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_FENCE && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_FENCE", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_FENCE", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___rg_next_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_FENCE && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_FENCE");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_SFENCE_VMA", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_SFENCE_VMA && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_SFENCE_VMA", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_finish_SFENCE_VMA", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___rg_next_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_finish_SFENCE_VMA && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_finish_SFENCE_VMA");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_WFI && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_WFI", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_WFI && RTL___cur_verbosity__h1827 ==4'd1)$display("instret:%0d  PC:0x%0h  instr:0x%0h  priv:%0d", RTL___csr_regfile$read_csr_minstret , RTL___near_mem$imem_pc , RTL___near_mem$imem_instr , RTL___rg_cur_priv );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_WFI && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU.rl_stage1_WFI");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_WFI_resume && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_WFI_resume", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_WFI_resume && RTL___cur_verbosity__h1827 !=4'd0)$display("    WFI resume");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_WFI_resume && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___rg_next_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_from_WFI && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_reset_from_WFI", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_trap_fetch && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("    CPU_Stage1.enq: 0x%08h", RTL___rg_next_pc );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_stage1_interrupt && RTL___NOT_IF_csr_regfile_read_csr_minstret__1_ULT_cf_ETC___d17 )$display("%0d: %m.rl_stage1_interrupt", RTL___csr_regfile$read_csr_mcycle );
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start )$display("================================================================");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start )$write("CPU: Bluespec  RISC-V  Piccolo  v3.0");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start )$display(" (RV32)");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start )$display("Copyright (c) 2016-2019 Bluespec, Inc. All Rights Reserved.");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start )$display("================================================================");
             if ( RTL___RST_N !=1'b0)
                 if ( RTL___WILL_FIRE_RL_rl_reset_start && RTL___cur_verbosity__h1827 !=4'd0)$display("%0d: %m.rl_reset_start", RTL___csr_regfile$read_csr_mcycle );
         end
  assign  RTL___RTL__DOT__s3_deq$D_IN = RTL___s3_deq$D_IN ; 
  assign  RTL___RTL__DOT__near_mem$dmem_exc = RTL___near_mem$dmem_exc ; 
  assign  RTL___RTL__DOT__near_mem$imem_pc = RTL___near_mem$imem_pc ; 
  assign  RTL___RTL__DOT__near_mem$imem_instr = RTL___near_mem$imem_instr ; 
  assign  RTL___RTL__DOT__near_mem$dmem_req_addr = RTL___near_mem$dmem_req_addr ; 
  assign  RTL___RTL__DOT__stage2_rg_stage2 = RTL___stage2_rg_stage2 ; 
  assign  RTL___RTL__DOT__rg_cur_priv = RTL___rg_cur_priv ; 
  assign  RTL___RTL__DOT__near_mem$EN_dmem_req = RTL___near_mem$EN_dmem_req ; 
  assign  RTL___RTL__DOT__near_mem$dmem_req_f3 = RTL___near_mem$dmem_req_f3 ; 
  assign  RTL___RTL__DOT__s1_to_s2$D_IN = RTL___s1_to_s2$D_IN ; 
  assign  RTL___RTL__DOT__near_mem$dmem_word64 = RTL___near_mem$dmem_word64 ; 
  assign  RTL___RTL__DOT__stage3_rg_full = RTL___stage3_rg_full ; 
  assign  RTL___RTL__DOT__rg_trap_instr = RTL___rg_trap_instr ; 
  assign  RTL___RTL__DOT__near_mem$dmem_req_op = RTL___near_mem$dmem_req_op ; 
  assign  RTL___RTL__DOT__s2_to_s3$D_IN = RTL___s2_to_s3$D_IN ; 
  assign  RTL___RTL__DOT__rg_retiring$EN = RTL___rg_retiring$EN ; 
  assign  RTL___RTL__DOT__rg_state = RTL___rg_state ; 
  assign  RTL___RTL__DOT__s3_deq$EN = RTL___s3_deq$EN ; 
  assign  RTL___RTL__DOT__s1_to_s2$EN = RTL___s1_to_s2$EN ; 
  assign  RTL___RTL__DOT__s2_to_s3$EN = RTL___s2_to_s3$EN ; 
  assign  RTL___RTL__DOT__rg_run_on_reset = RTL___rg_run_on_reset ; 
  assign  RTL___RTL__DOT__stage1_rg_full = RTL___stage1_rg_full ; 
  assign  RTL___RTL__DOT__stage2_rg_full = RTL___stage2_rg_full ; 
  assign  RTL___RTL__DOT__near_mem$dmem_req_store_value = RTL___near_mem$dmem_req_store_value ;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_4_;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__DOT__near_mem$dmem_req_op = RTL___RTL__DOT__near_mem$dmem_req_op;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__rg_trap_instr = RTL___RTL__DOT__rg_trap_instr;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__full_reg;
    assign RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__stage2_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem$dmem_req_store_value = RTL___RTL__DOT__near_mem$dmem_req_store_value;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_20_;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_word64 = RTL___RTL__DOT__near_mem$dmem_word64;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_5_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_addr;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__stage3_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__s1_to_s2$D_IN = RTL___RTL__DOT__s1_to_s2$D_IN;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_9_;
    assign RTL__DOT__stage2_rg_full = RTL___RTL__DOT__stage2_rg_full;
    assign RTL__DOT__csr_regfile__DOT__rg_state = RTL___RTL__DOT__csr_regfile__DOT__rg_state;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__DOT__stage1_rg_full = RTL___RTL__DOT__stage1_rg_full;
    assign RTL__DOT__stage1_f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__stage1_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_14_;
    assign RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__stage1_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__DOT__stage1_f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__stage1_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__rg_run_on_reset = RTL___RTL__DOT__rg_run_on_reset;
    assign RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__stage1_f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__stage3_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__s2_to_s3$EN = RTL___RTL__DOT__s2_to_s3$EN;
    assign RTL__DOT__near_mem$dmem_req_f3 = RTL___RTL__DOT__near_mem$dmem_req_f3;
    assign RTL__DOT__s1_to_s2$EN = RTL___RTL__DOT__s1_to_s2$EN;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_3_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_8_;
    assign RTL__DOT__s3_deq$EN = RTL___RTL__DOT__s3_deq$EN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__rg_state = RTL___RTL__DOT__rg_state;
    assign RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__gpr_regfile__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__rg_retiring$EN = RTL___RTL__DOT__rg_retiring$EN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_resp__DOT__empty_reg;
    assign RTL__DOT__s2_to_s3$D_IN = RTL___RTL__DOT__s2_to_s3$D_IN;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_11_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_18_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_24_;
    assign RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__stage2_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_2_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__DOT__stage2_f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__stage2_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_data__DOT__full_reg;
    assign RTL__DOT__stage3_f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__stage3_f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__stage3_rg_full = RTL___RTL__DOT__stage3_rg_full;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_28_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_17_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__full_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_21_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_22_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_23_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_25_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_27_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_29_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_31_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_6_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_1_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_10_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_7_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_12_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_15_;
    assign RTL__DOT__stage2_rg_stage2 = RTL___RTL__DOT__stage2_rg_stage2;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_19_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_13_;
    assign RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__csr_regfile__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__csr_regfile__DOT__rg_nmi = RTL___RTL__DOT__csr_regfile__DOT__rg_nmi;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__rg_pa;
    assign RTL__DOT__near_mem$EN_dmem_req = RTL___RTL__DOT__near_mem$EN_dmem_req;
    assign RTL__DOT__stage2_f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__stage2_f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__rg_cur_priv = RTL___RTL__DOT__rg_cur_priv;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_26_;
    assign RTL__DOT__f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__stage3_f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__f_reset_rsps__DOT__empty_reg = RTL___RTL__DOT__f_reset_rsps__DOT__empty_reg;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_30_;
    assign RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_ = RTL___RTL__DOT__gpr_regfile__DOT__regfile__DOT__arr_16_;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_wr_resp__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_req_addr = RTL___RTL__DOT__near_mem$dmem_req_addr;
    assign RTL__DOT__near_mem$imem_instr = RTL___RTL__DOT__near_mem$imem_instr;
    assign RTL__DOT__f_reset_reqs__DOT__full_reg = RTL___RTL__DOT__f_reset_reqs__DOT__full_reg;
    assign RTL__DOT__near_mem$imem_pc = RTL___RTL__DOT__near_mem$imem_pc;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_reset_rsps__DOT__full_reg;
    assign RTL__DOT__near_mem$dmem_exc = RTL___RTL__DOT__near_mem$dmem_exc;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_addr__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__f_fabric_write_reqs__DOT__empty_reg;
    assign RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__icache__DOT__master_xactor_f_wr_addr__DOT__full_reg;
    assign RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg = RTL___RTL__DOT__near_mem__DOT__dcache__DOT__master_xactor_f_rd_data__DOT__full_reg;
    assign RTL__DOT__s3_deq$D_IN = RTL___RTL__DOT__s3_deq$D_IN;
    assign RTL___CLK = clk;
    assign RTL___RST_N = ~rst;
    assign RTL___hart0_server_reset_request_put = __VLG_I_hart0_server_reset_request_put;
    assign RTL___EN_hart0_server_reset_request_put = __VLG_I_EN_hart0_server_reset_request_put;
    assign __VLG_O_RDY_hart0_server_reset_request_put = RTL___RDY_hart0_server_reset_request_put;
    assign RTL___EN_hart0_server_reset_response_get = __VLG_I_EN_hart0_server_reset_response_get;
    assign __VLG_O_hart0_server_reset_response_get = RTL___hart0_server_reset_response_get;
    assign __VLG_O_RDY_hart0_server_reset_response_get = RTL___RDY_hart0_server_reset_response_get;
    assign __VLG_O_imem_master_awvalid = RTL___imem_master_awvalid;
    assign __VLG_O_imem_master_awid = RTL___imem_master_awid;
    assign __VLG_O_imem_master_awaddr = RTL___imem_master_awaddr;
    assign __VLG_O_imem_master_awlen = RTL___imem_master_awlen;
    assign __VLG_O_imem_master_awsize = RTL___imem_master_awsize;
    assign __VLG_O_imem_master_awburst = RTL___imem_master_awburst;
    assign __VLG_O_imem_master_awlock = RTL___imem_master_awlock;
    assign __VLG_O_imem_master_awcache = RTL___imem_master_awcache;
    assign __VLG_O_imem_master_awprot = RTL___imem_master_awprot;
    assign __VLG_O_imem_master_awqos = RTL___imem_master_awqos;
    assign __VLG_O_imem_master_awregion = RTL___imem_master_awregion;
    assign RTL___imem_master_awready = __VLG_I_imem_master_awready;
    assign __VLG_O_imem_master_wvalid = RTL___imem_master_wvalid;
    assign __VLG_O_imem_master_wdata = RTL___imem_master_wdata;
    assign __VLG_O_imem_master_wstrb = RTL___imem_master_wstrb;
    assign __VLG_O_imem_master_wlast = RTL___imem_master_wlast;
    assign RTL___imem_master_wready = __VLG_I_imem_master_wready;
    assign RTL___imem_master_bvalid = __VLG_I_imem_master_bvalid;
    assign RTL___imem_master_bid = __VLG_I_imem_master_bid;
    assign RTL___imem_master_bresp = __VLG_I_imem_master_bresp;
    assign __VLG_O_imem_master_bready = RTL___imem_master_bready;
    assign __VLG_O_imem_master_arvalid = RTL___imem_master_arvalid;
    assign __VLG_O_imem_master_arid = RTL___imem_master_arid;
    assign __VLG_O_imem_master_araddr = RTL___imem_master_araddr;
    assign __VLG_O_imem_master_arlen = RTL___imem_master_arlen;
    assign __VLG_O_imem_master_arsize = RTL___imem_master_arsize;
    assign __VLG_O_imem_master_arburst = RTL___imem_master_arburst;
    assign __VLG_O_imem_master_arlock = RTL___imem_master_arlock;
    assign __VLG_O_imem_master_arcache = RTL___imem_master_arcache;
    assign __VLG_O_imem_master_arprot = RTL___imem_master_arprot;
    assign __VLG_O_imem_master_arqos = RTL___imem_master_arqos;
    assign __VLG_O_imem_master_arregion = RTL___imem_master_arregion;
    assign RTL___imem_master_arready = __VLG_I_imem_master_arready;
    assign RTL___imem_master_rvalid = __VLG_I_imem_master_rvalid;
    assign RTL___imem_master_rid = __VLG_I_imem_master_rid;
    assign RTL___imem_master_rdata = __VLG_I_imem_master_rdata;
    assign RTL___imem_master_rresp = __VLG_I_imem_master_rresp;
    assign RTL___imem_master_rlast = __VLG_I_imem_master_rlast;
    assign __VLG_O_imem_master_rready = RTL___imem_master_rready;
    assign __VLG_O_dmem_master_awvalid = RTL___dmem_master_awvalid;
    assign __VLG_O_dmem_master_awid = RTL___dmem_master_awid;
    assign __VLG_O_dmem_master_awaddr = RTL___dmem_master_awaddr;
    assign __VLG_O_dmem_master_awlen = RTL___dmem_master_awlen;
    assign __VLG_O_dmem_master_awsize = RTL___dmem_master_awsize;
    assign __VLG_O_dmem_master_awburst = RTL___dmem_master_awburst;
    assign __VLG_O_dmem_master_awlock = RTL___dmem_master_awlock;
    assign __VLG_O_dmem_master_awcache = RTL___dmem_master_awcache;
    assign __VLG_O_dmem_master_awprot = RTL___dmem_master_awprot;
    assign __VLG_O_dmem_master_awqos = RTL___dmem_master_awqos;
    assign __VLG_O_dmem_master_awregion = RTL___dmem_master_awregion;
    assign RTL___dmem_master_awready = __VLG_I_dmem_master_awready;
    assign __VLG_O_dmem_master_wvalid = RTL___dmem_master_wvalid;
    assign __VLG_O_dmem_master_wdata = RTL___dmem_master_wdata;
    assign __VLG_O_dmem_master_wstrb = RTL___dmem_master_wstrb;
    assign __VLG_O_dmem_master_wlast = RTL___dmem_master_wlast;
    assign RTL___dmem_master_wready = __VLG_I_dmem_master_wready;
    assign RTL___dmem_master_bvalid = __VLG_I_dmem_master_bvalid;
    assign RTL___dmem_master_bid = __VLG_I_dmem_master_bid;
    assign RTL___dmem_master_bresp = __VLG_I_dmem_master_bresp;
    assign __VLG_O_dmem_master_bready = RTL___dmem_master_bready;
    assign __VLG_O_dmem_master_arvalid = RTL___dmem_master_arvalid;
    assign __VLG_O_dmem_master_arid = RTL___dmem_master_arid;
    assign __VLG_O_dmem_master_araddr = RTL___dmem_master_araddr;
    assign __VLG_O_dmem_master_arlen = RTL___dmem_master_arlen;
    assign __VLG_O_dmem_master_arsize = RTL___dmem_master_arsize;
    assign __VLG_O_dmem_master_arburst = RTL___dmem_master_arburst;
    assign __VLG_O_dmem_master_arlock = RTL___dmem_master_arlock;
    assign __VLG_O_dmem_master_arcache = RTL___dmem_master_arcache;
    assign __VLG_O_dmem_master_arprot = RTL___dmem_master_arprot;
    assign __VLG_O_dmem_master_arqos = RTL___dmem_master_arqos;
    assign __VLG_O_dmem_master_arregion = RTL___dmem_master_arregion;
    assign RTL___dmem_master_arready = __VLG_I_dmem_master_arready;
    assign RTL___dmem_master_rvalid = __VLG_I_dmem_master_rvalid;
    assign RTL___dmem_master_rid = __VLG_I_dmem_master_rid;
    assign RTL___dmem_master_rdata = __VLG_I_dmem_master_rdata;
    assign RTL___dmem_master_rresp = __VLG_I_dmem_master_rresp;
    assign RTL___dmem_master_rlast = __VLG_I_dmem_master_rlast;
    assign __VLG_O_dmem_master_rready = RTL___dmem_master_rready;
    assign RTL___m_external_interrupt_req_set_not_clear = __VLG_II_m_external_interrupt_req_set_not_clear;
    assign RTL___s_external_interrupt_req_set_not_clear = __VLG_II_s_external_interrupt_req_set_not_clear;
    assign RTL___software_interrupt_req_set_not_clear = __VLG_II_software_interrupt_req_set_not_clear;
    assign RTL___timer_interrupt_req_set_not_clear = __VLG_II_timer_interrupt_req_set_not_clear;
    assign RTL___nmi_req_set_not_clear = __VLG_II_nmi_req_set_not_clear;
    assign RTL___set_verbosity_verbosity = __VLG_I_set_verbosity_verbosity;
    assign RTL___set_verbosity_logdelay = __VLG_I_set_verbosity_logdelay;
    assign RTL___EN_set_verbosity = __VLG_I_EN_set_verbosity;
    assign __VLG_O_RDY_set_verbosity = RTL___RDY_set_verbosity;
    
assign __all_assert_wire__ = (variable_map_assert__p118__) && (variable_map_assert__p119__) && (variable_map_assert__p120__) && (variable_map_assert__p121__) && (variable_map_assert__p122__) && (variable_map_assert__p123__) && (variable_map_assert__p124__) && (variable_map_assert__p125__) && (variable_map_assert__p126__) && (variable_map_assert__p127__) && (variable_map_assert__p128__) && (variable_map_assert__p129__) && (variable_map_assert__p130__) && (variable_map_assert__p131__) && (variable_map_assert__p132__) && (variable_map_assert__p133__) && (variable_map_assert__p134__) && (variable_map_assert__p135__) && (variable_map_assert__p136__) && (variable_map_assert__p137__) && (variable_map_assert__p138__) && (variable_map_assert__p139__) && (variable_map_assert__p140__) && (variable_map_assert__p141__) && (variable_map_assert__p142__) && (variable_map_assert__p143__) && (variable_map_assert__p144__) && (variable_map_assert__p145__) && (variable_map_assert__p146__) && (variable_map_assert__p147__) && (variable_map_assert__p148__) && (variable_map_assert__p149__) && (variable_map_assert__p150__) && (variable_map_assert__p151__) && (variable_map_assert__p152__) ;
normalassert: assert property ( __all_assert_wire__ ); // the only assertion 

assign __all_assume_wire__ = (input_map_assume___p0__)&& (invariant_assume__p1__)&& (invariant_assume__p2__)&& (invariant_assume__p3__)&& (invariant_assume__p4__)&& (invariant_assume__p5__)&& (invariant_assume__p6__)&& (invariant_assume__p7__)&& (invariant_assume__p8__)&& (invariant_assume__p9__)&& (invariant_assume__p10__)&& (invariant_assume__p11__)&& (invariant_assume__p12__)&& (invariant_assume__p13__)&& (invariant_assume__p14__)&& (invariant_assume__p15__)&& (invariant_assume__p16__)&& (invariant_assume__p17__)&& (invariant_assume__p18__)&& (invariant_assume__p19__)&& (invariant_assume__p20__)&& (invariant_assume__p21__)&& (invariant_assume__p22__)&& (invariant_assume__p23__)&& (invariant_assume__p24__)&& (invariant_assume__p25__)&& (invariant_assume__p26__)&& (invariant_assume__p27__)&& (invariant_assume__p28__)&& (invariant_assume__p29__)&& (invariant_assume__p30__)&& (invariant_assume__p31__)&& (invariant_assume__p32__)&& (issue_decode__p33__)&& (issue_valid__p34__)&& (noreset__p35__)&& (post_value_holder__p36__)&& (post_value_holder__p37__)&& (post_value_holder__p38__)&& (post_value_holder__p39__)&& (post_value_holder__p40__)&& (post_value_holder__p41__)&& (post_value_holder__p42__)&& (post_value_holder__p43__)&& (post_value_holder__p44__)&& (post_value_holder__p45__)&& (post_value_holder__p46__)&& (post_value_holder__p47__)&& (post_value_holder__p48__)&& (post_value_holder__p49__)&& (post_value_holder__p50__)&& (post_value_holder__p51__)&& (post_value_holder__p52__)&& (post_value_holder__p53__)&& (post_value_holder__p54__)&& (post_value_holder__p55__)&& (post_value_holder__p56__)&& (post_value_holder__p57__)&& (post_value_holder__p58__)&& (post_value_holder__p59__)&& (post_value_holder__p60__)&& (post_value_holder__p61__)&& (post_value_holder__p62__)&& (post_value_holder__p63__)&& (post_value_holder__p64__)&& (post_value_holder__p65__)&& (post_value_holder__p66__)&& (post_value_holder__p67__)&& (post_value_holder__p68__)&& (post_value_holder__p69__)&& (post_value_holder__p70__)&& (post_value_holder__p71__)&& (post_value_holder__p72__)&& (post_value_holder__p73__)&& (rfassumptions__p74__)&& (rfassumptions__p75__)&& (rfassumptions__p76__)&& (variable_map_assume___p77__)&& (variable_map_assume___p78__)&& (variable_map_assume___p79__)&& (variable_map_assume___p80__)&& (variable_map_assume___p81__)&& (variable_map_assume___p82__)&& (variable_map_assume___p83__)&& (variable_map_assume___p84__)&& (variable_map_assume___p85__)&& (variable_map_assume___p86__)&& (variable_map_assume___p87__)&& (variable_map_assume___p88__)&& (variable_map_assume___p89__)&& (variable_map_assume___p90__)&& (variable_map_assume___p91__)&& (variable_map_assume___p92__)&& (variable_map_assume___p93__)&& (variable_map_assume___p94__)&& (variable_map_assume___p95__)&& (variable_map_assume___p96__)&& (variable_map_assume___p97__)&& (variable_map_assume___p98__)&& (variable_map_assume___p99__)&& (variable_map_assume___p100__)&& (variable_map_assume___p101__)&& (variable_map_assume___p102__)&& (variable_map_assume___p103__)&& (variable_map_assume___p104__)&& (variable_map_assume___p105__)&& (variable_map_assume___p106__)&& (variable_map_assume___p107__)&& (variable_map_assume___p108__)&& (variable_map_assume___p109__)&& (variable_map_assume___p110__)&& (variable_map_assume___p111__)&& (variable_map_assume___p112__)&& (variable_map_assume___p113__)&& (variable_map_assume___p114__)&& (variable_map_assume___p115__)&& (variable_map_assume___p116__)&& (variable_map_assume___p117__) ;
all_assume: assume property ( __all_assume_wire__ ); // the only sanity assertion 

assign __sanitycheck_wire__ = (post_value_holder_overly_constrained__p153__) && (post_value_holder_overly_constrained__p154__) && (post_value_holder_overly_constrained__p155__) && (post_value_holder_overly_constrained__p156__) && (post_value_holder_overly_constrained__p157__) && (post_value_holder_overly_constrained__p158__) && (post_value_holder_overly_constrained__p159__) && (post_value_holder_overly_constrained__p160__) && (post_value_holder_overly_constrained__p161__) && (post_value_holder_overly_constrained__p162__) && (post_value_holder_overly_constrained__p163__) && (post_value_holder_overly_constrained__p164__) && (post_value_holder_overly_constrained__p165__) && (post_value_holder_overly_constrained__p166__) && (post_value_holder_overly_constrained__p167__) && (post_value_holder_overly_constrained__p168__) && (post_value_holder_overly_constrained__p169__) && (post_value_holder_overly_constrained__p170__) && (post_value_holder_overly_constrained__p171__) && (post_value_holder_overly_constrained__p172__) && (post_value_holder_overly_constrained__p173__) && (post_value_holder_overly_constrained__p174__) && (post_value_holder_overly_constrained__p175__) && (post_value_holder_overly_constrained__p176__) && (post_value_holder_overly_constrained__p177__) && (post_value_holder_overly_constrained__p178__) && (post_value_holder_overly_constrained__p179__) && (post_value_holder_overly_constrained__p180__) && (post_value_holder_overly_constrained__p181__) && (post_value_holder_overly_constrained__p182__) && (post_value_holder_overly_constrained__p183__) && (post_value_holder_overly_constrained__p184__) && (post_value_holder_overly_constrained__p185__) && (post_value_holder_overly_constrained__p186__) && (post_value_holder_overly_constrained__p187__) && (post_value_holder_overly_constrained__p188__) && (post_value_holder_overly_constrained__p189__) && (post_value_holder_overly_constrained__p190__) && (post_value_holder_triggered__p191__) && (post_value_holder_triggered__p192__) && (post_value_holder_triggered__p193__) && (post_value_holder_triggered__p194__) && (post_value_holder_triggered__p195__) && (post_value_holder_triggered__p196__) && (post_value_holder_triggered__p197__) && (post_value_holder_triggered__p198__) && (post_value_holder_triggered__p199__) && (post_value_holder_triggered__p200__) && (post_value_holder_triggered__p201__) && (post_value_holder_triggered__p202__) && (post_value_holder_triggered__p203__) && (post_value_holder_triggered__p204__) && (post_value_holder_triggered__p205__) && (post_value_holder_triggered__p206__) && (post_value_holder_triggered__p207__) && (post_value_holder_triggered__p208__) && (post_value_holder_triggered__p209__) && (post_value_holder_triggered__p210__) && (post_value_holder_triggered__p211__) && (post_value_holder_triggered__p212__) && (post_value_holder_triggered__p213__) && (post_value_holder_triggered__p214__) && (post_value_holder_triggered__p215__) && (post_value_holder_triggered__p216__) && (post_value_holder_triggered__p217__) && (post_value_holder_triggered__p218__) && (post_value_holder_triggered__p219__) && (post_value_holder_triggered__p220__) && (post_value_holder_triggered__p221__) && (post_value_holder_triggered__p222__) && (post_value_holder_triggered__p223__) && (post_value_holder_triggered__p224__) && (post_value_holder_triggered__p225__) && (post_value_holder_triggered__p226__) && (post_value_holder_triggered__p227__) && (post_value_holder_triggered__p228__) ;
sanitycheck: assert property ( __sanitycheck_wire__ ); // the only assumption 

always @(posedge clk) begin
   if(rst) begin
       __auxvar10__recorder <= ____auxvar10__recorder_init__;
       __auxvar10__recorder_sn_condmet <= 1'b0;
       __auxvar11__recorder <= ____auxvar11__recorder_init__;
       __auxvar11__recorder_sn_condmet <= 1'b0;
       __auxvar12__recorder <= ____auxvar12__recorder_init__;
       __auxvar12__recorder_sn_condmet <= 1'b0;
       __auxvar13__recorder <= ____auxvar13__recorder_init__;
       __auxvar13__recorder_sn_condmet <= 1'b0;
       __auxvar14__recorder <= ____auxvar14__recorder_init__;
       __auxvar14__recorder_sn_condmet <= 1'b0;
       __auxvar15__recorder <= ____auxvar15__recorder_init__;
       __auxvar15__recorder_sn_condmet <= 1'b0;
       __auxvar16__recorder <= ____auxvar16__recorder_init__;
       __auxvar16__recorder_sn_condmet <= 1'b0;
       __auxvar17__recorder <= ____auxvar17__recorder_init__;
       __auxvar17__recorder_sn_condmet <= 1'b0;
       __auxvar18__recorder <= ____auxvar18__recorder_init__;
       __auxvar18__recorder_sn_condmet <= 1'b0;
       __auxvar19__recorder <= ____auxvar19__recorder_init__;
       __auxvar19__recorder_sn_condmet <= 1'b0;
       __auxvar1__recorder <= ____auxvar1__recorder_init__;
       __auxvar1__recorder_sn_condmet <= 1'b0;
       __auxvar20__recorder <= ____auxvar20__recorder_init__;
       __auxvar20__recorder_sn_condmet <= 1'b0;
       __auxvar21__recorder <= ____auxvar21__recorder_init__;
       __auxvar21__recorder_sn_condmet <= 1'b0;
       __auxvar22__recorder <= ____auxvar22__recorder_init__;
       __auxvar22__recorder_sn_condmet <= 1'b0;
       __auxvar23__recorder <= ____auxvar23__recorder_init__;
       __auxvar23__recorder_sn_condmet <= 1'b0;
       __auxvar24__recorder <= ____auxvar24__recorder_init__;
       __auxvar24__recorder_sn_condmet <= 1'b0;
       __auxvar25__recorder <= ____auxvar25__recorder_init__;
       __auxvar25__recorder_sn_condmet <= 1'b0;
       __auxvar26__recorder <= ____auxvar26__recorder_init__;
       __auxvar26__recorder_sn_condmet <= 1'b0;
       __auxvar27__recorder <= ____auxvar27__recorder_init__;
       __auxvar27__recorder_sn_condmet <= 1'b0;
       __auxvar28__recorder <= ____auxvar28__recorder_init__;
       __auxvar28__recorder_sn_condmet <= 1'b0;
       __auxvar29__recorder <= ____auxvar29__recorder_init__;
       __auxvar29__recorder_sn_condmet <= 1'b0;
       __auxvar2__recorder <= ____auxvar2__recorder_init__;
       __auxvar2__recorder_sn_condmet <= 1'b0;
       __auxvar30__recorder <= ____auxvar30__recorder_init__;
       __auxvar30__recorder_sn_condmet <= 1'b0;
       __auxvar31__recorder <= ____auxvar31__recorder_init__;
       __auxvar31__recorder_sn_condmet <= 1'b0;
       __auxvar32__recorder <= ____auxvar32__recorder_init__;
       __auxvar32__recorder_sn_condmet <= 1'b0;
       __auxvar33__recorder <= ____auxvar33__recorder_init__;
       __auxvar33__recorder_sn_condmet <= 1'b0;
       __auxvar34__recorder <= ____auxvar34__recorder_init__;
       __auxvar34__recorder_sn_condmet <= 1'b0;
       __auxvar35__recorder <= ____auxvar35__recorder_init__;
       __auxvar35__recorder_sn_condmet <= 1'b0;
       __auxvar36__recorder <= ____auxvar36__recorder_init__;
       __auxvar36__recorder_sn_condmet <= 1'b0;
       __auxvar37__recorder <= ____auxvar37__recorder_init__;
       __auxvar37__recorder_sn_condmet <= 1'b0;
       __auxvar38__recorder <= ____auxvar38__recorder_init__;
       __auxvar38__recorder_sn_condmet <= 1'b0;
       __auxvar3__recorder <= ____auxvar3__recorder_init__;
       __auxvar3__recorder_sn_condmet <= 1'b0;
       __auxvar4__recorder <= ____auxvar4__recorder_init__;
       __auxvar4__recorder_sn_condmet <= 1'b0;
       __auxvar5__recorder <= ____auxvar5__recorder_init__;
       __auxvar5__recorder_sn_condmet <= 1'b0;
       __auxvar6__recorder <= ____auxvar6__recorder_init__;
       __auxvar6__recorder_sn_condmet <= 1'b0;
       __auxvar7__recorder <= ____auxvar7__recorder_init__;
       __auxvar7__recorder_sn_condmet <= 1'b0;
       __auxvar8__recorder <= ____auxvar8__recorder_init__;
       __auxvar8__recorder_sn_condmet <= 1'b0;
       __auxvar9__recorder <= ____auxvar9__recorder_init__;
       __auxvar9__recorder_sn_condmet <= 1'b0;
       __auxvar0__delay_d_1<= 0;
       monitor_s1_already<= 1'b0;
       monitor_s2<= 1'b0;
       monitor_s3<= 1'b0;
       monitor_s4<= 1'b0;
   end
   else if(1) begin
       __auxvar10__recorder <= __auxvar10__recorder;
       if (__auxvar10__recorder_sn_cond ) begin __auxvar10__recorder_sn_condmet <= 1'b1; __auxvar10__recorder_sn_vhold <= __auxvar10__recorder_sn_value; end
       __auxvar11__recorder <= __auxvar11__recorder;
       if (__auxvar11__recorder_sn_cond ) begin __auxvar11__recorder_sn_condmet <= 1'b1; __auxvar11__recorder_sn_vhold <= __auxvar11__recorder_sn_value; end
       __auxvar12__recorder <= __auxvar12__recorder;
       if (__auxvar12__recorder_sn_cond ) begin __auxvar12__recorder_sn_condmet <= 1'b1; __auxvar12__recorder_sn_vhold <= __auxvar12__recorder_sn_value; end
       __auxvar13__recorder <= __auxvar13__recorder;
       if (__auxvar13__recorder_sn_cond ) begin __auxvar13__recorder_sn_condmet <= 1'b1; __auxvar13__recorder_sn_vhold <= __auxvar13__recorder_sn_value; end
       __auxvar14__recorder <= __auxvar14__recorder;
       if (__auxvar14__recorder_sn_cond ) begin __auxvar14__recorder_sn_condmet <= 1'b1; __auxvar14__recorder_sn_vhold <= __auxvar14__recorder_sn_value; end
       __auxvar15__recorder <= __auxvar15__recorder;
       if (__auxvar15__recorder_sn_cond ) begin __auxvar15__recorder_sn_condmet <= 1'b1; __auxvar15__recorder_sn_vhold <= __auxvar15__recorder_sn_value; end
       __auxvar16__recorder <= __auxvar16__recorder;
       if (__auxvar16__recorder_sn_cond ) begin __auxvar16__recorder_sn_condmet <= 1'b1; __auxvar16__recorder_sn_vhold <= __auxvar16__recorder_sn_value; end
       __auxvar17__recorder <= __auxvar17__recorder;
       if (__auxvar17__recorder_sn_cond ) begin __auxvar17__recorder_sn_condmet <= 1'b1; __auxvar17__recorder_sn_vhold <= __auxvar17__recorder_sn_value; end
       __auxvar18__recorder <= __auxvar18__recorder;
       if (__auxvar18__recorder_sn_cond ) begin __auxvar18__recorder_sn_condmet <= 1'b1; __auxvar18__recorder_sn_vhold <= __auxvar18__recorder_sn_value; end
       __auxvar19__recorder <= __auxvar19__recorder;
       if (__auxvar19__recorder_sn_cond ) begin __auxvar19__recorder_sn_condmet <= 1'b1; __auxvar19__recorder_sn_vhold <= __auxvar19__recorder_sn_value; end
       __auxvar1__recorder <= __auxvar1__recorder;
       if (__auxvar1__recorder_sn_cond ) begin __auxvar1__recorder_sn_condmet <= 1'b1; __auxvar1__recorder_sn_vhold <= __auxvar1__recorder_sn_value; end
       __auxvar20__recorder <= __auxvar20__recorder;
       if (__auxvar20__recorder_sn_cond ) begin __auxvar20__recorder_sn_condmet <= 1'b1; __auxvar20__recorder_sn_vhold <= __auxvar20__recorder_sn_value; end
       __auxvar21__recorder <= __auxvar21__recorder;
       if (__auxvar21__recorder_sn_cond ) begin __auxvar21__recorder_sn_condmet <= 1'b1; __auxvar21__recorder_sn_vhold <= __auxvar21__recorder_sn_value; end
       __auxvar22__recorder <= __auxvar22__recorder;
       if (__auxvar22__recorder_sn_cond ) begin __auxvar22__recorder_sn_condmet <= 1'b1; __auxvar22__recorder_sn_vhold <= __auxvar22__recorder_sn_value; end
       __auxvar23__recorder <= __auxvar23__recorder;
       if (__auxvar23__recorder_sn_cond ) begin __auxvar23__recorder_sn_condmet <= 1'b1; __auxvar23__recorder_sn_vhold <= __auxvar23__recorder_sn_value; end
       __auxvar24__recorder <= __auxvar24__recorder;
       if (__auxvar24__recorder_sn_cond ) begin __auxvar24__recorder_sn_condmet <= 1'b1; __auxvar24__recorder_sn_vhold <= __auxvar24__recorder_sn_value; end
       __auxvar25__recorder <= __auxvar25__recorder;
       if (__auxvar25__recorder_sn_cond ) begin __auxvar25__recorder_sn_condmet <= 1'b1; __auxvar25__recorder_sn_vhold <= __auxvar25__recorder_sn_value; end
       __auxvar26__recorder <= __auxvar26__recorder;
       if (__auxvar26__recorder_sn_cond ) begin __auxvar26__recorder_sn_condmet <= 1'b1; __auxvar26__recorder_sn_vhold <= __auxvar26__recorder_sn_value; end
       __auxvar27__recorder <= __auxvar27__recorder;
       if (__auxvar27__recorder_sn_cond ) begin __auxvar27__recorder_sn_condmet <= 1'b1; __auxvar27__recorder_sn_vhold <= __auxvar27__recorder_sn_value; end
       __auxvar28__recorder <= __auxvar28__recorder;
       if (__auxvar28__recorder_sn_cond ) begin __auxvar28__recorder_sn_condmet <= 1'b1; __auxvar28__recorder_sn_vhold <= __auxvar28__recorder_sn_value; end
       __auxvar29__recorder <= __auxvar29__recorder;
       if (__auxvar29__recorder_sn_cond ) begin __auxvar29__recorder_sn_condmet <= 1'b1; __auxvar29__recorder_sn_vhold <= __auxvar29__recorder_sn_value; end
       __auxvar2__recorder <= __auxvar2__recorder;
       if (__auxvar2__recorder_sn_cond ) begin __auxvar2__recorder_sn_condmet <= 1'b1; __auxvar2__recorder_sn_vhold <= __auxvar2__recorder_sn_value; end
       __auxvar30__recorder <= __auxvar30__recorder;
       if (__auxvar30__recorder_sn_cond ) begin __auxvar30__recorder_sn_condmet <= 1'b1; __auxvar30__recorder_sn_vhold <= __auxvar30__recorder_sn_value; end
       __auxvar31__recorder <= __auxvar31__recorder;
       if (__auxvar31__recorder_sn_cond ) begin __auxvar31__recorder_sn_condmet <= 1'b1; __auxvar31__recorder_sn_vhold <= __auxvar31__recorder_sn_value; end
       __auxvar32__recorder <= __auxvar32__recorder;
       if (__auxvar32__recorder_sn_cond ) begin __auxvar32__recorder_sn_condmet <= 1'b1; __auxvar32__recorder_sn_vhold <= __auxvar32__recorder_sn_value; end
       __auxvar33__recorder <= __auxvar33__recorder;
       if (__auxvar33__recorder_sn_cond ) begin __auxvar33__recorder_sn_condmet <= 1'b1; __auxvar33__recorder_sn_vhold <= __auxvar33__recorder_sn_value; end
       __auxvar34__recorder <= __auxvar34__recorder;
       if (__auxvar34__recorder_sn_cond ) begin __auxvar34__recorder_sn_condmet <= 1'b1; __auxvar34__recorder_sn_vhold <= __auxvar34__recorder_sn_value; end
       __auxvar35__recorder <= __auxvar35__recorder;
       if (__auxvar35__recorder_sn_cond ) begin __auxvar35__recorder_sn_condmet <= 1'b1; __auxvar35__recorder_sn_vhold <= __auxvar35__recorder_sn_value; end
       __auxvar36__recorder <= __auxvar36__recorder;
       if (__auxvar36__recorder_sn_cond ) begin __auxvar36__recorder_sn_condmet <= 1'b1; __auxvar36__recorder_sn_vhold <= __auxvar36__recorder_sn_value; end
       __auxvar37__recorder <= __auxvar37__recorder;
       if (__auxvar37__recorder_sn_cond ) begin __auxvar37__recorder_sn_condmet <= 1'b1; __auxvar37__recorder_sn_vhold <= __auxvar37__recorder_sn_value; end
       __auxvar38__recorder <= __auxvar38__recorder;
       if (__auxvar38__recorder_sn_cond ) begin __auxvar38__recorder_sn_condmet <= 1'b1; __auxvar38__recorder_sn_vhold <= __auxvar38__recorder_sn_value; end
       __auxvar3__recorder <= __auxvar3__recorder;
       if (__auxvar3__recorder_sn_cond ) begin __auxvar3__recorder_sn_condmet <= 1'b1; __auxvar3__recorder_sn_vhold <= __auxvar3__recorder_sn_value; end
       __auxvar4__recorder <= __auxvar4__recorder;
       if (__auxvar4__recorder_sn_cond ) begin __auxvar4__recorder_sn_condmet <= 1'b1; __auxvar4__recorder_sn_vhold <= __auxvar4__recorder_sn_value; end
       __auxvar5__recorder <= __auxvar5__recorder;
       if (__auxvar5__recorder_sn_cond ) begin __auxvar5__recorder_sn_condmet <= 1'b1; __auxvar5__recorder_sn_vhold <= __auxvar5__recorder_sn_value; end
       __auxvar6__recorder <= __auxvar6__recorder;
       if (__auxvar6__recorder_sn_cond ) begin __auxvar6__recorder_sn_condmet <= 1'b1; __auxvar6__recorder_sn_vhold <= __auxvar6__recorder_sn_value; end
       __auxvar7__recorder <= __auxvar7__recorder;
       if (__auxvar7__recorder_sn_cond ) begin __auxvar7__recorder_sn_condmet <= 1'b1; __auxvar7__recorder_sn_vhold <= __auxvar7__recorder_sn_value; end
       __auxvar8__recorder <= __auxvar8__recorder;
       if (__auxvar8__recorder_sn_cond ) begin __auxvar8__recorder_sn_condmet <= 1'b1; __auxvar8__recorder_sn_vhold <= __auxvar8__recorder_sn_value; end
       __auxvar9__recorder <= __auxvar9__recorder;
       if (__auxvar9__recorder_sn_cond ) begin __auxvar9__recorder_sn_condmet <= 1'b1; __auxvar9__recorder_sn_vhold <= __auxvar9__recorder_sn_value; end
       __auxvar0__delay_d_1 <= __auxvar0__delay_d_0 ;
       if(monitor_s1_already_enter_cond) begin monitor_s1_already <= 1'b1;
       end
       else if(monitor_s1_already_exit_cond) begin monitor_s1_already <= 1'b0;
       end
       if(monitor_s2_enter_cond) begin monitor_s2 <= 1'b1;
       end
       else if(monitor_s2_exit_cond) begin monitor_s2 <= 1'b0;
       end
       if(monitor_s3_enter_cond) begin monitor_s3 <= 1'b1;
       end
       else if(monitor_s3_exit_cond) begin monitor_s3 <= 1'b0;
       end
       if(monitor_s4_enter_cond) begin monitor_s4 <= 1'b1;
       end
       else if(monitor_s4_exit_cond) begin monitor_s4 <= 1'b0;
       end
   end
end
endmodule