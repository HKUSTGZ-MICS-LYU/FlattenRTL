module dma_axi64_core0_top #(
        parameter dma_axi64_core0_dma_axi64_core0_arbiter_rd_CH_LAST=1-1,
        parameter dma_axi64_core0_dma_axi64_core0_arbiter_wr_CH_LAST=1-1,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE=3'd0,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD=3'd1,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_CLR=3'd2,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY=3'd3,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL=3'd4,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE=3'd0,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD=3'd1,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_CLR=3'd2,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY=3'd3,
        parameter dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL=3'd4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AXI_WORD_SIZE=0?2'b10:2'b11,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AXI_3=0?2:3,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_SIZE_BITS=4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_DELAY=2,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_DELAY=2,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_SIZE_BITS,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL=2,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH=7+4+2+1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_FULL=4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH=8+4+7+2,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_FULL=4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH=64,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_FULL=5+2,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_DEPTH=3,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_CMD_DEPTH=4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP_SLVERR=2'b10,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP_DECERR=2'b11,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH=7,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_FULL=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_CMD_DEPTH,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AXI_WORD_SIZE=0?2'b10:2'b11,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AXI_3=0?2:3,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_CMD_DEPTH=4,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP_SLVERR=2'b10,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP_DECERR=2'b11,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH=7,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_FULL=dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_CMD_DEPTH,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_SINGLE=dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_FULL==1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH=dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_SINGLE?1:dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_FULL-1,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_BITS=(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=2)?1:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=4)?2:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=8)?3:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=16)?4:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=32)?5:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=64)?6:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=128)?7:(dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH<=256)?8:0,
        parameter dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_LAST_LINE=dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH-1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH=32,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH=64,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH=31,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH=31,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH=3,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH=3,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH=32,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH=6,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH=6,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH=32,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT=0?32:0,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE0=8'h00,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE1=8'h04,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE2=8'h08,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE3=8'h0C,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE0=8'h10,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE1=8'h14,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE2=8'h18,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE3=8'h1C,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE4=8'h20,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RESTRICT=8'h2C,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RD_OFFSETS=8'h30,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_WR_OFFSETS=8'h34,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_FIFO_FULLNESS=8'h38,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_OUTS=8'h3C,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ENABLE=8'h40,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_START=8'h44,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ACTIVE=8'h48,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_CMD_COUNTER=8'h50,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_RAWSTAT=8'hA0,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_CLEAR=8'hA4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_ENABLE=8'hA8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_STATUS=8'hAC,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST=0?64:128,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES=32/2,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_LARGE_FIFO=32>dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_SMALL_FIFO=32==16,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_MAX_BURST=0?64:128,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES=32/2,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_LARGE_FIFO=32>dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_SMALL_FIFO=32==16,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE=13,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_READ=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_SINGLE_SIZE=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_READ=0,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_SINGLE_SIZE=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_READ=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_CMD_SIZE=16,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_READ=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_CMD_SIZE=16,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH=8,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE=!dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE=3'd0,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE=3'd1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT=3'd2,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY=3'd3,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS=3'd4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ=3'd5,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK=3'd6,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH=3'd7,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ=dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE=!dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE=3'd0,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE=3'd1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT=3'd2,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY=3'd3,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS=3'd4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ=3'd5,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK=3'd6,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH=3'd7,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_WIDTH=4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_WIDTH=4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_DELAY=2,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_DELAY=1,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_WIDTH=4,
        parameter dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_DELAY=1) (
            input clk,
            input reset,
            input scan_en,
            output idle,
            output [8*1-1:0] ch_int_all_proc,
            input [7:0] ch_start,
            input [3:0] clkdiv,
            input [31:1] periph_tx_req,
            output [31:1] periph_tx_clr,
            input [31:1] periph_rx_req,
            output [31:1] periph_rx_clr,
            input pclken,
            input psel,
            input penable,
            input [10:0] paddr,
            input pwrite,
            input [31:0] pwdata,
            output [31:0] prdata,
            output pslverr,
            output pready,
            output rd_port_num,
            output wr_port_num,
            input joint_mode,
            input joint_remote,
            input rd_prio_top,
            input rd_prio_high,
            input [2:0] rd_prio_top_num,
            input [2:0] rd_prio_high_num,
            input wr_prio_top,
            input wr_prio_high,
            input [2:0] wr_prio_top_num,
            input [2:0] wr_prio_high_num,
            output [31:0] AWADDR,
            output [4-1:0] AWLEN,
            output [2-1:0] AWSIZE,
            output AWVALID,
            input AWREADY,
            output [63:0] WDATA,
            output [64/8-1:0] WSTRB,
            output WLAST,
            output WVALID,
            input WREADY,
            input [1:0] BRESP,
            input BVALID,
            output BREADY,
            output [31:0] ARADDR,
            output [4-1:0] ARLEN,
            output [2-1:0] ARSIZE,
            output ARVALID,
            input ARREADY,
            input [63:0] RDATA,
            input [1:0] RRESP,
            input RLAST,
            input RVALID,
            output RREADY) ;
    wire [31:0] slow_AWADDR ;
    wire [4-1:0] slow_AWLEN ;
    wire [2-1:0] slow_AWSIZE ;
    wire slow_AWVALID ;
    wire slow_AWREADY ;
    wire [63:0] slow_WDATA ;
    wire [64/8-1:0] slow_WSTRB ;
    wire slow_WLAST ;
    wire slow_WVALID ;
    wire slow_WREADY ;
    wire [1:0] slow_BRESP ;
    wire slow_BVALID ;
    wire slow_BREADY ;
    wire [31:0] slow_ARADDR ;
    wire [4-1:0] slow_ARLEN ;
    wire [2-1:0] slow_ARSIZE ;
    wire slow_ARVALID ;
    wire slow_ARREADY ;
    wire [63:0] slow_RDATA ;
    wire [1:0] slow_RRESP ;
    wire slow_RLAST ;
    wire slow_RVALID ;
    wire slow_RREADY ;
    wire clk_out ;
    wire clken ;
    wire bypass ;
    assign clk_out=clk;
    assign clken=1'b1;
    assign AWADDR=slow_AWADDR;
    assign AWLEN=slow_AWLEN;
    assign AWSIZE=slow_AWSIZE;
    assign AWVALID=slow_AWVALID;
    assign WDATA=slow_WDATA;
    assign WSTRB=slow_WSTRB;
    assign WLAST=slow_WLAST;
    assign WVALID=slow_WVALID;
    assign BREADY=slow_BREADY;
    assign ARADDR=slow_ARADDR;
    assign ARLEN=slow_ARLEN;
    assign ARSIZE=slow_ARSIZE;
    assign ARVALID=slow_ARVALID;
    assign RREADY=slow_RREADY;
    assign slow_AWREADY=AWREADY;
    assign slow_WREADY=WREADY;
    assign slow_BRESP=BRESP;
    assign slow_BVALID=BVALID;
    assign slow_ARREADY=ARREADY;
    assign slow_RDATA=RDATA;
    assign slow_RRESP=RRESP;
    assign slow_RLAST=RLAST;
    assign slow_RVALID=RVALID;

    wire  dma_axi64_core0_clk;
    wire  dma_axi64_core0_reset;
    wire  dma_axi64_core0_scan_en;
    wire  dma_axi64_core0_idle;
    wire [8*1-1:0] dma_axi64_core0_ch_int_all_proc;
    wire [7:0] dma_axi64_core0_ch_start;
    wire [31:1] dma_axi64_core0_periph_tx_req;
    wire [31:1] dma_axi64_core0_periph_tx_clr;
    wire [31:1] dma_axi64_core0_periph_rx_req;
    wire [31:1] dma_axi64_core0_periph_rx_clr;
    wire  dma_axi64_core0_pclk;
    wire  dma_axi64_core0_clken;
    wire  dma_axi64_core0_pclken;
    wire  dma_axi64_core0_psel;
    wire  dma_axi64_core0_penable;
    wire [10:0] dma_axi64_core0_paddr;
    wire  dma_axi64_core0_pwrite;
    wire [31:0] dma_axi64_core0_pwdata;
    wire [31:0] dma_axi64_core0_prdata;
    wire  dma_axi64_core0_pslverr;
    wire  dma_axi64_core0_rd_port_num;
    wire  dma_axi64_core0_wr_port_num;
    wire  dma_axi64_core0_joint_mode_in;
    wire  dma_axi64_core0_joint_remote;
    wire  dma_axi64_core0_rd_prio_top;
    wire  dma_axi64_core0_rd_prio_high;
    wire [2:0] dma_axi64_core0_rd_prio_top_num;
    wire [2:0] dma_axi64_core0_rd_prio_high_num;
    wire  dma_axi64_core0_wr_prio_top;
    wire  dma_axi64_core0_wr_prio_high;
    wire [2:0] dma_axi64_core0_wr_prio_top_num;
    wire [2:0] dma_axi64_core0_wr_prio_high_num;
    wire [31:0] dma_axi64_core0_AWADDR;
    wire [4-1:0] dma_axi64_core0_AWLEN;
    wire [2-1:0] dma_axi64_core0_AWSIZE;
    wire  dma_axi64_core0_AWVALID;
    wire  dma_axi64_core0_AWREADY;
    wire [63:0] dma_axi64_core0_WDATA;
    wire [64/8-1:0] dma_axi64_core0_WSTRB;
    wire  dma_axi64_core0_WLAST;
    wire  dma_axi64_core0_WVALID;
    wire  dma_axi64_core0_WREADY;
    wire [1:0] dma_axi64_core0_BRESP;
    wire  dma_axi64_core0_BVALID;
    wire  dma_axi64_core0_BREADY;
    wire [31:0] dma_axi64_core0_ARADDR;
    wire [4-1:0] dma_axi64_core0_ARLEN;
    wire [2-1:0] dma_axi64_core0_ARSIZE;
    wire  dma_axi64_core0_ARVALID;
    wire  dma_axi64_core0_ARREADY;
    wire [63:0] dma_axi64_core0_RDATA;
    wire [1:0] dma_axi64_core0_RRESP;
    wire  dma_axi64_core0_RLAST;
    wire  dma_axi64_core0_RVALID;
    wire  dma_axi64_core0_RREADY;

    wire  dma_axi64_core0_wdt_timeout  ;
    wire[2:0]  dma_axi64_core0_wdt_ch_num  ;
    wire  dma_axi64_core0_rd_ch_go_joint  ;
    wire  dma_axi64_core0_rd_ch_go_null  ;
    wire  dma_axi64_core0_rd_ch_go  ;
    wire[2:0]  dma_axi64_core0_rd_ch_num  ;
    wire  dma_axi64_core0_rd_ch_last  ;
    wire  dma_axi64_core0_wr_ch_go_joint  ;
    wire  dma_axi64_core0_wr_ch_go  ;
    wire[2:0]  dma_axi64_core0_wr_ch_num_joint  ;
    wire[2:0]  dma_axi64_core0_wr_ch_num  ;
    wire  dma_axi64_core0_wr_ch_last  ;
    wire  dma_axi64_core0_wr_ch_last_joint  ;
    wire  dma_axi64_core0_load_req_in_prog  ;
    wire[7:0]  dma_axi64_core0_ch_idle  ;
    wire[7:0]  dma_axi64_core0_ch_active  ;
    wire[7:0]  dma_axi64_core0_ch_active_joint  ;
    wire[7:0]  dma_axi64_core0_ch_rd_active  ;
    wire[7:0]  dma_axi64_core0_ch_wr_active  ;
    wire  dma_axi64_core0_wr_last_cmd  ;
    wire  dma_axi64_core0_rd_line_cmd  ;
    wire  dma_axi64_core0_wr_line_cmd  ;
    wire  dma_axi64_core0_rd_go_next_line  ;
    wire  dma_axi64_core0_wr_go_next_line  ;
    wire[7:0]  dma_axi64_core0_ch_rd_ready_joint  ;
    wire[7:0]  dma_axi64_core0_ch_rd_ready  ;
    wire  dma_axi64_core0_rd_ready  ;
    wire  dma_axi64_core0_rd_ready_joint  ;
    wire[32-1:0]  dma_axi64_core0_rd_burst_addr  ;
    wire[8-1:0]  dma_axi64_core0_rd_burst_size  ;
    wire[6-1:0]  dma_axi64_core0_rd_tokens  ;
    wire[3-1:0]  dma_axi64_core0_rd_periph_delay  ;
    wire  dma_axi64_core0_rd_clr_valid  ;
    wire[2:0]  dma_axi64_core0_rd_transfer_num  ;
    wire  dma_axi64_core0_rd_transfer  ;
    wire[4-1:0]  dma_axi64_core0_rd_transfer_size  ;
    wire  dma_axi64_core0_rd_clr_stall  ;
    wire[7:0]  dma_axi64_core0_ch_wr_ready  ;
    wire  dma_axi64_core0_wr_ready  ;
    wire  dma_axi64_core0_wr_ready_joint  ;
    wire[32-1:0]  dma_axi64_core0_wr_burst_addr  ;
    wire[8-1:0]  dma_axi64_core0_wr_burst_size  ;
    wire[6-1:0]  dma_axi64_core0_wr_tokens  ;
    wire[3-1:0]  dma_axi64_core0_wr_periph_delay  ;
    wire  dma_axi64_core0_wr_clr_valid  ;
    wire  dma_axi64_core0_wr_clr_stall  ;
    wire[7:0]  dma_axi64_core0_ch_joint_req  ;
    wire  dma_axi64_core0_joint_req  ;
    wire  dma_axi64_core0_joint_mode  ;
    wire  dma_axi64_core0_joint_ch_go  ;
    wire  dma_axi64_core0_joint_stall  ;
    wire  dma_axi64_core0_rd_burst_start  ;
    wire  dma_axi64_core0_rd_finish_joint  ;
    wire  dma_axi64_core0_rd_finish  ;
    wire  dma_axi64_core0_rd_ctrl_busy  ;
    wire  dma_axi64_core0_wr_burst_start_joint  ;
    wire  dma_axi64_core0_wr_burst_start  ;
    wire  dma_axi64_core0_wr_finish  ;
    wire  dma_axi64_core0_wr_ctrl_busy  ;
    wire  dma_axi64_core0_wr_cmd_split  ;
    wire[2:0]  dma_axi64_core0_wr_cmd_num  ;
    wire  dma_axi64_core0_wr_cmd_pending_joint  ;
    wire  dma_axi64_core0_wr_cmd_pending  ;
    wire  dma_axi64_core0_wr_cmd_full_joint  ;
    wire  dma_axi64_core0_ch_fifo_rd  ;
    wire[4-1:0]  dma_axi64_core0_ch_fifo_rsize  ;
    wire[2:0]  dma_axi64_core0_ch_fifo_rd_num  ;
    wire[2:0]  dma_axi64_core0_wr_transfer_num  ;
    wire  dma_axi64_core0_wr_transfer  ;
    wire[4-1:0]  dma_axi64_core0_wr_transfer_size  ;
    wire[4-1:0]  dma_axi64_core0_wr_next_size  ;
    wire  dma_axi64_core0_wr_clr_line  ;
    wire[2:0]  dma_axi64_core0_wr_clr_line_num  ;
    wire  dma_axi64_core0_wr_cmd_full  ;
    wire  dma_axi64_core0_wr_slverr  ;
    wire  dma_axi64_core0_wr_decerr  ;
    wire  dma_axi64_core0_wr_clr  ;
    wire  dma_axi64_core0_wr_clr_last  ;
    wire[2:0]  dma_axi64_core0_wr_ch_num_resp  ;
    wire  dma_axi64_core0_timeout_aw  ;
    wire  dma_axi64_core0_timeout_w  ;
    wire[2:0]  dma_axi64_core0_timeout_num_aw  ;
    wire[2:0]  dma_axi64_core0_timeout_num_w  ;
    wire  dma_axi64_core0_wr_hold_ctrl  ;
    wire  dma_axi64_core0_wr_hold  ;
    wire  dma_axi64_core0_joint_in_prog  ;
    wire  dma_axi64_core0_joint_not_in_prog  ;
    wire  dma_axi64_core0_joint_mux_in_prog  ;
    wire  dma_axi64_core0_wr_page_cross  ;
    wire  dma_axi64_core0_load_wr  ;
    wire[2:0]  dma_axi64_core0_load_wr_num  ;
    wire[1:0]  dma_axi64_core0_load_wr_cycle  ;
    wire[64-1:0]  dma_axi64_core0_load_wdata  ;
    wire  dma_axi64_core0_rd_cmd_split  ;
    wire  dma_axi64_core0_rd_cmd_line  ;
    wire[2:0]  dma_axi64_core0_rd_cmd_num  ;
    wire  dma_axi64_core0_rd_cmd_pending_joint  ;
    wire  dma_axi64_core0_rd_cmd_pending  ;
    wire  dma_axi64_core0_rd_cmd_full_joint  ;
    wire  dma_axi64_core0_ch_fifo_wr  ;
    wire[64-1:0]  dma_axi64_core0_ch_fifo_wdata  ;
    wire[4-1:0]  dma_axi64_core0_ch_fifo_wsize  ;
    wire[2:0]  dma_axi64_core0_ch_fifo_wr_num  ;
    wire  dma_axi64_core0_rd_clr_line  ;
    wire[2:0]  dma_axi64_core0_rd_clr_line_num  ;
    wire  dma_axi64_core0_rd_burst_cmd  ;
    wire  dma_axi64_core0_rd_cmd_full  ;
    wire  dma_axi64_core0_rd_slverr  ;
    wire  dma_axi64_core0_rd_decerr  ;
    wire  dma_axi64_core0_rd_clr  ;
    wire  dma_axi64_core0_rd_clr_last  ;
    wire  dma_axi64_core0_rd_clr_load  ;
    wire[2:0]  dma_axi64_core0_rd_ch_num_resp  ;
    wire  dma_axi64_core0_timeout_ar  ;
    wire[2:0]  dma_axi64_core0_timeout_num_ar  ;
    wire  dma_axi64_core0_rd_hold_joint  ;
    wire  dma_axi64_core0_rd_hold_ctrl  ;
    wire  dma_axi64_core0_rd_hold  ;
    wire  dma_axi64_core0_joint_hold  ;
    wire  dma_axi64_core0_rd_page_cross  ;
    wire  dma_axi64_core0_joint_page_cross  ;
    wire  dma_axi64_core0_rd_arbiter_en  ;
    wire  dma_axi64_core0_wr_arbiter_en  ;
    wire  dma_axi64_core0_rd_cmd_port  ;
    wire  dma_axi64_core0_wr_cmd_port  ;
    wire[64-1:0]  dma_axi64_core0_ch_fifo_rdata  ;
    wire  dma_axi64_core0_ch_fifo_rd_valid  ;
    wire  dma_axi64_core0_ch_fifo_wr_ready  ;
    wire  dma_axi64_core0_FIFO_WR  ;
    wire  dma_axi64_core0_FIFO_RD  ;
    wire[3+5-3-1:0]  dma_axi64_core0_FIFO_WR_ADDR  ;
    wire[3+5-3-1:0]  dma_axi64_core0_FIFO_RD_ADDR  ;
    wire[64-1:0]  dma_axi64_core0_FIFO_DIN  ;
    wire[8-1:0]  dma_axi64_core0_FIFO_BSEL  ;
    wire[64-1:0]  dma_axi64_core0_FIFO_DOUT  ;
    wire  dma_axi64_core0_clk_en  ;
    wire  dma_axi64_core0_gclk  ;
    assign   dma_axi64_core0_joint_mode  =  dma_axi64_core0_joint_mode_in  &1'b1;
    assign   dma_axi64_core0_rd_arbiter_en  =1'b1;
    assign   dma_axi64_core0_wr_arbiter_en  =!  dma_axi64_core0_joint_mode  ;
    assign   dma_axi64_core0_rd_ready  =  dma_axi64_core0_ch_rd_ready  [  dma_axi64_core0_rd_ch_num  ];
    assign   dma_axi64_core0_wr_ready  =  dma_axi64_core0_ch_wr_ready  [  dma_axi64_core0_wr_ch_num_joint  ];
    assign   dma_axi64_core0_rd_ready_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_rd_ready  &  dma_axi64_core0_wr_ready  :  dma_axi64_core0_rd_ready  ;
    assign   dma_axi64_core0_wr_ready_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_rd_ready  &  dma_axi64_core0_wr_ready  :  dma_axi64_core0_wr_ready  ;
    assign   dma_axi64_core0_ch_active_joint  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_ch_rd_active  |  dma_axi64_core0_ch_wr_active  :  dma_axi64_core0_ch_rd_active  ;
    assign   dma_axi64_core0_joint_page_cross  =(  dma_axi64_core0_rd_page_cross  &  dma_axi64_core0_rd_ready  )|(  dma_axi64_core0_wr_page_cross  &  dma_axi64_core0_wr_ready  );
    assign   dma_axi64_core0_joint_req  =  dma_axi64_core0_ch_joint_req  [  dma_axi64_core0_rd_ch_num  ];
    assign   dma_axi64_core0_ch_rd_ready_joint  =  dma_axi64_core0_joint_mode   ? (  dma_axi64_core0_ch_joint_req  &  dma_axi64_core0_ch_rd_ready  &  dma_axi64_core0_ch_wr_ready  )|((~  dma_axi64_core0_ch_joint_req  )&(  dma_axi64_core0_ch_rd_ready  |  dma_axi64_core0_ch_wr_ready  )):  dma_axi64_core0_ch_rd_ready  ;
    assign   dma_axi64_core0_wr_burst_start_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_rd_burst_start  :  dma_axi64_core0_wr_burst_start  ;
    assign   dma_axi64_core0_joint_hold  =  dma_axi64_core0_joint_mux_in_prog  |(  dma_axi64_core0_joint_in_prog  &(~  dma_axi64_core0_joint_req  ))|(  dma_axi64_core0_joint_not_in_prog  &  dma_axi64_core0_joint_req  )|  dma_axi64_core0_joint_stall  |(  dma_axi64_core0_joint_req  &  dma_axi64_core0_joint_page_cross  );
    assign   dma_axi64_core0_rd_hold_ctrl  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_rd_hold  |  dma_axi64_core0_joint_hold  |(  dma_axi64_core0_joint_in_prog  &  dma_axi64_core0_wr_hold  ):  dma_axi64_core0_rd_hold  ;
    assign   dma_axi64_core0_rd_hold_joint  =  dma_axi64_core0_joint_mode  &(  dma_axi64_core0_rd_hold_ctrl  |  dma_axi64_core0_rd_ctrl_busy  |  dma_axi64_core0_wr_ctrl_busy  );
    assign   dma_axi64_core0_wr_hold_ctrl  =  dma_axi64_core0_joint_mode  &(  dma_axi64_core0_joint_req  |  dma_axi64_core0_joint_in_prog  ) ?   dma_axi64_core0_wr_hold  |  dma_axi64_core0_joint_hold  :  dma_axi64_core0_wr_hold  ;
    assign   dma_axi64_core0_rd_ch_go_joint  =  dma_axi64_core0_rd_ch_go  &  dma_axi64_core0_ch_rd_ready  [  dma_axi64_core0_rd_ch_num  ]&(~  dma_axi64_core0_rd_ctrl_busy  );
    assign   dma_axi64_core0_wr_ch_go_joint  =  dma_axi64_core0_joint_mode   ? (  dma_axi64_core0_wr_ready  &(~  dma_axi64_core0_wr_ctrl_busy  )&(  dma_axi64_core0_joint_req   ?   dma_axi64_core0_rd_ch_go_joint  :  dma_axi64_core0_rd_ch_go  &(~  dma_axi64_core0_rd_ch_go_joint  ))):  dma_axi64_core0_wr_ch_go  ;
    assign   dma_axi64_core0_rd_ch_go_null  =  dma_axi64_core0_rd_ch_go  &(~  dma_axi64_core0_rd_ch_go_joint  )&(  dma_axi64_core0_joint_mode   ? (~  dma_axi64_core0_wr_ch_go_joint  ):1'b1);
    assign   dma_axi64_core0_wr_ch_num_joint  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_rd_ch_num  :  dma_axi64_core0_wr_ch_num  ;
    assign   dma_axi64_core0_wr_ch_last_joint  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_rd_ch_last  :  dma_axi64_core0_wr_ch_last  ;
    assign   dma_axi64_core0_rd_finish_joint  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_rd_finish  |  dma_axi64_core0_wr_finish  |  dma_axi64_core0_rd_ch_go_null  :  dma_axi64_core0_rd_finish  |  dma_axi64_core0_rd_ch_go_null  ;
    assign   dma_axi64_core0_rd_cmd_full_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_wr_cmd_full  |  dma_axi64_core0_rd_cmd_full  :  dma_axi64_core0_rd_cmd_full  ;
    assign   dma_axi64_core0_wr_cmd_full_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_wr_cmd_full  |  dma_axi64_core0_rd_cmd_full  :  dma_axi64_core0_wr_cmd_full  ;
    assign   dma_axi64_core0_rd_cmd_pending_joint  =  dma_axi64_core0_joint_mode   ?   dma_axi64_core0_rd_cmd_pending  |  dma_axi64_core0_wr_cmd_pending  :  dma_axi64_core0_rd_cmd_pending  ;
    assign   dma_axi64_core0_wr_cmd_pending_joint  =  dma_axi64_core0_joint_mode  &  dma_axi64_core0_joint_req   ?   dma_axi64_core0_rd_cmd_pending  |  dma_axi64_core0_wr_cmd_pending  :  dma_axi64_core0_wr_cmd_pending  ;
    assign   dma_axi64_core0_idle  =&  dma_axi64_core0_ch_idle  ;
    assign   dma_axi64_core0_gclk  =  dma_axi64_core0_clk  ;

    wire  dma_axi64_core0_dma_axi64_core0_wdt_clk;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_reset;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_wdt_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_rd_burst_start;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_wdt_rd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_wr_burst_start;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_wdt_wr_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_wdt_timeout;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num;

    reg[11-1:0]  dma_axi64_core0_dma_axi64_core0_wdt_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_current_ch_active  ;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_current_burst_start  ;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_advance  ;
    wire  dma_axi64_core0_dma_axi64_core0_wdt_idle  ;
    assign   dma_axi64_core0_dma_axi64_core0_wdt_idle  =  dma_axi64_core0_dma_axi64_core0_wdt_ch_active  ==8'd0;
    assign   dma_axi64_core0_dma_axi64_core0_wdt_current_ch_active  =  dma_axi64_core0_dma_axi64_core0_wdt_ch_active  [  dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num  ];
    assign   dma_axi64_core0_dma_axi64_core0_wdt_current_burst_start  =(  dma_axi64_core0_dma_axi64_core0_wdt_rd_burst_start  &(  dma_axi64_core0_dma_axi64_core0_wdt_rd_ch_num  ==  dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num  ))|(  dma_axi64_core0_dma_axi64_core0_wdt_wr_burst_start  &(  dma_axi64_core0_dma_axi64_core0_wdt_wr_ch_num  ==  dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num  ));
    assign   dma_axi64_core0_dma_axi64_core0_wdt_advance  =(!  dma_axi64_core0_dma_axi64_core0_wdt_current_ch_active  )|  dma_axi64_core0_dma_axi64_core0_wdt_current_burst_start  |  dma_axi64_core0_dma_axi64_core0_wdt_wdt_timeout  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_wdt_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_wdt_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_wdt_reset  )
            dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num   <=3'd0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_wdt_advance  )
                dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num   <=  dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num  +1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_wdt_wdt_timeout  =(  dma_axi64_core0_dma_axi64_core0_wdt_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_wdt_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_wdt_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_wdt_reset  )
            dma_axi64_core0_dma_axi64_core0_wdt_counter   <={11{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_wdt_advance  |  dma_axi64_core0_dma_axi64_core0_wdt_idle  )
                dma_axi64_core0_dma_axi64_core0_wdt_counter   <={11{1'b1}};
            else
                dma_axi64_core0_dma_axi64_core0_wdt_counter   <=  dma_axi64_core0_dma_axi64_core0_wdt_counter  -1'b1;

    assign dma_axi64_core0_dma_axi64_core0_wdt_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_wdt_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_wdt_ch_active = dma_axi64_core0_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_wdt_rd_burst_start = dma_axi64_core0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_wdt_rd_ch_num = dma_axi64_core0_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_wdt_wr_burst_start = dma_axi64_core0_wr_burst_start_joint;
    assign dma_axi64_core0_dma_axi64_core0_wdt_wr_ch_num = dma_axi64_core0_wr_ch_num_joint;
    assign dma_axi64_core0_wdt_timeout = dma_axi64_core0_dma_axi64_core0_wdt_wdt_timeout;
    assign dma_axi64_core0_wdt_ch_num = dma_axi64_core0_dma_axi64_core0_wdt_wdt_ch_num;


    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_enable;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_top;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_high;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_top_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_high_num;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_hold;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_ready;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_finish;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_out;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_last;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_enable;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_top;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_high;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_top_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_high_num;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_hold;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_ready;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_finish;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_out;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_last;

    reg[7:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_current_active  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_current_ready_only  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_last_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ready0  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ready1  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_top_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_high_ready  ;
    reg  dma_axi64_core0_dma_axi64_core0_arbiter_rd_in_prog  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_pre_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_top_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_high_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_top  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_high  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_next  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_hold_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_rd_advance_next  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_num_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num0_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num0_pre2  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num0  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num1_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num1_pre2  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num1  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_rd_next_ch_num_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_out  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_last  ='d1;



    reg[7:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_current_active  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_current_ready_only  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_last_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ready0  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ready1  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_top_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_high_ready  ;
    reg  dma_axi64_core0_dma_axi64_core0_arbiter_wr_in_prog  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_pre_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_top_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_high_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_top  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_high  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_next  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_hold_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_arbiter_wr_advance_next  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_num_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num0_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num0_pre2  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num0  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num1_pre  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num1_pre2  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num1  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_arbiter_wr_next_ch_num_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_out  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_last  ='d1;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_enable = dma_axi64_core0_rd_arbiter_en;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_joint_mode = dma_axi64_core0_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_page_cross = dma_axi64_core0_joint_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_top = dma_axi64_core0_rd_prio_top;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_high = dma_axi64_core0_rd_prio_high;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_top_num = dma_axi64_core0_rd_prio_top_num;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_prio_high_num = dma_axi64_core0_rd_prio_high_num;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_hold = dma_axi64_core0_rd_hold_joint;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_ready = dma_axi64_core0_ch_rd_ready_joint;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_active = dma_axi64_core0_ch_active_joint;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_rd_finish = dma_axi64_core0_rd_finish_joint;
    assign dma_axi64_core0_rd_ch_go = dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_go_out;
    assign dma_axi64_core0_rd_ch_num = dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_num;
    assign dma_axi64_core0_rd_ch_last = dma_axi64_core0_dma_axi64_core0_arbiter_rd_ch_last;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_enable = dma_axi64_core0_wr_arbiter_en;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_joint_mode = dma_axi64_core0_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_page_cross = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_top = dma_axi64_core0_wr_prio_top;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_high = dma_axi64_core0_wr_prio_high;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_top_num = dma_axi64_core0_wr_prio_top_num;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_prio_high_num = dma_axi64_core0_wr_prio_high_num;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_hold = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_ready = dma_axi64_core0_ch_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_active = dma_axi64_core0_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_arbiter_wr_finish = dma_axi64_core0_wr_finish;
    assign dma_axi64_core0_wr_ch_go = dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_go_out;
    assign dma_axi64_core0_wr_ch_num = dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_num;
    assign dma_axi64_core0_wr_ch_last = dma_axi64_core0_dma_axi64_core0_arbiter_wr_ch_last;


    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_req;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_clr_stall;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_rd_burst_start;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_busy;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_hold;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_req;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_clr_stall;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_wr_burst_start;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_busy;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_hold;

    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  ;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain_reg  ;
    reg[6-1:0]  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall  ;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_ch  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last_ch  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line_d  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_busy  =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps  !=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_ch  =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid  &  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr  &(  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num  ==  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num_resp  );
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last_ch  =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid  &  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last  &(  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num  ==  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num_resp  );
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line_d  =1'b0;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish  )
                dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl_reg   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl_reg   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_req  ;

    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl  =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  =(|  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter  )|  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter   <={6{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go  )
                dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_burst_start  &(|  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter  ))
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_counter  -1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter   <={3{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_ch  )
                dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_delay  ;
            else
                if (|  dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter  -1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall  =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_pending  |  dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_full  |  dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line_d  ;
    always @(                  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go                                        or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last                        or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready                       or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_clr_stall                      or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter                     or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line_d                    or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_hold                   or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl                  or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_req                 or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_ch                or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last_ch               or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid              or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_delay             or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps            or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall           or    dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain   )
    begin
        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
        dma_axi64_core0_dma_axi64_core0_ctrl_rd_burst_start   =1'b0;
        dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b0;
        case (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps  )
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go  )
                begin
                    if (!  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                    end
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall  )
                            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL  ;
                        else
                            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD  ;
                end
                else
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_req  ^  dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_ctrl  )
                begin
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                end
                else
                    if ((  dma_axi64_core0_dma_axi64_core0_ctrl_rd_clr_stall  |  dma_axi64_core0_dma_axi64_core0_ctrl_rd_hold  )&  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  )
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready  &  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  )
                        begin
                            if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall  )
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL  ;
                            else
                            begin
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_burst_start   =1'b1;
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_CLR  ;
                            end
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last  &(~  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready  ))
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD  ;
                            else
                            begin
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                                dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                            end
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_CLR   :
            begin
                if ((|  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_delay  )&  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid  )
                begin
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last_ch  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                    end
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_ch  )
                            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY  ;
                        else
                            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_CLR  ;
                end
                else
                    if (!  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                    end
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line_d  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_delay_counter  =='d0)
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_WAIT_DELAY  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready  &  dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens_remain  )
                begin
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_stall  )
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_STALL  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD  ;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last  &(~  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready  ))
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_CMD  ;
                    else
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish   =1'b1;
                    end
            end
            default :
            begin
                dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
            end
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_IDLE  ;
        else
            dma_axi64_core0_dma_axi64_core0_ctrl_rd_ps   <=  dma_axi64_core0_dma_axi64_core0_ctrl_rd_ns  ;




    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  ;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain_reg  ;
    reg[6-1:0]  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall  ;
    reg  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_ch  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last_ch  ;
    wire  dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line_d  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_busy  =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps  !=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_ch  =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid  &  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr  &(  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num  ==  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num_resp  );
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last_ch  =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid  &  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last  &(  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num  ==  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num_resp  );
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line_d  =1'b0;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish  )
                dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl_reg   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl_reg   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_req  ;

    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl  =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  =(|  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter  )|  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter   <={6{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go  )
                dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_burst_start  &(|  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter  ))
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_counter  -1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter   <={3{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_ch  )
                dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_delay  ;
            else
                if (|  dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter  -1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall  =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_pending  |  dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_full  |  dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line_d  ;
    always @(                  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go                                        or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last                        or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready                       or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_clr_stall                      or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter                     or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line_d                    or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_hold                   or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl                  or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_req                 or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_ch                or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last_ch               or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid              or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_delay             or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps            or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall           or    dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain   )
    begin
        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
        dma_axi64_core0_dma_axi64_core0_ctrl_wr_burst_start   =1'b0;
        dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b0;
        case (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps  )
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go  )
                begin
                    if (!  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                    end
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall  )
                            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL  ;
                        else
                            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD  ;
                end
                else
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_req  ^  dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_ctrl  )
                begin
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                end
                else
                    if ((  dma_axi64_core0_dma_axi64_core0_ctrl_wr_clr_stall  |  dma_axi64_core0_dma_axi64_core0_ctrl_wr_hold  )&  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  )
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready  &  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  )
                        begin
                            if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall  )
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL  ;
                            else
                            begin
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_burst_start   =1'b1;
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_CLR  ;
                            end
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last  &(~  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready  ))
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD  ;
                            else
                            begin
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                                dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                            end
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_CLR   :
            begin
                if ((|  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_delay  )&  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid  )
                begin
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last_ch  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                    end
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_ch  )
                            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY  ;
                        else
                            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_CLR  ;
                end
                else
                    if (!  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                    end
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line_d  )
                    dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_delay_counter  =='d0)
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_WAIT_DELAY  ;
            end
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready  &  dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens_remain  )
                begin
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_stall  )
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_STALL  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD  ;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last  &(~  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready  ))
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_CMD  ;
                    else
                    begin
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish   =1'b1;
                    end
            end
            default :
            begin
                dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns   =  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
            end
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_IDLE  ;
        else
            dma_axi64_core0_dma_axi64_core0_ctrl_wr_ps   <=  dma_axi64_core0_dma_axi64_core0_ctrl_wr_ns  ;

    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_go = dma_axi64_core0_rd_ch_go_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_full = dma_axi64_core0_rd_cmd_full_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_cmd_pending = dma_axi64_core0_rd_cmd_pending_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num = dma_axi64_core0_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_num_resp = dma_axi64_core0_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_go_next_line = dma_axi64_core0_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_valid = dma_axi64_core0_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr = dma_axi64_core0_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_clr_last = dma_axi64_core0_rd_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_periph_delay = dma_axi64_core0_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_clr_stall = dma_axi64_core0_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_tokens = dma_axi64_core0_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_ready = dma_axi64_core0_rd_ready_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_ch_last = dma_axi64_core0_rd_ch_last;
    assign dma_axi64_core0_rd_burst_start = dma_axi64_core0_dma_axi64_core0_ctrl_rd_burst_start;
    assign dma_axi64_core0_rd_finish = dma_axi64_core0_dma_axi64_core0_ctrl_rd_finish;
    assign dma_axi64_core0_rd_ctrl_busy = dma_axi64_core0_dma_axi64_core0_ctrl_rd_busy;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_rd_hold = dma_axi64_core0_rd_hold_ctrl;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_go = dma_axi64_core0_wr_ch_go_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_full = dma_axi64_core0_wr_cmd_full_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_cmd_pending = dma_axi64_core0_wr_cmd_pending_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num = dma_axi64_core0_wr_ch_num_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_num_resp = dma_axi64_core0_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_go_next_line = dma_axi64_core0_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_valid = dma_axi64_core0_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr = dma_axi64_core0_wr_clr;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_clr_last = dma_axi64_core0_wr_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_periph_delay = dma_axi64_core0_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_clr_stall = dma_axi64_core0_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_tokens = dma_axi64_core0_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_ready = dma_axi64_core0_wr_ready_joint;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_ch_last = dma_axi64_core0_wr_ch_last_joint;
    assign dma_axi64_core0_wr_burst_start = dma_axi64_core0_dma_axi64_core0_ctrl_wr_burst_start;
    assign dma_axi64_core0_wr_finish = dma_axi64_core0_dma_axi64_core0_ctrl_wr_finish;
    assign dma_axi64_core0_wr_ctrl_busy = dma_axi64_core0_dma_axi64_core0_ctrl_wr_busy;
    assign dma_axi64_core0_dma_axi64_core0_ctrl_wr_hold = dma_axi64_core0_wr_hold_ctrl;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_port;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_line_cmd;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_split;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_valid;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_wr_ready;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_last;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_page_cross;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_AWADDR;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_AWPORT;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_AWLEN;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_AWSIZE;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_AWVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_AWREADY;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_WDATA;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_WSTRB;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_WLAST;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_WVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_WREADY;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_BREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_joint_stall;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_w;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_aw;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_w;

    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_AWID  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_AJOINT  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID_d  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_BID  ;
    reg[1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_wr_resp_full  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_BREADY  =1'b1;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_din = dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID_d = dma_axi64_core0_dma_axi64_core0_axim_wr_delay_bvalid_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP_d   <=2'b00;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP_d   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP  ;
            end


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_end_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_extra_bit;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_port;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_pending;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_split;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross;
    reg [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_APORT;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN;
    reg [1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AWVALID;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout;

    reg[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_pre  ;
    wire[32-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR_pre  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE_pre  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_length  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_line_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr  ;
    wire[8:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach_pre  ;
    reg[8:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_cross  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start_d  ;
    wire[8:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst  ;
    reg[8:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst_d  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr  [11:8]==4'hf;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr  [7:0]+  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach  >{1'b1,{8{1'b0}}});
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst  ={1'b1,{8{1'b0}}}-  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr  [7:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_full  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach   <={9{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_reach_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst   <=1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst_d   <={9{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst_d   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start_d  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size  -  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst_d  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_split  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start_d  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_num  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_line_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID  [6];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_pending  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY  )&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_pending   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_pending   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst  ))
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_pending   <=1'b0;



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_high_addr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_high_addr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cross_start_d = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cross_start_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_line_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_line = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_delay_cmd_line_dout;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_pre  ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_end_line_cmd  ,  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE_pre  [1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_extra_bit  ,  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ch_num  [2:0]};
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  =='d1 ? 2'b00:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  =='d2 ? 2'b01:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  =='d4 ? 2'b10:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AXI_WORD_SIZE  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_length  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst   ?   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_size  :  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross   ?   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_max_burst  :  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_length  [8-1:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AXI_3  ]=='d0 ? {4{1'b0}}:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_length  [8-1:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AXI_3  ]-1'b1;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE   <={2{1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT   <=1'b0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE_pre  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_req  ;
            end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg   <={7{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_pre  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID   =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg  ;
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID   [6]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg  [6]&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst  );
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID   [3]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID_reg  [3]&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst  );
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR   <={32{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR  [32-1:12],{12{1'b1}}}+1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_APORT   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_APORT   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_port  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg   <=1'b0;
            else
                if ((  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size  >'d0))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_next_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg   <=1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT   ?   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AWVALID  ):  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID_reg  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_VALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_READY;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_ID;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout;

    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout_num  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_ID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout  =(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter   <={10{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_VALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_READY  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter   <={10{1'b1}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_VALID  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_counter  -1'b1;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_VALID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_READY = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_ID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_dma_axi64_axim_timeout_axim_timeout;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ch_num = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_start = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_addr = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_burst_size = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_end_line_cmd = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_extra_bit = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_port = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_joint_req = dma_axi64_core0_dma_axi64_core0_axim_wr_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_page_cross = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWADDR = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AADDR;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWPORT = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_APORT;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWLEN = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ALEN;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWSIZE = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_ASIZE;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AREADY = dma_axi64_core0_dma_axi64_core0_axim_wr_AWREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AWVALID = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AJOINT = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_AJOINT;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_aw = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_aw = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wcmd_axim_timeout;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rsize;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_valid;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_wr_ready;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_num;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_resp_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_stall;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWID;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWADDR;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWLEN;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWSIZE;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AJOINT;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WDATA;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLAST;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY;

    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_pre  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_pre  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_pre  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_data  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_data  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_data  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_valid_last  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_pre  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size_pre  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_last_channel  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_cmd  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_cmd  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_ready  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness_pre  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_fifo_rd_valid  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_req_out  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_joint  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size_joint  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_full  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_full  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_full  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_full  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end_num  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_ready  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_valid  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness  +  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_ready  -  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness   <=3'd0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_ready  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness_pre  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_SIZE_BITS -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_ch_fifo_rd;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_data_fullness_pre;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_HOLD;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd_valid;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_SIZE_BITS -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size_joint;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_pre  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_rd_stall_num  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_rd_stall  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_DELAY  -1];

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo  +  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint  -  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_ch_fifo_rd  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo   <=3'd0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_ch_fifo_rd  ))
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out  &((  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  >'d2)|((  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  =='d2)&(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_data_fullness_pre  >'d1))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_HOLD  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_data_fullness_pre  >'d1)&(~(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_pre  ));
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_reg   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_count_ch_fifo_pre  =='d0)
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_reg   <=1'b0;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall_reg  |(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_HOLD  );


    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_DELAY  -1];


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_full;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_fullness  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_stall;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_pend  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_pend  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_stall  ))
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count  -1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_din  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_stall  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count  +1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_pend  =(|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_count  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_dout  =(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_din  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_pend  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_stall  );
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_stall = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_stall_joint_fifo_rd_dout;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_req_out = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_req_out;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_ch_fifo_rd = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_data_fullness_pre = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fullness_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_HOLD = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size_joint = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size_joint;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_stall = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_stall;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY  );


    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_DELAY  -1];

    always @(   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_cmd   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_cmd  )
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size   =4'd1;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size   =4'd2;
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size   =4'd4;
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size   =4'd8;
        endcase
    end

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_fifo_rd_valid  |((~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_empty  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall  )&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_wr_ready  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rsize  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_fifo_rd_valid   ?   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size_joint  :  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [5:4]==2'b00 ? 4'd1:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [5:4]==2'b01 ? 4'd2:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [5:4]==2'b10 ? 4'd4:4'd8;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_num  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [2:0];


    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_last_channel   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_last_channel   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_pre  [2:0];

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  [5:4]==2'b00 ? 4'd1:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  [5:4]==2'b01 ? 4'd2:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  [5:4]==2'b10 ? 4'd4:4'd8;


    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num   <=3'd0;
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size   <=3'd0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num_pre  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size_pre  ;
            end

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_valid_last  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_cmd  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_empty  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_valid_last  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_num   <=3'd0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_num   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end_num  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_pre  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_num  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end_num  );


    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_fifo_rd_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_not_ready = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_delay_joint_not_ready_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pending = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_pending_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop_d = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_cmd_pop_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_wr_transfer_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_stall = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_stall_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_delay_clr_line_dout;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_cmd_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_full  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_full  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_resp_full  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_valid_last  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWID  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWLEN  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWSIZE  ;
    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWADDR            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWSIZE   )
    begin
        case ({  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWSIZE  [1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWADDR  [2:0]})
            { 2'b00,3'b000}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_0001;
            { 2'b00,3'b001}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_0010;
            { 2'b00,3'b010}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_0100;
            { 2'b00,3'b011}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_1000;
            { 2'b00,3'b100}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0001_0000;
            { 2'b00,3'b101}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0010_0000;
            { 2'b00,3'b110}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0100_0000;
            { 2'b00,3'b111}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b1000_0000;
            { 2'b01,3'b000}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_0011;
            { 2'b01,3'b010}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_1100;
            { 2'b01,3'b100}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0011_0000;
            { 2'b01,3'b110}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b1100_0000;
            { 2'b10,3'b000}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b0000_1111;
            { 2'b10,3'b100}:
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b1111_0000;
            default :
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre   =8'b1111_1111;
        endcase
    end



    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_fullness  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [6];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_line_end_num  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd  [2:0];
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count   <={4{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_out_count  +1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_push  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLAST  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB  =(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count  [0] ? {  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_data  [3:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_data  [7:4]}:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_data  )&{8{  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  }};
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_fullness  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count   <={4{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count  +1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_valid  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_pre  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_fullness  ;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_joint;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_joint_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_size_joint = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_gen_joint_stall_rd_transfer_fifo_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_push;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_din = {dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AJOINT};
    assign {dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_cmd,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_cmd,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_cmd,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_req_out} = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_empty = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_empty;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_fifo_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_push;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_din = {dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_pre,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_pre};
    assign {dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_data,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSIZE_data,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB_data,dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID_data} = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_empty = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_empty;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_fifo_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_push;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WDATA = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_empty = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_empty;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_fifo_full;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_data_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLAST  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_in_count  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLEN_data  )&(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_cmd_data_empty  );

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_VALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_READY;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_ID;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout;

    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout_num  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_ID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout  =(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter   <={10{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_VALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_READY  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter   <={10{1'b1}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_VALID  )
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_counter  -1'b1;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_VALID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_READY = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_ID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_dma_axi64_axim_timeout_axim_timeout;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer = dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rsize = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rdata = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_ch_fifo_rd_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_next_size = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_resp_full = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_resp_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_cmd_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line_num = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_wr_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_joint_stall = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_joint_stall;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_w = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_w = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_axim_timeout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWID = dma_axi64_core0_dma_axi64_core0_axim_wr_AWID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWADDR = dma_axi64_core0_dma_axi64_core0_axim_wr_AWADDR;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWLEN = dma_axi64_core0_dma_axi64_core0_axim_wr_AWLEN;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWSIZE = dma_axi64_core0_dma_axi64_core0_axim_wr_AWSIZE;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_AWVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AWREADY = dma_axi64_core0_dma_axi64_core0_axim_wr_AWREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_AJOINT = dma_axi64_core0_dma_axi64_core0_axim_wr_AJOINT;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_WDATA = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WDATA;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_WSTRB = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WSTRB;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_WLAST = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WLAST;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_WVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wdata_WREADY = dma_axi64_core0_dma_axi64_core0_axim_wr_WREADY;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_full;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AREADY;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_VALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_READY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_LAST;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_VALID  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_READY  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_LAST  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_pop  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP_SLVERR  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP_DECERR  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last_pre  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ID  [3];

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_clr_last_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_slverr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_delay_decerr_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp_pre  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_full;

    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_fullness  ;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_push;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_din = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_empty = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_empty;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_fifo_full;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clk = dma_axi64_core0_dma_axi64_core0_axim_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_reset = dma_axi64_core0_dma_axi64_core0_axim_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_slverr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_slverr;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_decerr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_decerr;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_last = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num_resp = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_resp_full = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_resp_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AID = dma_axi64_core0_dma_axi64_core0_axim_wr_AWID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_AWVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_AREADY = dma_axi64_core0_dma_axi64_core0_axim_wr_AWREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_RESP = dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_BID = dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_ID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_VALID = dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_READY = dma_axi64_core0_dma_axi64_core0_axim_wr_BREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_dma_axi64_axim_wresp_LAST = 1'b1;

    assign dma_axi64_core0_dma_axi64_core0_axim_wr_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_port = dma_axi64_core0_wr_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_last_cmd = dma_axi64_core0_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_line_cmd = dma_axi64_core0_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num = dma_axi64_core0_wr_ch_num_joint;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_start = dma_axi64_core0_wr_burst_start_joint;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_addr = dma_axi64_core0_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_wr_burst_size = dma_axi64_core0_wr_burst_size;
    assign dma_axi64_core0_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_pending;
    assign dma_axi64_core0_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_split;
    assign dma_axi64_core0_wr_cmd_num = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer = dma_axi64_core0_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_rd_transfer_size = dma_axi64_core0_rd_transfer_size;
    assign dma_axi64_core0_ch_fifo_rd = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rdata = dma_axi64_core0_ch_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_valid = dma_axi64_core0_ch_fifo_rd_valid;
    assign dma_axi64_core0_ch_fifo_rsize = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_wr_ready = dma_axi64_core0_ch_fifo_wr_ready;
    assign dma_axi64_core0_ch_fifo_rd_num = dma_axi64_core0_dma_axi64_core0_axim_wr_ch_fifo_rd_num;
    assign dma_axi64_core0_wr_transfer_num = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_num;
    assign dma_axi64_core0_wr_transfer = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer;
    assign dma_axi64_core0_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_transfer_size;
    assign dma_axi64_core0_wr_next_size = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_next_size;
    assign dma_axi64_core0_wr_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_cmd_full;
    assign dma_axi64_core0_wr_clr_line = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line;
    assign dma_axi64_core0_wr_clr_line_num = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_line_num;
    assign dma_axi64_core0_wr_slverr = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_slverr;
    assign dma_axi64_core0_wr_decerr = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_decerr;
    assign dma_axi64_core0_wr_clr = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr;
    assign dma_axi64_core0_wr_clr_last = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_clr_last;
    assign dma_axi64_core0_wr_ch_num_resp = dma_axi64_core0_dma_axi64_core0_axim_wr_wr_ch_num_resp;
    assign dma_axi64_core0_wr_page_cross = dma_axi64_core0_dma_axi64_core0_axim_wr_page_cross;
    assign dma_axi64_core0_AWADDR = dma_axi64_core0_dma_axi64_core0_axim_wr_AWADDR;
    assign dma_axi64_core0_wr_port_num = dma_axi64_core0_dma_axi64_core0_axim_wr_AWPORT;
    assign dma_axi64_core0_AWLEN = dma_axi64_core0_dma_axi64_core0_axim_wr_AWLEN;
    assign dma_axi64_core0_AWSIZE = dma_axi64_core0_dma_axi64_core0_axim_wr_AWSIZE;
    assign dma_axi64_core0_AWVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_AWVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_AWREADY = dma_axi64_core0_AWREADY;
    assign dma_axi64_core0_WDATA = dma_axi64_core0_dma_axi64_core0_axim_wr_WDATA;
    assign dma_axi64_core0_WSTRB = dma_axi64_core0_dma_axi64_core0_axim_wr_WSTRB;
    assign dma_axi64_core0_WLAST = dma_axi64_core0_dma_axi64_core0_axim_wr_WLAST;
    assign dma_axi64_core0_WVALID = dma_axi64_core0_dma_axi64_core0_axim_wr_WVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_WREADY = dma_axi64_core0_WREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_BRESP = dma_axi64_core0_BRESP;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_BVALID = dma_axi64_core0_BVALID;
    assign dma_axi64_core0_BREADY = dma_axi64_core0_dma_axi64_core0_axim_wr_BREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_wr_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_joint_stall = dma_axi64_core0_dma_axi64_core0_axim_wr_joint_stall;
    assign dma_axi64_core0_timeout_aw = dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_aw;
    assign dma_axi64_core0_timeout_w = dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_w;
    assign dma_axi64_core0_timeout_num_aw = dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_aw;
    assign dma_axi64_core0_timeout_num_w = dma_axi64_core0_dma_axi64_core0_axim_wr_axim_timeout_num_w;


    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_num;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_joint_stall;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_port;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wsize;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_last;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_page_cross;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ARADDR;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_ARPORT;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ARLEN;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_ARSIZE;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_ARVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_ARREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_AWVALID;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY_out;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_ar;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_num_ar;

    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_ARID  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID_d  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_RID  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA_d  ;
    reg[1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP_d  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr  =  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_pre  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_last  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_load  =  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_last  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_din = dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY_out;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_delay_ready_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_din = dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID_d = dma_axi64_core0_dma_axi64_core0_axim_rd_delay_rvalid_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP_d   <=2'b00;
            dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA_d   <={64{1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST_d   <=1'b0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP_d   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP  ;
                dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA_d   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA  ;
                dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST_d   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST  ;
            end

    always @(   dma_axi64_core0_dma_axi64_core0_axim_rd_RID   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_axim_rd_RID  [5:4])
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size   =4'd1;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size   =4'd2;
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size   =4'd4;
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size   =4'd8;
        endcase
    end


    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_end_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_extra_bit;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_port;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_pending;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_full;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_split;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross;
    reg [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_APORT;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN;
    reg [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AWVALID;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AJOINT;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout;

    reg[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg  ;
    wire[7-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_pre  ;
    wire[32-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR_pre  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE_pre  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_length  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr  ;
    wire[8:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach_pre  ;
    reg[8:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_cross  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start_d  ;
    wire[8:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst  ;
    reg[8:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst_d  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr  [11:8]==4'hf;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr  [7:0]+  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr  &(  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach  >{1'b1,{8{1'b0}}});
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst  ={1'b1,{8{1'b0}}}-  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr  [7:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg  )&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_full  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach   <={9{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_reach_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst   <=1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst_d   <={9{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst_d   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start_d  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size  -  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst_d  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_split  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start_d  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_num  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID  [6];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_pending  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY  )&  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AJOINT  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_pending   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_pending   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst  ))
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_pending   <=1'b0;



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_high_addr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_high_addr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cross_start_d = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cross_start_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_delay_cmd_line_dout;

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_pre  ={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_end_line_cmd  ,  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE_pre  [1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_extra_bit  ,  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ch_num  [2:0]};
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  =='d1 ? 2'b00:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  =='d2 ? 2'b01:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  =='d4 ? 2'b10:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AXI_WORD_SIZE  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_length  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst   ?   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_size  :  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross   ?   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_max_burst  :  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_length  [8-1:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AXI_3  ]=='d0 ? {4{1'b0}}:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_length  [8-1:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AXI_3  ]-1'b1;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE   <={2{1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AJOINT   <=1'b0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE_pre  ;
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AJOINT   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_req  ;
            end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg   <={7{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_pre  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg            or    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID   =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg  ;
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID   [6]=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg  [6]&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst  );
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID   [3]=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID_reg  [3]&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst  );
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR   <={32{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR  [32-1:12],{12{1'b1}}}+1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_APORT   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_APORT   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_port  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  |  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg   <=1'b0;
            else
                if ((  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start  &(  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size  >'d0))|  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_next_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg   <=1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AJOINT   ?   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AWVALID  ):  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID_reg  ;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_VALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_READY;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_ID;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout;

    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout_num  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_ID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout  =(  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter   <={10{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_VALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_READY  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter   <={10{1'b1}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_VALID  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_counter  -1'b1;

    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_VALID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_READY = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_ID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_dma_axi64_axim_timeout_axim_timeout;

    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ch_num = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_start = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_addr = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_burst_size = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_end_line_cmd = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_extra_bit = dma_axi64_core0_dma_axi64_core0_axim_rd_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_port = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_joint_req = dma_axi64_core0_dma_axi64_core0_axim_rd_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_pending = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_cmd_line;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_page_cross = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARADDR = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AADDR;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARPORT = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_APORT;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARLEN = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ALEN;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARSIZE = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_ASIZE;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_ARREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_AWVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_AWVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_num_ar = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_ar = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rcmd_axim_timeout;


    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_joint_stall;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wsize;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_burst_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_num;
    reg [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARREADY;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARID;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RDATA;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RLAST;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY_out;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_cmd_id  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre_d  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num_d  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_cmd_id  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [3];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY_out  =(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre  )&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre_d  )&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_joint_stall  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_num  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_cmd_id  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_burst_cmd  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [5];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wdata  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RDATA  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wsize  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RLAST  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [6]&(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [3]);

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre_d = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_delay_clr2_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num_d   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num_d   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_num   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_pre_d  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_num   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num_d  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_cmd_id  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_num  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wdata  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RDATA  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle   <=2'b00;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle  [0]&1'b1)
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle   <=2'b00;
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr  )
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle  +1'b1;

    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_joint_stall = dma_axi64_core0_dma_axi64_core0_axim_rd_joint_stall;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wdata = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wsize = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ch_fifo_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_cmd = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_burst_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_load_wdata = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line_num = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_rd_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_ARVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_ARREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_ARID = dma_axi64_core0_dma_axi64_core0_axim_rd_ARID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RID = dma_axi64_core0_dma_axi64_core0_axim_rd_RID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RDATA = dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RLAST = dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY_out = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rdata_RREADY_out;


    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last;
    reg [2:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_full;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AVALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AREADY;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP;
    wire [7-1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_VALID;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_READY;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_LAST;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_push  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AVALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AREADY  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_pop  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_VALID  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_READY  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_LAST  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_pop  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ID  [2:0];
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP  ==  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP_SLVERR  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP  ==  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP_DECERR  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last_pre  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ID  [3];

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_din;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_dout  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_clr_last_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_slverr_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr_pre;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_delay_decerr_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_pre  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp_pre  ;


    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_push;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_pop;
    wire [ dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_din;
    reg [ dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_empty;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_full;

    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_pop  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_out  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  -1:0];
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_next  ;
    reg  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in  ;
    reg[  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_BITS  -1:0]  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_push  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_push  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_empty  &(  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty  |  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_pop  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_pop  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_pop  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  =!  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_push  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_push  );
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  =!  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_SINGLE  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_pop  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_pop  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_push  )
            begin
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_din  ;
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty   <=1'b0;
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reg_pop  )
                begin
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_WIDTH  {1'b0}};
                    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty   <=1'b1;
                end
                else
                    if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo  [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out  ];
                        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty   <=1'b0;
                    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in  ==  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH_BITS  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out   <=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out  ==  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_LAST_LINE   ? 0:  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out  +1'b1;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo   [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in  ]<=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_din  ;

    always @(    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push            or    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_in   ={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_in   [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_in  ]=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  ;
    end

    always @(    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop            or    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out   )
    begin
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_out   ={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  {1'b0}};
        dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_out   [  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_ptr_out  ]=  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  ;
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset  )
            dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness   <={  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_DEPTH  {1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_push  |  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_pop  )
                dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness   <=(  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness  &(~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_out  ))|  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness_in  ;

    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_next  =|  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_empty  =~  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_next  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_empty  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fifo_empty  &  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_full  =  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_SINGLE   ? !  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout_empty  :&  dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_fullness  ;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_push = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_push;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_pop = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_pop;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_din = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_dout;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_empty = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_empty;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_full = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_fifo_full;

    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clk = dma_axi64_core0_dma_axi64_core0_axim_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_reset = dma_axi64_core0_dma_axi64_core0_axim_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_slverr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_slverr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_decerr = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_decerr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_pre = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_last = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num_resp = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_resp_full;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AID = dma_axi64_core0_dma_axi64_core0_axim_rd_ARID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_ARVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_AREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_ARREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_RESP = dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RID = dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_ID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_VALID = dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID_d;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_READY = dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_dma_axi64_axim_rresp_LAST = dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST_d;

    assign dma_axi64_core0_dma_axi64_core0_axim_rd_clk = dma_axi64_core0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_load_wr = dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr;
    assign dma_axi64_core0_load_wr_num = dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_num;
    assign dma_axi64_core0_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_axim_rd_load_wr_cycle;
    assign dma_axi64_core0_load_wdata = dma_axi64_core0_dma_axi64_core0_axim_rd_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_joint_stall = dma_axi64_core0_joint_stall;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_joint_req = dma_axi64_core0_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_line_cmd = dma_axi64_core0_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_load_req_in_prog = dma_axi64_core0_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_port = dma_axi64_core0_rd_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num = dma_axi64_core0_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_start = dma_axi64_core0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_addr = dma_axi64_core0_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_size = dma_axi64_core0_rd_burst_size;
    assign dma_axi64_core0_rd_cmd_pending = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_pending;
    assign dma_axi64_core0_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_split;
    assign dma_axi64_core0_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_line;
    assign dma_axi64_core0_rd_cmd_num = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_num;
    assign dma_axi64_core0_rd_cmd_full = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_cmd_full;
    assign dma_axi64_core0_ch_fifo_wr = dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr;
    assign dma_axi64_core0_ch_fifo_wdata = dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wdata;
    assign dma_axi64_core0_ch_fifo_wsize = dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wsize;
    assign dma_axi64_core0_ch_fifo_wr_num = dma_axi64_core0_dma_axi64_core0_axim_rd_ch_fifo_wr_num;
    assign dma_axi64_core0_rd_transfer_num = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_num;
    assign dma_axi64_core0_rd_transfer = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer;
    assign dma_axi64_core0_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_transfer_size;
    assign dma_axi64_core0_rd_burst_cmd = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_burst_cmd;
    assign dma_axi64_core0_rd_clr_line = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line;
    assign dma_axi64_core0_rd_clr_line_num = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_line_num;
    assign dma_axi64_core0_rd_slverr = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_slverr;
    assign dma_axi64_core0_rd_decerr = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_decerr;
    assign dma_axi64_core0_rd_clr = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr;
    assign dma_axi64_core0_rd_clr_load = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_load;
    assign dma_axi64_core0_rd_clr_last = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_clr_last;
    assign dma_axi64_core0_rd_ch_num_resp = dma_axi64_core0_dma_axi64_core0_axim_rd_rd_ch_num_resp;
    assign dma_axi64_core0_rd_page_cross = dma_axi64_core0_dma_axi64_core0_axim_rd_page_cross;
    assign dma_axi64_core0_ARADDR = dma_axi64_core0_dma_axi64_core0_axim_rd_ARADDR;
    assign dma_axi64_core0_rd_port_num = dma_axi64_core0_dma_axi64_core0_axim_rd_ARPORT;
    assign dma_axi64_core0_ARLEN = dma_axi64_core0_dma_axi64_core0_axim_rd_ARLEN;
    assign dma_axi64_core0_ARSIZE = dma_axi64_core0_dma_axi64_core0_axim_rd_ARSIZE;
    assign dma_axi64_core0_ARVALID = dma_axi64_core0_dma_axi64_core0_axim_rd_ARVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_ARREADY = dma_axi64_core0_ARREADY;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_AWVALID = dma_axi64_core0_AWVALID;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RDATA = dma_axi64_core0_RDATA;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RRESP = dma_axi64_core0_RRESP;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RLAST = dma_axi64_core0_RLAST;
    assign dma_axi64_core0_dma_axi64_core0_axim_rd_RVALID = dma_axi64_core0_RVALID;
    assign dma_axi64_core0_RREADY = dma_axi64_core0_dma_axi64_core0_axim_rd_RREADY_out;
    assign dma_axi64_core0_timeout_ar = dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_ar;
    assign dma_axi64_core0_timeout_num_ar = dma_axi64_core0_dma_axi64_core0_axim_rd_axim_timeout_num_ar;

    assign   dma_axi64_core0_rd_hold  =1'b0;
    assign   dma_axi64_core0_wr_hold  =1'b0;

    wire  dma_axi64_core0_dma_axi64_core0_channels_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_penable;
    wire [10:0] dma_axi64_core0_dma_axi64_core0_channels_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_pending;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_load_wr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_load_wr_num;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_load_req_in_prog;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_decerr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num_resp;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_clr_last;
    wire [8*1-1:0] dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_start;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_idle;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_active;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_timeout_ar;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_timeout_num_aw;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_timeout_num_w;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_timeout_num_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wdt_timeout;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wdt_ch_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_fifo_wr_ready;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_port;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_rd_periph_delay;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_port;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_joint_mux_in_prog;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req;

    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_psel  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr  ;
    wire[32*8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_prdata  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_joint_end  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start  ;
    wire[8*32-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr  ;
    wire[8*8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size  ;
    wire[8*6-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num  ;
    wire[8*3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start  ;
    wire[8*32-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr  ;
    wire[8*8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size  ;
    wire[8*6-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num  ;
    wire[8*3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid  ;
    wire[8*31-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr  ;
    wire[8*31-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid  ;
    wire[8*64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_penable;
    wire [10:8] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pslverr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_psel;
    wire [32*8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_prdata;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_pslverr;

    wire[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d   <=3'b000;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_psel  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_penable  ))
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel  ;
            else
                if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_psel  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pclken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d   <=3'b000;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr  [10:8];

    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x;

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x  ;
        endcase
    end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_psel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_psel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_psel_ch_x;


    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x;

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_WIDTH  -1:0];
        endcase
    end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_prdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_mux_prdata_x;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pslverr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_pslverr  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr_sel_d  ];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_clk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_psel = dma_axi64_core0_dma_axi64_core0_channels_psel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[10:8];
    assign dma_axi64_core0_dma_axi64_core0_channels_prdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_pslverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_psel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_psel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_prdata = dma_axi64_core0_dma_axi64_core0_channels_ch_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_apb_mux_ch_pslverr = dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr;


    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd_valid;
    wire [8*64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rdata;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rdata;
    wire [8*31-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_rx_clr;
    wire [30:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_rx_clr;
    wire [8*31-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_tx_clr;
    wire [30:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_tx_clr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_page_cross;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_ar;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_aw;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_w;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_timeout;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_ch_num;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_aw;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_w;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_ar;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_mux_in_prog;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_in_prog;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_not_in_prog;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_pending;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_pending;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_port;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_stall;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_req_in_prog;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_line_cmd;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_go_next_line;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_start;
    wire [8*32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_addr;
    wire [8*8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_size;
    wire [8*6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_tokens;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_port_num;
    wire [8*3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_periph_delay;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_valid;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_split;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_line;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_stall;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_wr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_transfer;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_line;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_load;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_slverr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_decerr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_load;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_port;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_stall;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_last_cmd;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_line_cmd;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_go_next_line;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_start;
    wire [8*32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_addr;
    wire [8*8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_size;
    wire [8*6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_tokens;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_port_num;
    wire [8*3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_periph_delay;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_valid;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_split;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_stall;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer_num;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_line_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_ready;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_transfer;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_line;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr_ready;
    wire [2:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_last;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_slverr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_decerr;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_last;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr;


    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_x;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_x;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_WIDTH  *7];



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_WIDTH  *7];



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_WIDTH  *7];



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_WIDTH  *7];


    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_sel;
    wire [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x;

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_WIDTH  -1:0];
        endcase
    end



    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_sel;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x;
    reg [8* dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x;

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x  ;
        endcase
    end




    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_WIDTH  *7];



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_WIDTH  *7];



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_x  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *0]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *1]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *2]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *3]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *4]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *5]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *6]|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_WIDTH  *7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_2_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_3_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_rx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_4_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_tx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_5_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_55_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_not_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_56_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_mux_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_57_x;



    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x  ;
        endcase
    end


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_go_next_line  ='d0;


    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_WIDTH  -1:0];
        endcase
    end


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_port  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_port  ='d0;


    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x  ;
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_sel            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   ={8*  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  {1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  *7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_WIDTH  -1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x  ;
        endcase
    end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_6_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_7_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_8_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_9_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_60_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_11_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_13_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_15_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_16_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_17_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_39_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_20_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_42_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_58_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_59_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_18_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_load;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_19_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_21_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_34_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_37_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_38_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_40_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_41_ch_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_43_ch_x;



    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_WIDTH  -1:0];
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_sel   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_sel  )
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *1];
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *2];
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *3:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *3];
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *4];
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *5:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *5];
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *6:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *6];
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1+  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *7:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  *7];
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_WIDTH  -1:0];
        endcase
    end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_30_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_51_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_33_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_53_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_23_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_26_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_27_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_28_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_49_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_31_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_last_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_44_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_47_x;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_sel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_ch_x = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_mux_48_x;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_rx_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_periph_rx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_periph_tx_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_periph_tx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_wr_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_timeout_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_timeout_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_timeout_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_aw = dma_axi64_core0_dma_axi64_core0_channels_timeout_num_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_w = dma_axi64_core0_dma_axi64_core0_channels_timeout_num_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_timeout_num_ar = dma_axi64_core0_dma_axi64_core0_channels_timeout_num_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_wdt_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wdt_ch_num = dma_axi64_core0_dma_axi64_core0_channels_wdt_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_timeout_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wdt_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_joint_not_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_joint_mux_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_not_in_prog = dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_joint_mux_in_prog = dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num = dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_num = dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_port = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_tokens = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_port_num = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_cmd_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr_num = dma_axi64_core0_dma_axi64_core0_channels_load_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_load_wr = dma_axi64_core0_dma_axi64_core0_channels_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_num = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer_num = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_line_num = dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_ch_num_resp = dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_rd_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_rd_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_rd_clr_load;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_rd_clr_load;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num = dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_num = dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_last_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_port = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_port;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_last_cmd = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_tokens = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_port_num = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd_num = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer_num = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_line_num = dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_ch_num_resp = dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_wr_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_wr_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_wr_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_wr_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_channels_mux_ch_wr_clr;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req;

    wire[32-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_addr  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_in_prog  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  ;
    wire[32-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_start_addr  ;
    wire[32-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_start_addr  ;
    wire[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size  ;
    wire[10-8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_y_size  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_block  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_frame_width  ;
    wire[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_width_align  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_block  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_block  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_max  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_max  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_limit  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_limit  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_incr  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_max_size  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_max_size  ;
    wire[4:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_num  ;
    wire[4:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_num  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outstanding  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outstanding  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_retry_wait  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_in_prog  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_end_swap  ;
    wire[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_offset  ;
    wire[10-8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_y_offset  ;
    wire[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_remain  ;
    wire[10-8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_remain  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ch_end  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_empty  ;
    wire[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_align  ;
    wire[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_offset  ;
    wire[10-8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_y_offset  ;
    wire[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_remain  ;
    wire[10-8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_remain  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_line_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_empty  ;
    wire[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_align  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end_pre  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end_reg  ;
    wire[5:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_gap  ;
    wire[5:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_fullness  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_outs  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_stall  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_rresp  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_outs  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_empty  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_wresp  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_last  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_flush  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_burst_req  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_last  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_single  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_flush  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_line_req  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_overflow  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_underflow  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_block_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_block  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_block_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_block  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_mux  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_line_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_allow_line_cmd  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_cmd  ;
    wire[4:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_bus  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_flush  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_page_cross  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port0_mux  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port1_mux  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk_en  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_active  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_in_prog  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_empty  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start  );

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog   <=(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  );
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_empty  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog   <=(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  );
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_empty  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_empty  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_empty  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_page_cross  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg   <=1'b1;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_not_in_prog  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg   <=1'b0;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_page_cross  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_page_cross  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_page_cross  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_in_prog  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_in_prog  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_not_in_prog  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_not_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_not_in_prog  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port0_mux  =((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_port_num  ==1'b0)|((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_port_num  ==1'b0)))&0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port1_mux  =((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_port_num  ==1'b1)|((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_port_num  ==1'b1)))&0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mux_in_prog  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_in_prog  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port0_mux  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_access_port1_mux  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_ready  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_flush  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_flush  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_block  =1'b1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_block  =1'b1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_mux  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_stall  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_stall  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_allow_line_cmd  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_cmd  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_line_cmd  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_block  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_retry_wait  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_block  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_retry_wait  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ready  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_stall  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_stall  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_rd_active  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_ready  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_ready  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ready  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_stall  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_wr_active  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_ready  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_last_cmd  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_empty  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_cmd  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_outs  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_split  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_outs  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_split  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_load  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_bus  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_aw  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_w  ,{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_wresp  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_aw  )},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_ar  ,{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_rresp  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_ar  )}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk_en  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_active  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update  |(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty  )|(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_ready  )|(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_ready  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle_pre  =!  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk_en  ;


    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_outs_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_outs_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_rd_clr_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_wr_clr_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_delay_idle_dout;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata;
    reg [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr;
    wire [4:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_bus;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_decerr;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_wr_active;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_in_prog;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_x_offset;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_y_offset;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_x_offset;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_y_offset;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_fullness;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_gap;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_overflow;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_underflow;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_x_size;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_y_size;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_line_cmd;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_width_align;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_block;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_block;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_outs_empty;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wait_limit;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_wait_limit;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr;
    wire [4:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num;
    wire [4:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_flush;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap;

    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog_reg  ;
    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size  ;
    reg[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mux  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_auto_retry_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_auto_retry  ;
    reg[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap_reg  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_rd  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_pre  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_block_reg  ;
    reg[6-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens_reg  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_port_num_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num_cfg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_port_num  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding_cfg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr_reg  ;
    reg[4:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num_reg  ;
    reg[12-1:4]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wait_limit_reg  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_rd  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_pre  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_reg  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_block_reg  ;
    reg[6-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens_reg  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding_cfg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr_reg  ;
    reg[4:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num_reg  ;
    reg[12-1:4]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_wait_limit_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_allow_full_fifo  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_allow_full_fifo  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_burst  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_joint_burst  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int_reg  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last_reg  ;
    reg[32-1:2]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr_reg  ;
    reg[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last  ;
    wire[32-1:2]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_set  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_clear  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_int  ;
    wire[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_proc_num  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_proc_num_reg  ;
    wire[13-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_bus  ;
    wire[13-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_rawstat  ;
    reg[13-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable  ;
    wire[13-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_status  ;
    wire[7:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_all_proc_bus  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line0  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line1  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line3  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line0  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line1  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line3  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line4  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_enable  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_start  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_rawstat  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_clear  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_enable  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_frame_width  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line0  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line1  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line2  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line3  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_enable  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_rawstat  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_enable  ;
    reg[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_status  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle0  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle1  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle3  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr0  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr1  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr3  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_last  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_aw  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_w  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_b  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_ar  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_r  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait_pre  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_int  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_paddr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_penable  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwrite  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_penable  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwrite  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line0  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE0  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line1  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE1  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line2  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE2  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line3  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE3  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line0  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE0  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line1  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE1  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line2  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE2  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line3  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE3  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line4  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE4  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_enable  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ENABLE  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_start  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_START  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_start  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_rawstat  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_RAWSTAT  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_clear  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_CLEAR  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_enable  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_ENABLE  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle0  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle  ==2'd0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle1  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle  ==2'd1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle2  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle  ==2'd2;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle3  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle  ==2'd3;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr0  =0 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle0  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle0  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr1  =0 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle1  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle0  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr2  =0 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle2  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle1  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr3  =0 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle3  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle1  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_last  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr3  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr   <={32{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line0  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [32-1:0];
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr0  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [32-1:0];
                end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr   <={32{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line1  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [32-1:0];
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr1  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [32+32-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  -1:32-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  ];
                end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size   <={10{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line2  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [10-1:0];
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr2  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [10-1:0];
                end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int_reg   <=1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last_reg   <=1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr_reg   <={30{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_cmd_line3  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [0];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [1];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [32-1:2];
            end
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr3  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [32-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  ];
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [33-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  ];
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata  [32+32-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  -1:34-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_DATA_SHIFT  ];
                end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg   <={12{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_start  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg   <={12{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg  +1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_start  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg   <={4{1'b0}};
            else
                if ((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_int  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_clear  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg  +(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_int  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )-  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_clear  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_x_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block   ? {{10-8{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size  [8-1:0]}:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_y_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size  [10-1:8]:'d1;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg   <='d0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens_reg   <='d1;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max_reg   <={4{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr_reg   <='d1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line0  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [8-1:0];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [6+16-1:16];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [4+24-1:24];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [31];
            end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_reg   <='d0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens_reg   <='d1;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max_reg   <={4{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr_reg   <='d1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line1  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [8-1:0];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [6+16-1:16];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [4+24-1:24];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [31];
            end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding_cfg  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding_cfg  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mux   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens_reg  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mux   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max_reg  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_allow_full_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr  [5-1:0]=='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_allow_full_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr  [5-1:0]=='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_allow_full_fifo  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_allow_full_fifo  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mux   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_pre  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_joint_burst  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_flush  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_page_cross  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_cross  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_burst  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_joint_burst  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_d  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_DELAY  -1];


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_update;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_start_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_reg;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_other;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_burst;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_fifo;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_joint_flush;
    reg [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_update;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_start_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_reg;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_other;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_burst;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_fifo;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_joint_flush;
    reg [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size;

    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_fifo  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_burst  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_LARGE_FIFO   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_joint_flush  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_SMALL_FIFO   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES  :(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_other  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES  )&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_reg  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES  )&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_other  !=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_reg  ) ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_fifo   ? 32:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_HALF_BYTES  ;

    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_min;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_min;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_b  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_pre  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_MAX_BURST  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_pre  ;




    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_fifo  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_burst  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_LARGE_FIFO   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_MAX_BURST  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_joint_flush  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_SMALL_FIFO   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES  :(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_other  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES  )&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_reg  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES  )&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_other  !=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_reg  ) ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_fifo   ? 32:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_HALF_BYTES  ;


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_b  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_reg;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_min2_max_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_reg;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_min2_max_min;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_pre  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_MAX_BURST   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_MAX_BURST  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_pre  ;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_reg = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size_other = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_burst = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_burst;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_allow_full_fifo = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_rd_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_reg = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_reg;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size_other = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_burst = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_allow_full_fifo = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_dma_axi64_core0_ch_reg_size_wr_burst_max_size;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg   <=1'b1;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap_reg   <=2'b00;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line2  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [16];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [29:28];
            end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem   <=(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num  =='d0)&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num  =='d0)&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_line_cmd  );

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mode  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem  &1'b1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mux  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_port_num  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num_cfg  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width  ={12{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_width_align  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width  [3-1:0];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wait_limit  ={12-4{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_wait_limit  ={12-4{1'b0}};
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num_reg   <='d0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay_reg   <='d0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num_reg   <='d0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay_reg   <='d0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_static_line4  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [4:0];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [3+8-1:8];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [20:16];
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [3+24-1:24];
            end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_block  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_block  =1'b0;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable   <=1'b1;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_enable  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [0];
            end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_in_prog   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_underflow  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_overflow  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog   <=1'b0;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_underflow  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_overflow  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog   <=1'b0;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog_reg   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog_reg   <=1'b0;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog_reg   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_cmd  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog_reg   <=1'b0;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_auto_retry  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_start  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_last  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_pre  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update   <=1'b1;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update   <=1'b0;



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_burst_max_size_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_max_size_update_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_delay_ch_update_dout;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last  ))|(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_x_size  =='d0));
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_addr  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr  [32-1:2],2'b00};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_clr_last  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_int  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_rd_active  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_wr_active  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_in_prog  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_set  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_clear  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_clear  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [0];
    assign {  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_aw  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_w  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_b  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_ar  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_r  }=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_bus  [4:0];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_bus  ={13{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken  }}&{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wdt_timeout  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_aw  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_w  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_b  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_ar  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_r  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_underflow  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_overflow  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_decerr  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_decerr  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_slverr  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_slverr  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_end_set  };

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_pwdata;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_int_bus;
    reg [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_rawstat;

    wire[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write_bus  ;
    wire[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear_bus  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write_bus  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE  {  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_pwdata  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear_bus  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE  {  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_pwdata  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_rawstat   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_SIZE  {1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_rawstat   <=(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_rawstat  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_int_bus  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write_bus  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear_bus  );

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_clear = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_clear;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_write = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_rawstat;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_pwdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata[13-1:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_int_bus = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_bus;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_rawstat = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rawstat_rawstat;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable   <={13{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_int_enable  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata  [13-1:0];

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_status  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_rawstat  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_int  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_status  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_proc_num  =3'd0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_all_proc  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_int  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_rd  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_rd  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_reg  ;
    always @(                                                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_burst                                                                                                                            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo                                                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_joint_burst                                                                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_line_cmd                                                                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_auto_retry                                                               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block                                                              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size                                                             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable                                                            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_rd_active                                                           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_wr_active                                                          or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter                                                         or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last                                                        or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr                                                       or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_port_num                                                      or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int                                                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap                                                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width                                                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter                                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable                                                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_proc_num                                                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_rawstat                                               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_status                                              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg                                             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_allow_full_fifo                                            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_rd                                           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_gap                                          or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr                                         or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs                                        or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max                                       or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding                                      or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding_cfg                                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_block_reg                                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay                                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num_cfg                                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr                                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens                               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wait_limit                              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_x_offset                             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_y_offset                            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem                           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_allow_full_fifo                          or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_rd                         or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_fullness                        or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr                       or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs                      or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding_cfg                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_block_reg                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_wait_limit            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_x_offset           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_y_offset   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line0   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line1   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line2   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line3   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_enable   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_rawstat   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_enable   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_status   ={32{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line0   [32-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line1   [32-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line2   [10-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_buff_size  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3   [0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_set_int  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3   [1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_last  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3   [32-1:2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_next_addr  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   [8-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size_rd  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   [6+16-1:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   [4+24-1:24]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   [30]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding_cfg  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0   [31]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   [8-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size_rd  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   [6+16-1:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   [4+24-1:24]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   [30]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding_cfg  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1   [31]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [12-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [15]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_reg  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [17]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_auto_retry  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [20]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_port_num  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [21]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num_cfg  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [22]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [26:24]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_proc_num  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2   [29:28]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4   [4:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4   [3+8-1:8]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4   [20:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4   [3+24-1:24]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_allow_full_fifo  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_allow_full_fifo  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [2]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_fifo  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [3]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_full_burst  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [4]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_joint_burst  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [5]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [6]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [7]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_line_cmd  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict   [8]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_simple_mem  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets   [10-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_x_offset  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets   [10-8+16-1:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_y_offset  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets   [10-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_x_offset  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets   [10-8+16-1:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_y_offset  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness   [5:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_gap  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness   [5+16:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_fullness  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs   [4-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs   [4-1+8:8]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_enable   [0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_enable  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active   [0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_rd_active  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active   [1]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_wr_active  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter   [12-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_cmd_counter  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter   [4-1+16:16]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_counter  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_rawstat   [13-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_rawstat  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_enable   [13-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_enable  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_status   [13-1:0]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_status  ;
    end

    always @(                       dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr                                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active                             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_enable                            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter                           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line0                          or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line1                         or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line2                        or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3                       or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs                      or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_enable                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_rawstat                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_status                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line3            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   ={32{1'b0}};
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE0   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line0  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE1   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line1  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE2   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line2  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE3   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_line3  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE0   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line0  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE1   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line1  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE2   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line2  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE3   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line3  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE4   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_static_line4  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RESTRICT   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_restrict  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RD_OFFSETS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_rd_offsets  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_WR_OFFSETS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wr_offsets  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_FIFO_FULLNESS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_fifo_fullness  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_OUTS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_outs  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ENABLE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_enable  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_START   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   ={32{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ACTIVE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_active  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_CMD_COUNTER   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_cmd_counter  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_RAWSTAT   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_rawstat  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_CLEAR   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   ={32{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_ENABLE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_enable  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_STATUS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_int_status  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre   ={32{1'b0}};
        endcase
    end

    always @(      dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpaddr  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE0   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE1   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE2   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_LINE3   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE0   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE1   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE2   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE3   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_STATIC_LINE4   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RESTRICT   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_RD_OFFSETS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_WR_OFFSETS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_FIFO_FULLNESS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CMD_OUTS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ENABLE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_START   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_ACTIVE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_CH_CMD_COUNTER   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_RAWSTAT   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_CLEAR   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_ENABLE   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_INT_STATUS   :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  ;
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel  ;
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata   <={32{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata_pre  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata   <={32{1'b0}};

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr   <=1'b0;
        else
            if ((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpread  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_gpwrite  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr_pre  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr   <=1'b0;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_clken = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pclken = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_psel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_psel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_penable = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_paddr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_paddr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwrite = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pwdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_prdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pslverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_timeout_bus = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_bus;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wdt_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_load_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_int_all_proc = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_rd_active = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_wr_active = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_x_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_y_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_y_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_x_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_y_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_y_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_fullness = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_fullness;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_gap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_gap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_overflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_overflow;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_fifo_underflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_underflow;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_x_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_y_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_y_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_block = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_block;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_allow_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_allow_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_frame_width = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_frame_width;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_width_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_width_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_block = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_block;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_block = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_block;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_tokens = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_port_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_port_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_max = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs_max;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_max = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs_max;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outs = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outs = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_limit = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_wait_limit;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_limit = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_wait_limit;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_periph_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_periph_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_wr_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_rd_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_retry_wait = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_ch_retry_wait;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_reg_end_swap;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_last;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_load_req_in_prog;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_size;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_y_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_offset;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_y_offset;
    reg [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clr_remain;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_line_empty;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_empty;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_start_align;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_width_align;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_align;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_last;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_load_req_in_prog;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_size;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_y_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_offset;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_y_offset;
    reg [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain;
    wire [10-8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clr_remain;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_line_empty;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_empty;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_start_align;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_width_align;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_align;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_update_line  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_line_end_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_update_d  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_start  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_last  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_go_next_line  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_line_empty  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_empty  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end_pre  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end_pre  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end   <=1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain   <={10{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_go_next_line  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_size  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_start  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_load_req_in_prog  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_size  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_offset  ={10{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_y_offset  ={10-8{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clr_remain  ={10-8{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_align  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_start_align  ;



    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_update_line  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_line_end_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_update_d  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_start  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_last  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_go_next_line  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_line_empty  =1'b0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_empty  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end_pre  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end_pre  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end   <=1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain   <={10{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_go_next_line  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_size  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_start  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_load_req_in_prog  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_size  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_offset  ={10{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_y_offset  ={10-8{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clr_remain  ={10-8{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_align  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_start_align  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_y_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_y_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_y_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_y_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clr_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_line_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_start_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_start_addr[3-1:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_width_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_width_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_rd_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_load_req_in_prog = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_y_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_y_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_y_offset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_y_offset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clr_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_line_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_line_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_start_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_start_addr[3-1:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_width_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_width_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_offsets_wr_align;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_start;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_start;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_line_cmd_valid  ;
    reg[5+1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg  ;
    reg[5+1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_qual  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_qual  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size_valid  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size_valid  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size_valid  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size_valid  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_line_cmd_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_line_cmd  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_start  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_qual  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_start  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_load_req_in_prog  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_qual  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_start  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size_valid   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_qual  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size_valid   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size  ;
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size_valid   <={8{1'b0}};

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size_valid   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_qual  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size_valid   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size  ;
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size_valid   <={8{1'b0}};

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size_valid  ={4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size_valid  ={4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg   <={1'b0,1'b1,{5{1'b0}}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg   <={1'b0,1'b1,{5{1'b0}}};
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size_valid  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size_valid  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg  [5+1] ? 'd0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap_reg  [5:0];
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg   <={5+1{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg   <={5+1{1'b0}};
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size_valid  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size_valid  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg  [5+1] ? 'd0:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness_reg  [5:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_gap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_rd_gap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_fullness = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_remain_wr_fullness;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clr;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_max;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_empty;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clr;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_max;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_empty;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_timeout;

    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_pre  ;
    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_empty  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs  =='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_cmd  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clr  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs   <='d0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_cmd  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_stall   <=1'b0;
        else
            if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_max  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_stall   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs  >=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_max  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_timeout  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter   <={10{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter   <={10{1'b1}};
            else
                if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_counter  -1'b1;




    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_pre  ;
    reg[10-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_empty  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs  =='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_cmd  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clr  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs   <='d0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_cmd  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_stall   <=1'b0;
        else
            if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_max  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_stall   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs  >=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_max  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_timeout  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter  =='d0);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter   <={10{1'b1}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter   <={10{1'b1}};
            else
                if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_counter  -1'b1;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_max = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_max;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_stall = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_rresp = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_rd_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_cmd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_max = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_max;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_wresp = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_outs_wr_timeout;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_stall_pre  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req  );

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_req_in_prog;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_outs_empty;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_max_size;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_start_addr;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_frame_width;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_last;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_ready;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_single;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_req_in_prog;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_outs_empty;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_max_size;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_start_addr;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_frame_width;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_last;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_ready;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_single;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_burst_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_burst_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush_in;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d3  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_DELAY  -1];

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_single   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_start  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_single   <=(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_size  <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_SINGLE_SIZE  );


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_ch_update_d;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_in_prog;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_incr;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_start_addr;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_x_size;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_size;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_ch_update_d;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_in_prog;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_addr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_incr;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_start_addr;
    wire [12-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_x_size;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_size;
    reg [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_go_next_line_d  ;
    reg[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width_diff_reg  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width_diff  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width_diff  ={12{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_go_next_line_d  =1'b0;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr   <={32{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_in_prog  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_addr  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_ch_update_d  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_start_addr  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_start  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_incr  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_size  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_go_next_line_d  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_incr  )
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width_diff  ;



    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d2;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d3;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_outs_empty;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_max_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_last;
    reg [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d2;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d3;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_req_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_outs_empty;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_max_size;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_last;
    reg [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_out;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush_in;

    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain_fifo  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_max_burst_align  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_update  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_wait  ;
    reg[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_size  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_size  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_buffer_small  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_release_fifo  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain_fifo  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain  [10-1:8] ? {1'b1,{8-1{1'b0}}}:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain  [8-1:0];

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_reset;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_c;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_reset;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_c;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min;

    wire[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab_pre  ;
    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab  ;
    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_c  ;

    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_min;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_min;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_min;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_min;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_b  ;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_b  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_c   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_WIDTH  {1'b0}};
        end
        else
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab_pre  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_c   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_c  ;
        end


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_max_burst_align  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [0] ? 'd1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [2] ? 'd4:{1'b1,{8-1{1'b0}}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  [8-1:3] ? {  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  [8-1:3],3'b000}:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  [2] ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre  [0] ? 'd1:'d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready_pre  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_remain  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_release_fifo  );

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  -1];

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_last  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d2  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d3  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_req_in_prog  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                else
                    if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_buffer_small  ))
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready_pre  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_wait  |(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_page_cross  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size  !=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  )))
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready   <=|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_req_in_prog  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_CMD_SIZE  ;
            else
                if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_size  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_buffer_small  ))
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_size  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_update  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d2  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush_in  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_in  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg  [0] ? 2'b11:2'b01;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush_in  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_in  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [2:0]==3'd0 ? 4'd8:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [1:0]==2'd0 ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [0]==1'd0 ? 'd2:'d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [0] ? 'd1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr  [2]&(!0) ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req  [1] ? 'd32:'d16;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty;
    wire [10-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready;
    wire [5:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small;

    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  )&(|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain  )|(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain  <'d8);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=1'b0;
        else
            if ((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end  ))
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=1'b0;
            else
                if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  ;

    always @(               dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE  )
                                begin
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b1;
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                                end
                                else
                                begin
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                                end
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
                    end
                    else
                    begin
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                    end
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS  ;
                else
                    if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK  ;
                        end
                        else
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b1;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ  )
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
                end
                else
                    if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )|(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                    begin
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain  <='d16))
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain  =='d0)
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ  ;
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        end
                        else
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
                    end
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush   =1'b1;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
            end
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns  ;


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_release_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_out  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_cross  );




    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d3  ;


    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc0_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc1_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d3 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_delay_calc2_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc0_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc1_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d3 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_delay_calc2_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_single   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_start  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_single   <=(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_size  <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_SINGLE_SIZE  );



    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_go_next_line_d  ;
    reg[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width_diff_reg  ;
    wire[12-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width_diff  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width_diff  ={12{1'b0}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_go_next_line_d  =1'b0;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr   <={32{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_in_prog  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_addr  ;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_ch_update_d  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_start_addr  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_start  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_incr  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_size  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_go_next_line_d  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_incr  )
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width_diff  ;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_load_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_frame_width = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_frame_width;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_addr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_load_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_frame_width = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_frame_width;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_addr_burst_addr;



    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain_fifo  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_max_burst_align  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_update  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_wait  ;
    reg[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg  ;
    wire[1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_size  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_size  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_buffer_small  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_release_fifo  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain_fifo  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain  [10-1:8] ? {1'b1,{8-1{1'b0}}}:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain  [8-1:0];


    wire[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab_pre  ;
    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab  ;
    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH  -1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_c  ;


    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_b  ;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_b  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_a;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_b;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_ab_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_ab;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min_c;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min2_abc_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_a;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_b;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_ab_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_c;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min2_abc_min;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH  {1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_c   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_WIDTH  {1'b0}};
        end
        else
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_ab_pre  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min_c   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_c  ;
        end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_max_burst_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_c = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_min3_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_max_burst_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_c = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_min3_min;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_max_burst_align  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [0] ? 'd1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [2] ? 'd4:{1'b1,{8-1{1'b0}}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  =|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  [8-1:3] ? {  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  [8-1:3],3'b000}:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  [2] ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre  [0] ? 'd1:'d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready_pre  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_remain  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_release_fifo  );


    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_delay_fifo_not_ready_dout;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_last  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d2  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d3  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_req_in_prog  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                else
                    if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_buffer_small  ))
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b1;
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_in_prog  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready_pre  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_wait  |(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_page_cross  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size  !=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  )))
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=1'b0;
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready   <=|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size   <={8{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_req_in_prog  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_CMD_SIZE  ;
            else
                if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_size  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_buffer_small  ))
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_size  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_update  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d2  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush_in  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg   <=2'b00;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_in  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg  [0] ? 2'b11:2'b01;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush_in  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_start  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b0;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_in  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg   <=1'b1;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_reg  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [2:0]==3'd0 ? 4'd8:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [1:0]==2'd0 ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [0]==1'd0 ? 'd2:'d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_size  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [0] ? 'd1:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [1] ? 'd2:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr  [2]&(!0) ? 'd4:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req  [1] ? 'd32:'d16;


    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps  ;
    reg[2:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  )&(|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size  >  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain  )|(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain  <'d8);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=1'b0;
        else
            if ((  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end  ))
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=1'b0;
            else
                if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end  )&(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out_pre  ;

    always @(               dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush                                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready                     or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain                    or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready                   or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small                  or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross                 or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr               or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out             or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush   =1'b0;
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE  )
                                begin
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b1;
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                                end
                                else
                                begin
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                                end
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr  )
                    begin
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
                    end
                    else
                    begin
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                    end
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS  ;
                else
                    if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b0;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK  ;
                        end
                        else
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
                    else
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_WRITE  )
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req   =1'b1;
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        end
                        else
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READ  )
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_RECHK  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  )
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait   =1'b1;
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY_OUT  ;
                end
                else
                    if ((~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  )|(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in  )|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_READY  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS   :
            begin
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty  )
                    begin
                        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain  <='d16))
                        begin
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain  =='d0)
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ  ;
                            else
                                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
                        end
                        else
                            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
                    end
                    else
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_CROSS  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_BURST_REQ   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req   =1'b1;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_REQ_LINE  ;
            end
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH   :
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush   =1'b1;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_FLUSH  ;
            end
            default :
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_IDLE  ;
            else
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ps   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ns  ;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size_pre2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_not_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_wait = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_buffer_small = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_ch_end_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_size_pre2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size_pre2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_not_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_not_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_line_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_burst_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_wait = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_wait;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_buffer_small = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_dma_axi64_core0_ch_calc_joint_joint_buffer_small;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_release_fifo  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_in  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_out  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_cross  );
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_update_d3 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update_d3;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_ch_end_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_burst_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_line_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_burst_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_dma_axi64_ch_calc_size_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d2 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d2;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_update_d3 = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update_d3;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_ch_end_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_burst_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_line_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_burst_req_in;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_burst_req_out = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_burst_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_dma_axi64_ch_calc_size_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush_in;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_load_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_ch_end_flush = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_wr_cmd_pending = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_frame_width = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_frame_width;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size[8-1:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_gap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_burst_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_line_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_in = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_burst_req = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_burst_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_rd_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_req_in_prog = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_load_addr = {32{1'b0}};
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_ch_end_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ch_end;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_outs_empty = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_outs_empty;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_max_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_max_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_start_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_start_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_frame_width = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_frame_width;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_x_size[8-1:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_x_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_x_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_wr_ready = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_fifo_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_fullness;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_last = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_last;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_burst_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_single = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_single;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_ready_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_joint_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_in = 1'b0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_line_req = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_burst_req_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_burst_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_line_req_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_cross = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_joint_flush = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_calc_wr_joint_flush_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_flush;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_wait_ready  =1'b1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_wait_ready  =1'b1;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clken;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req;
    reg [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready;
    wire [4:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clken;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req;
    reg [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready;
    wire [4:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_num;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr;

    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req_full  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready_pre  ;
    always @(      dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clken                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr_valid           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_num   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_clr   ={31{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_clr   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_num  ]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr_valid  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clken  ;
    end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req_full  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req  ,1'b1};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req_full  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_num  ];

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_DELAY  -1];




    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req_full  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready_pre  ;
    always @(      dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clken                or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr_valid           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_num   )
    begin
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_clr   ={31{1'b0}};
        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_clr   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_num  ]=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr_valid  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clken  ;
    end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req_full  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req  ,1'b1};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req_full  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_num  ];


    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_delay_ready_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_delay_ready_dout;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clken = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_req = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_periph_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_gclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clken = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_req = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_periph_num = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_periph_mux_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_mux;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_reset;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_end_swap;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wsize;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_align;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rsize;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_align;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_single;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_burst_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_clr_line;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_overflow;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_underflow;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_fifo  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_ptr  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_bsel  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wdata  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wsize  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rdata  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rsize  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_ptr  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_valid  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_ptr  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_ptr  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_line_remain  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_joint_delay  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_DOUT  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_d  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_valid  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata_valid  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rdata  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rdata  &{64{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_valid  }};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_valid  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wsize;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align;
    wire [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_incr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_end_swap;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_fifo;
    reg [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr;
    reg [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel;
    reg [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize;

    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append_wsize  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_direct_wsize  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  ;
    wire[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align_valid  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  ;
    reg[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_pre  ;
    wire[8-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_swap  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre_d  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_swap  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain   <=4'd8;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_clr_line  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain   <=4'd8;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain   <=4'd8;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size  +  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wsize  ;

    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_min;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_min;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_b  ;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_b  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_b = 4'd8;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_append_min;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_line_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_direct_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_min2_direct_min;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   <=1'b0;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   <=1'b0;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   <=1'b1;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size   <={4{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append_wsize  ;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_join_wsize  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_direct_wsize  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d   <={64{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align_valid  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_incr   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr  [3-1:0];
    always @(     dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align_valid           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align_valid  [3-1:0])
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:8]};
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [15:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:16]};
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [23:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:24]};
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [31:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:32]};
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [39:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:40]};
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [47:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:48]};
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [55:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata  [63:56]};
        endcase
    end

    always @(     dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size  [3-1:0])
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:8],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [7:0]};
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [15:0]};
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:24],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [23:0]};
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:32],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [31:0]};
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:40],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [39:0]};
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:48],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [47:0]};
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  [63:56],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata_d  [55:0]};
        endcase
    end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd1 ? 8'b00000001:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd2 ? 8'b00000011:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd3 ? 8'b00000111:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd4 ? 8'b00001111:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd5 ? 8'b00011111:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd6 ? 8'b00111111:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd7 ? 8'b01111111:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize  ==4'd8 ? 8'b11111111:{8{1'b0}};
    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr  [3-1:0])
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  ;
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [6:0],1'b0};
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [5:0],2'b0};
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [4:0],3'b0};
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [3:0],4'b0};
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [2:0],5'b0};
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [1:0],6'b0};
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_dec  [0],7'b0};
        endcase
    end

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  )&(|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wr   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_size  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append_wsize  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_direct_wsize  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_append   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_next_wdata  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_align_wdata  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_bsel_shift  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr0_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_fifo = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_delay_wr_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize   <={4{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre_d   <={64{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_pre  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize_pre  ;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre_d   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre  ;
            end


    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap;
    wire [63:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in;
    wire [63:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out;

    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_low  ;
    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_high  ;
    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_low  ;
    wire[31:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_high  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_low  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_high  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_low  ;
    wire[3:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_high  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_low  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap  ==2'b11 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in  [63:32]:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in  [31:0];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_high  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap  ==2'b11 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in  [31:0]:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in  [63:32];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_low  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap  ==2'b11 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in  [7:4]:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in  [3:0];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_high  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap  ==2'b11 ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in  [3:0]:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in  [7:4];

    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in;
    reg [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out;
    wire [3:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in;
    reg [3:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in;
    reg [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out;
    wire [3:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in;
    reg [3:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out;

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap  [1:0])
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  ;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [31:24],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [15:8]};
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [15:8],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [31:24]};
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [15:8],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in  [31:24]};
        endcase
    end

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap  [1:0])
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  ;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [3],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [1]};
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [1],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [3]};
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [1],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in  [3]};
        endcase
    end




    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap  [1:0])
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  ;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [31:24],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [15:8]};
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [15:8],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [31:24]};
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [15:8],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [23:16],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in  [31:24]};
        endcase
    end

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap  [1:0])
            2 'b00:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  ;
            2 'b01:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [3],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [1]};
            2 'b10:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [1],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [3]};
            2 'b11:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [1],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [2],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in  [3]};
        endcase
    end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_low;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_low = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_data_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_low;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_low = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_low_bsel_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in_high;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_high = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_data_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in_high;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_high = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_swap32_high_bsel_out;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_high  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out_low  };
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out  ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_high  ,  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out_low  };
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_end_swap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_pre_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_data_out;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_in = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_swap64_bsel_out;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata   <={64{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr   <={5{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel   <={8{1'b0}};
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata_swap  ;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr_pre  ;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel_swap  ;
            end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_wr_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_rd_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_end_swap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_fifo = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wr_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_bsel = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_bsel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_wr_slicer_slice_wsize;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rsize;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align;
    wire [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_ptr;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_line_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_single;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd;
    reg [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rsize;
    wire [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_ptr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_valid;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd_d  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_d  ;
    wire[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid_pre  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid  ;
    reg[3-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_d  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre  ;
    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize_pre  ;
    reg[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize_reg  ;
    wire[4-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rd  ;

    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_dout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_DELAY  -1];



    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd0_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd_d;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd_valid_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_pre;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd1_dout;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_delay_fifo_rd2_dout;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid_pre  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_incr  )&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_single   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_ptr  [3-1:0]:  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid   <={3{1'b0}};
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_d   <={3{1'b0}};
        end
        else
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid_pre  ;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_d   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid  ;
        end

    always @(     dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata              or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata           or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_d   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_d  [3-1:0])
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [63:0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [55:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [7:0]};
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [47:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [15:0]};
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [39:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [23:0]};
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [31:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [31:0]};
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [23:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [39:0]};
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [15:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [47:0]};
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata   ={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [7:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata  [55:0]};
        endcase
    end

    always @(    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata            or    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid   )
    begin
        case (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align_valid  [3-1:0])
            3 'd0:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:0];
            3 'd1:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{56{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:56]};
            3 'd2:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{48{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:48]};
            3 'd3:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{40{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:40]};
            3 'd4:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{32{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:32]};
            3 'd5:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{24{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:24]};
            3 'd6:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{16{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:16]};
            3 'd7:
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre   ={{8{1'b0}},  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata  [63:8]};
        endcase
    end

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata   <={64{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_d  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rdata_pre  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  +({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rsize  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  |(|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  ))
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize_pre  ;


    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_a;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_b;
    wire [ dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_WIDTH -1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_min;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_min  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_a  <  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_b   ?   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_a  :  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_b  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_a = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_line_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_b = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_actual_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_min_rsize_min;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize_reg   <={4{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rd  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize_reg   <={4{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  +({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rsize  );

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize_reg  -({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd_d  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rsize  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rd  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  )&(|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rsize  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_next_rd  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_ptr  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_ptr  ;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_DOUT;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_rd_line_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_line_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_wr_single = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_single;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_rd_slicer_slice_rd_valid;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_outstanding;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr_fifo;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_clr_line;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_next_size;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_burst_size;
    reg [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr;
    reg [5-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr;
    reg [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_wr_ready;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow;

    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr_pre  ;
    wire[5-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr_pre  ;
    wire[5+1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness_pre  ;
    reg[5+1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog_d  ;
    reg  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay_reg  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow_pre  ;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow_pre  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr  +({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wsize  );
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr  +({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rsize  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr   <={5{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr   <={5{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr   <={5{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr   <={5{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr_pre  ;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain   <=4'd8;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_clr_line  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain   <=4'd8;
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd  &(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain  ==  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rsize  ))
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain   <=4'd8;
                else
                    if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd  )
                        dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain  -  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rsize  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  +({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wsize  )-({4{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rd  }}&  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rsize  );
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness   <={5+2{1'b0}};
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness   <={5+2{1'b0}};
            else
                if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rd  |  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness_pre  ;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_din;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_dout;

    reg[  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_DELAY  :0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_shift_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_DELAY  +1{1'b0}};
        else
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_shift_reg   <={  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_DELAY  -1:0],  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_din  };

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_dout  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_shift_reg  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_DELAY  -1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_din = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog_d = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_delay_joint_in_prog_dout;

    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay_reg   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog  &(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog_d  ))
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay_reg   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  >32-4'd8;
            else
                if (~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay_reg   <=1'b0;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay_reg  ;
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_wr_ready   <=1'b0;
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog  )
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_wr_ready   <=1'b0;
            else
                if (|  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_next_size  )
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_wr_ready   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness_pre  >=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_next_size  ;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow_pre  =  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  [5+1];
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow_pre  =(~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  [5+1])&(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fullness  [5:0]>32);
    always @(  posedge    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk          or  posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset  )
        begin
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow   <=1'b0;
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow   <=1'b0;
        end
        else
            if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update  )
            begin
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow   <=1'b0;
                dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow   <=1'b0;
            end
            else
                if ((!  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow  )&(!  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow  ))
                begin
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow_pre  ;
                    dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow_pre  ;
                end

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wr_fifo = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_slice_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_ptr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_wr_ptr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_line_remain = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_rd_line_remain;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_joint_delay = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_joint_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_overflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_overflow;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_underflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_ptr_fifo_underflow;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_CLK;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD;
    wire [5-3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR_ADDR;
    wire [5-3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD_ADDR;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL;
    reg [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DOUT;

    reg[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_Mem  [4-1:0];
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BitSEL  ;
    wire[64-1:0]  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN_BitSEL  ;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BitSEL  ={{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [7]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [6]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [5]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [4]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [3]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [2]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [1]}},{8{  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL  [0]}}};
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN_BitSEL  =(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_Mem  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR_ADDR  ]&~  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BitSEL  )|(  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN  &  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BitSEL  );
    always @( posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_CLK  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_Mem   [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR_ADDR  ]<=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN_BitSEL  ;

    always @( posedge   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_CLK  )
        if (  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD  )
            dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DOUT   <=  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_Mem  [  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD_ADDR  ];

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_CLK = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_fifo;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_WR_ADDR = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wr_ptr[5-1:3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_RD_ADDR = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_rd_ptr[5-1:3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DIN = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_BSEL = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_slice_bsel;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_DOUT = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_dma_axi64_ch_fifo_DOUT;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_clk = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_reset = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_end_swap = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_end_swap;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_outstanding = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_outstanding;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_ch_update = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_update;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_align = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_align;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_incr = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_incr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_single = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_single;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_overflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_overflow;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_underflow = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_dma_axi64_ch_fifo_ctrl_fifo_underflow;

    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*0:32*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*0+31-1:31*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*0+31-1:31*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*0):1*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*0:32*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*0:8*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*0:6*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*0:3*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*0:32*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*0:8*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*0:6*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*0:3*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*0:64*0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[0];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[0] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch0_joint_req;


    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_req;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_clk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_reset;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_scan_en;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pclk;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_clken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pclken;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_psel;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_penable;
    wire [7:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_paddr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pwrite;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pwdata;
    wire [31:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_prdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pslverr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_tx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_tx_clr;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_rx_req;
    wire [31:1] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_rx_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_cmd_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_load;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_cmd_split;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_cmd_pending;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_last;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_slverr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_decerr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wr;
    wire [1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wr_cycle;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_req_in_prog;
    wire [1-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_int_all_proc;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_start;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_idle;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_rd_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_wr_active;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_last_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_line_cmd;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_go_next_line;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_transfer_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_start;
    wire [32-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_addr;
    wire [8-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_size;
    wire [6-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_tokens;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_port_num;
    wire [3-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_periph_delay;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_valid;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_transfer;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_transfer_size;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_next_size;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_stall;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_incr;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_aw;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_w;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_ar;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wdt_timeout;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wr;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wdata;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rd;
    wire [4-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rsize;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rd_valid;
    wire [64-1:0] dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rdata;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wr_ready;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_mode;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_remote;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_page_cross;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_not_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_mux_in_prog;
    wire  dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_req;

    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_req  ='d0;



    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_prdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pslverr  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_tx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_rx_clr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_req_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_int_all_proc  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_idle  ='d1;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_rd_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_wr_active  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_last_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_line_cmd  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_go_next_line  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_addr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_size  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_tokens  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_port_num  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_periph_delay  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_stall  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_incr  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rd_valid  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rdata  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wr_ready  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_not_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_mux_in_prog  ='d0;
    assign   dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_req  ='d0;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*1:32*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*1+31-1:31*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*1+31-1:31*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*1):1*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*1:32*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*1:8*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*1:6*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*1:3*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*1:32*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*1:8*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*1:6*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*1:3*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*1:64*1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[1];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[1] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty1_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*2:32*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*2+31-1:31*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*2+31-1:31*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*2):1*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*2:32*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*2:8*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*2:6*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*2:3*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*2:32*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*2:8*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*2:6*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*2:3*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*2:64*2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[2];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[2] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty2_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*3:32*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*3+31-1:31*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*3+31-1:31*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*3):1*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*3:32*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*3:8*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*3:6*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*3:3*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*3:32*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*3:8*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*3:6*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*3:3*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*3:64*3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[3];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[3] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty3_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*4:32*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*4+31-1:31*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*4+31-1:31*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*4):1*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*4:32*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*4:8*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*4:6*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*4:3*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*4:32*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*4:8*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*4:6*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*4:3*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*4:64*4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[4];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[4] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty4_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*5:32*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*5+31-1:31*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*5+31-1:31*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*5):1*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*5:32*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*5:8*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*5:6*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*5:3*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*5:32*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*5:8*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*5:6*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*5:3*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*5:64*5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[5];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[5] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty5_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*6:32*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*6+31-1:31*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*6+31-1:31*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*6):1*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*6:32*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*6:8*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*6:6*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*6:3*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*6:32*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*6:8*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*6:6*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*6:3*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*6:64*6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[6];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[6] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty6_joint_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_clk = dma_axi64_core0_dma_axi64_core0_channels_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_reset = dma_axi64_core0_dma_axi64_core0_channels_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_scan_en = dma_axi64_core0_dma_axi64_core0_channels_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pclk = dma_axi64_core0_dma_axi64_core0_channels_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_clken = dma_axi64_core0_dma_axi64_core0_channels_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pclken = dma_axi64_core0_dma_axi64_core0_channels_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_psel = dma_axi64_core0_dma_axi64_core0_channels_ch_psel[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_penable = dma_axi64_core0_dma_axi64_core0_channels_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_paddr = dma_axi64_core0_dma_axi64_core0_channels_paddr[7:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pwrite = dma_axi64_core0_dma_axi64_core0_channels_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pwdata = dma_axi64_core0_dma_axi64_core0_channels_pwdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_prdata[31+32*7:32*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_prdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_pslverr[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_tx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_tx_clr[31*7+31-1:31*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_rx_req = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_periph_rx_clr[31*7+31-1:31*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_periph_rx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_split[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_cmd_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_cmd_line[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_line[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_load = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_load[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_slverr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_decerr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_cmd_split = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_split[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_cmd_pending = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_cmd_pending[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_line = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_line[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_last = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_last[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_slverr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_slverr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_decerr = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_decerr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_load_wr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wr_cycle = dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_wdata = dma_axi64_core0_dma_axi64_core0_channels_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_load_req_in_prog[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc[1-1+(1*7):1*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_start = dma_axi64_core0_dma_axi64_core0_channels_ch_start[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_idle[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_idle;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_active[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_rd_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_ch_wr_active;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_last_cmd[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_line_cmd[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_line_cmd[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_line_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_go_next_line[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_go_next_line[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_start[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_addr[32-1+32*7:32*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_burst_size[8-1+8*7:8*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_tokens[6-1+6*7:6*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_port_num[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_periph_delay[3-1+3*7:3*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_valid[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_transfer[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_rd_clr_stall[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_start = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_start[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_addr[32-1+32*7:32*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_addr;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_burst_size[8-1+8*7:8*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_burst_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_tokens[6-1+6*7:6*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_tokens;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_port_num[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_port_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_periph_delay[3-1+3*7:3*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_valid[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_transfer = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_transfer[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_transfer_size = dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_next_size = dma_axi64_core0_dma_axi64_core0_channels_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_wr_clr_stall[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_aw = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_aw[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_w = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_w[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_timeout_ar = dma_axi64_core0_dma_axi64_core0_channels_ch_timeout_ar[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wdt_timeout = dma_axi64_core0_dma_axi64_core0_channels_ch_wdt_timeout[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wr = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rd = dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rsize = dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_valid[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rd_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rdata[(64-1)+64*7:64*7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_rdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_ready[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_fifo_wr_ready;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_mode = dma_axi64_core0_dma_axi64_core0_channels_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_remote = dma_axi64_core0_dma_axi64_core0_channels_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_rd_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_page_cross[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_wr_page_cross = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_page_cross[7];
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_in_prog[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_not_in_prog[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_not_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_mux_in_prog[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_mux_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req[7] = dma_axi64_core0_dma_axi64_core0_channels_dma_axi64_core0_ch_empty7_joint_req;

    assign dma_axi64_core0_dma_axi64_core0_channels_clk = dma_axi64_core0_clk;
    assign dma_axi64_core0_dma_axi64_core0_channels_reset = dma_axi64_core0_reset;
    assign dma_axi64_core0_dma_axi64_core0_channels_scan_en = dma_axi64_core0_scan_en;
    assign dma_axi64_core0_dma_axi64_core0_channels_pclk = dma_axi64_core0_pclk;
    assign dma_axi64_core0_dma_axi64_core0_channels_clken = dma_axi64_core0_clken;
    assign dma_axi64_core0_dma_axi64_core0_channels_pclken = dma_axi64_core0_pclken;
    assign dma_axi64_core0_dma_axi64_core0_channels_psel = dma_axi64_core0_psel;
    assign dma_axi64_core0_dma_axi64_core0_channels_penable = dma_axi64_core0_penable;
    assign dma_axi64_core0_dma_axi64_core0_channels_paddr = dma_axi64_core0_paddr[10:0];
    assign dma_axi64_core0_dma_axi64_core0_channels_pwrite = dma_axi64_core0_pwrite;
    assign dma_axi64_core0_dma_axi64_core0_channels_pwdata = dma_axi64_core0_pwdata;
    assign dma_axi64_core0_prdata = dma_axi64_core0_dma_axi64_core0_channels_prdata;
    assign dma_axi64_core0_pslverr = dma_axi64_core0_dma_axi64_core0_channels_pslverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_periph_tx_req = dma_axi64_core0_periph_tx_req;
    assign dma_axi64_core0_periph_tx_clr = dma_axi64_core0_dma_axi64_core0_channels_periph_tx_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_periph_rx_req = dma_axi64_core0_periph_rx_req;
    assign dma_axi64_core0_periph_rx_clr = dma_axi64_core0_dma_axi64_core0_channels_periph_rx_clr;
    assign dma_axi64_core0_rd_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_rd_clr_valid;
    assign dma_axi64_core0_wr_clr_valid = dma_axi64_core0_dma_axi64_core0_channels_wr_clr_valid;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr = dma_axi64_core0_rd_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr_load = dma_axi64_core0_rd_clr_load;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr = dma_axi64_core0_wr_clr;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_split = dma_axi64_core0_rd_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_line = dma_axi64_core0_rd_cmd_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_num = dma_axi64_core0_rd_cmd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_split = dma_axi64_core0_wr_cmd_split;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_pending = dma_axi64_core0_wr_cmd_pending;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_num = dma_axi64_core0_wr_cmd_num;
    assign dma_axi64_core0_rd_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_rd_clr_stall;
    assign dma_axi64_core0_wr_clr_stall = dma_axi64_core0_dma_axi64_core0_channels_wr_clr_stall;
    assign dma_axi64_core0_dma_axi64_core0_channels_load_wr = dma_axi64_core0_load_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_load_wr_num = dma_axi64_core0_load_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_load_wr_cycle = dma_axi64_core0_load_wr_cycle;
    assign dma_axi64_core0_dma_axi64_core0_channels_load_wdata = dma_axi64_core0_load_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num = dma_axi64_core0_rd_ch_num;
    assign dma_axi64_core0_load_req_in_prog = dma_axi64_core0_dma_axi64_core0_channels_load_req_in_prog;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num = dma_axi64_core0_wr_ch_num_joint;
    assign dma_axi64_core0_wr_last_cmd = dma_axi64_core0_dma_axi64_core0_channels_wr_last_cmd;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_slverr = dma_axi64_core0_rd_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_decerr = dma_axi64_core0_rd_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_slverr = dma_axi64_core0_wr_slverr;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_decerr = dma_axi64_core0_wr_decerr;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_ch_num_resp = dma_axi64_core0_rd_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_ch_num_resp = dma_axi64_core0_wr_ch_num_resp;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr_last = dma_axi64_core0_wr_clr_last;
    assign dma_axi64_core0_ch_int_all_proc = dma_axi64_core0_dma_axi64_core0_channels_ch_int_all_proc;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_start = dma_axi64_core0_ch_start;
    assign dma_axi64_core0_ch_idle = dma_axi64_core0_dma_axi64_core0_channels_ch_idle;
    assign dma_axi64_core0_ch_active = dma_axi64_core0_dma_axi64_core0_channels_ch_active;
    assign dma_axi64_core0_ch_rd_active = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_active;
    assign dma_axi64_core0_ch_wr_active = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_active;
    assign dma_axi64_core0_rd_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_rd_line_cmd;
    assign dma_axi64_core0_wr_line_cmd = dma_axi64_core0_dma_axi64_core0_channels_wr_line_cmd;
    assign dma_axi64_core0_rd_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_rd_go_next_line;
    assign dma_axi64_core0_wr_go_next_line = dma_axi64_core0_dma_axi64_core0_channels_wr_go_next_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_aw = dma_axi64_core0_timeout_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_w = dma_axi64_core0_timeout_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_ar = dma_axi64_core0_timeout_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_num_aw = dma_axi64_core0_timeout_num_aw;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_num_w = dma_axi64_core0_timeout_num_w;
    assign dma_axi64_core0_dma_axi64_core0_channels_timeout_num_ar = dma_axi64_core0_timeout_num_ar;
    assign dma_axi64_core0_dma_axi64_core0_channels_wdt_timeout = dma_axi64_core0_wdt_timeout;
    assign dma_axi64_core0_dma_axi64_core0_channels_wdt_ch_num = dma_axi64_core0_wdt_ch_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_wr_num = dma_axi64_core0_ch_fifo_wr_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_num = dma_axi64_core0_rd_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_burst_start = dma_axi64_core0_rd_burst_start;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_transfer = dma_axi64_core0_rd_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_transfer_size = dma_axi64_core0_rd_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line = dma_axi64_core0_rd_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_clr_line_num = dma_axi64_core0_rd_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_rd = dma_axi64_core0_ch_fifo_rd;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_rsize = dma_axi64_core0_ch_fifo_rsize;
    assign dma_axi64_core0_ch_fifo_rd_valid = dma_axi64_core0_dma_axi64_core0_channels_fifo_rd_valid;
    assign dma_axi64_core0_ch_fifo_rdata = dma_axi64_core0_dma_axi64_core0_channels_fifo_rdata;
    assign dma_axi64_core0_ch_fifo_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_fifo_wr_ready;
    assign dma_axi64_core0_ch_rd_ready = dma_axi64_core0_dma_axi64_core0_channels_ch_rd_ready;
    assign dma_axi64_core0_rd_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_rd_burst_addr;
    assign dma_axi64_core0_rd_burst_size = dma_axi64_core0_dma_axi64_core0_channels_rd_burst_size;
    assign dma_axi64_core0_rd_tokens = dma_axi64_core0_dma_axi64_core0_channels_rd_tokens;
    assign dma_axi64_core0_rd_cmd_port = dma_axi64_core0_dma_axi64_core0_channels_rd_cmd_port;
    assign dma_axi64_core0_rd_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_rd_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_ch_fifo_rd_num = dma_axi64_core0_ch_fifo_rd_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_num = dma_axi64_core0_wr_transfer_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_burst_start = dma_axi64_core0_wr_burst_start_joint;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_transfer = dma_axi64_core0_wr_transfer;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_transfer_size = dma_axi64_core0_wr_transfer_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_next_size = dma_axi64_core0_wr_next_size;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line = dma_axi64_core0_wr_clr_line;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_clr_line_num = dma_axi64_core0_wr_clr_line_num;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_wr = dma_axi64_core0_ch_fifo_wr;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_wdata = dma_axi64_core0_ch_fifo_wdata;
    assign dma_axi64_core0_dma_axi64_core0_channels_fifo_wsize = dma_axi64_core0_ch_fifo_wsize;
    assign dma_axi64_core0_ch_wr_ready = dma_axi64_core0_dma_axi64_core0_channels_ch_wr_ready;
    assign dma_axi64_core0_wr_burst_addr = dma_axi64_core0_dma_axi64_core0_channels_wr_burst_addr;
    assign dma_axi64_core0_wr_burst_size = dma_axi64_core0_dma_axi64_core0_channels_wr_burst_size;
    assign dma_axi64_core0_wr_tokens = dma_axi64_core0_dma_axi64_core0_channels_wr_tokens;
    assign dma_axi64_core0_wr_cmd_port = dma_axi64_core0_dma_axi64_core0_channels_wr_cmd_port;
    assign dma_axi64_core0_wr_periph_delay = dma_axi64_core0_dma_axi64_core0_channels_wr_periph_delay;
    assign dma_axi64_core0_dma_axi64_core0_channels_joint_mode = dma_axi64_core0_joint_mode;
    assign dma_axi64_core0_dma_axi64_core0_channels_joint_remote = dma_axi64_core0_joint_remote;
    assign dma_axi64_core0_dma_axi64_core0_channels_rd_page_cross = dma_axi64_core0_rd_page_cross;
    assign dma_axi64_core0_dma_axi64_core0_channels_wr_page_cross = dma_axi64_core0_wr_page_cross;
    assign dma_axi64_core0_joint_in_prog = dma_axi64_core0_dma_axi64_core0_channels_joint_in_prog;
    assign dma_axi64_core0_joint_not_in_prog = dma_axi64_core0_dma_axi64_core0_channels_joint_not_in_prog;
    assign dma_axi64_core0_joint_mux_in_prog = dma_axi64_core0_dma_axi64_core0_channels_joint_mux_in_prog;
    assign dma_axi64_core0_ch_joint_req = dma_axi64_core0_dma_axi64_core0_channels_ch_joint_req;

    assign dma_axi64_core0_clk = clk_out;
    assign dma_axi64_core0_reset = reset;
    assign dma_axi64_core0_scan_en = scan_en;
    assign idle = dma_axi64_core0_idle;
    assign ch_int_all_proc = dma_axi64_core0_ch_int_all_proc;
    assign dma_axi64_core0_ch_start = ch_start;
    assign dma_axi64_core0_periph_tx_req = periph_tx_req;
    assign periph_tx_clr = dma_axi64_core0_periph_tx_clr;
    assign dma_axi64_core0_periph_rx_req = periph_rx_req;
    assign periph_rx_clr = dma_axi64_core0_periph_rx_clr;
    assign dma_axi64_core0_pclk = clk;
    assign dma_axi64_core0_clken = clken;
    assign dma_axi64_core0_pclken = pclken;
    assign dma_axi64_core0_psel = psel;
    assign dma_axi64_core0_penable = penable;
    assign dma_axi64_core0_paddr = paddr[10:0];
    assign dma_axi64_core0_pwrite = pwrite;
    assign dma_axi64_core0_pwdata = pwdata;
    assign prdata = dma_axi64_core0_prdata;
    assign pslverr = dma_axi64_core0_pslverr;
    assign rd_port_num = dma_axi64_core0_rd_port_num;
    assign wr_port_num = dma_axi64_core0_wr_port_num;
    assign dma_axi64_core0_joint_mode_in = joint_mode;
    assign dma_axi64_core0_joint_remote = joint_remote;
    assign dma_axi64_core0_rd_prio_top = rd_prio_top;
    assign dma_axi64_core0_rd_prio_high = rd_prio_high;
    assign dma_axi64_core0_rd_prio_top_num = rd_prio_top_num;
    assign dma_axi64_core0_rd_prio_high_num = rd_prio_high_num;
    assign dma_axi64_core0_wr_prio_top = wr_prio_top;
    assign dma_axi64_core0_wr_prio_high = wr_prio_high;
    assign dma_axi64_core0_wr_prio_top_num = wr_prio_top_num;
    assign dma_axi64_core0_wr_prio_high_num = wr_prio_high_num;
    assign slow_AWADDR = dma_axi64_core0_AWADDR;
    assign slow_AWLEN = dma_axi64_core0_AWLEN;
    assign slow_AWSIZE = dma_axi64_core0_AWSIZE;
    assign slow_AWVALID = dma_axi64_core0_AWVALID;
    assign dma_axi64_core0_AWREADY = slow_AWREADY;
    assign slow_WDATA = dma_axi64_core0_WDATA;
    assign slow_WSTRB = dma_axi64_core0_WSTRB;
    assign slow_WLAST = dma_axi64_core0_WLAST;
    assign slow_WVALID = dma_axi64_core0_WVALID;
    assign dma_axi64_core0_WREADY = slow_WREADY;
    assign dma_axi64_core0_BRESP = slow_BRESP;
    assign dma_axi64_core0_BVALID = slow_BVALID;
    assign slow_BREADY = dma_axi64_core0_BREADY;
    assign slow_ARADDR = dma_axi64_core0_ARADDR;
    assign slow_ARLEN = dma_axi64_core0_ARLEN;
    assign slow_ARSIZE = dma_axi64_core0_ARSIZE;
    assign slow_ARVALID = dma_axi64_core0_ARVALID;
    assign dma_axi64_core0_ARREADY = slow_ARREADY;
    assign dma_axi64_core0_RDATA = slow_RDATA;
    assign dma_axi64_core0_RRESP = slow_RRESP;
    assign dma_axi64_core0_RLAST = slow_RLAST;
    assign dma_axi64_core0_RVALID = slow_RVALID;
    assign slow_RREADY = dma_axi64_core0_RREADY;

endmodule
