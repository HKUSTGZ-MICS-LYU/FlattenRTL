module RocketTile(
  input         clock,
                reset,
                auto_buffer_out_a_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_a_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_buffer_out_a_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_buffer_out_a_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [1:0]  auto_buffer_out_a_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_buffer_out_a_bits_address,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_a_bits_user_amba_prot_bufferable,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_modifiable,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_readalloc,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_writealloc,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_privileged,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_secure,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_a_bits_user_amba_prot_fetch,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [7:0]  auto_buffer_out_a_bits_mask,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [63:0] auto_buffer_out_a_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_a_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_b_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_b_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [2:0]  auto_buffer_out_b_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [1:0]  auto_buffer_out_b_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [3:0]  auto_buffer_out_b_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [1:0]  auto_buffer_out_b_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [31:0] auto_buffer_out_b_bits_address,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [7:0]  auto_buffer_out_b_bits_mask,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [63:0] auto_buffer_out_b_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_b_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_c_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_buffer_out_c_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_buffer_out_c_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [1:0]  auto_buffer_out_c_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_buffer_out_c_bits_address,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_c_bits_user_amba_prot_bufferable,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_modifiable,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_readalloc,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_writealloc,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_privileged,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_secure,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_c_bits_user_amba_prot_fetch,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [63:0] auto_buffer_out_c_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_c_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_d_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [2:0]  auto_buffer_out_d_bits_opcode,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [1:0]  auto_buffer_out_d_bits_param,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [3:0]  auto_buffer_out_d_bits_size,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [1:0]  auto_buffer_out_d_bits_source,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_d_bits_sink,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_bits_denied,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [63:0] auto_buffer_out_d_bits_data,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_buffer_out_d_bits_corrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_buffer_out_e_ready,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_buffer_out_e_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [1:0]  auto_buffer_out_e_bits_sink,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_broadcast_out_insns_0_valid,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [33:0] auto_broadcast_out_insns_0_iaddr,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_broadcast_out_insns_0_insn,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [2:0]  auto_broadcast_out_insns_0_priv,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_broadcast_out_insns_0_exception,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_broadcast_out_insns_0_interrupt,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [63:0] auto_broadcast_out_insns_0_cause,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [33:0] auto_broadcast_out_insns_0_tval,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [63:0] auto_broadcast_out_time,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_wfi_out_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_cease_out_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_halt_out_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_int_local_in_2_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_1_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_1_1,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_int_local_in_0_0,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_trace_core_source_out_group_0_iretire,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_trace_core_source_out_group_0_iaddr,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_trace_core_source_out_group_0_itype,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output        auto_trace_core_source_out_group_0_ilastsize,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [3:0]  auto_trace_core_source_out_priv,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  output [31:0] auto_trace_core_source_out_tval,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_trace_core_source_out_cause,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_nmi_in_rnmi,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input  [31:0] auto_nmi_in_rnmi_interrupt_vector,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_nmi_in_rnmi_exception_vector,	// src/main/scala/diplomacy/LazyModule.scala:374:18
                auto_reset_vector_in,	// src/main/scala/diplomacy/LazyModule.scala:374:18
  input         auto_hartid_in	// src/main/scala/diplomacy/LazyModule.scala:374:18
);

  wire [1:0]  buffer_auto_in_e_bits_sink;
  wire        buffer_auto_in_e_valid;
  wire        buffer_auto_in_e_ready;
  wire        buffer_auto_in_d_bits_corrupt;
  wire [63:0] buffer_auto_in_d_bits_data;
  wire        buffer_auto_in_d_bits_denied;
  wire [1:0]  buffer_auto_in_d_bits_sink;
  wire [1:0]  buffer_auto_in_d_bits_source;
  wire [3:0]  buffer_auto_in_d_bits_size;
  wire [1:0]  buffer_auto_in_d_bits_param;
  wire [2:0]  buffer_auto_in_d_bits_opcode;
  wire        buffer_auto_in_d_valid;
  wire        buffer_auto_in_d_ready;
  wire        buffer_auto_in_c_bits_corrupt;
  wire [63:0] buffer_auto_in_c_bits_data;
  wire        buffer_auto_in_c_bits_user_amba_prot_fetch;
  wire        buffer_auto_in_c_bits_user_amba_prot_secure;
  wire        buffer_auto_in_c_bits_user_amba_prot_privileged;
  wire        buffer_auto_in_c_bits_user_amba_prot_writealloc;
  wire        buffer_auto_in_c_bits_user_amba_prot_readalloc;
  wire        buffer_auto_in_c_bits_user_amba_prot_modifiable;
  wire        buffer_auto_in_c_bits_user_amba_prot_bufferable;
  wire [31:0] buffer_auto_in_c_bits_address;
  wire [1:0]  buffer_auto_in_c_bits_source;
  wire [3:0]  buffer_auto_in_c_bits_size;
  wire [2:0]  buffer_auto_in_c_bits_param;
  wire [2:0]  buffer_auto_in_c_bits_opcode;
  wire        buffer_auto_in_c_valid;
  wire        buffer_auto_in_c_ready;
  wire        buffer_auto_in_b_bits_corrupt;
  wire [63:0] buffer_auto_in_b_bits_data;
  wire [7:0]  buffer_auto_in_b_bits_mask;
  wire [31:0] buffer_auto_in_b_bits_address;
  wire [1:0]  buffer_auto_in_b_bits_source;
  wire [3:0]  buffer_auto_in_b_bits_size;
  wire [1:0]  buffer_auto_in_b_bits_param;
  wire [2:0]  buffer_auto_in_b_bits_opcode;
  wire        buffer_auto_in_b_valid;
  wire        buffer_auto_in_b_ready;
  wire        buffer_auto_in_a_bits_corrupt;
  wire [63:0] buffer_auto_in_a_bits_data;
  wire [7:0]  buffer_auto_in_a_bits_mask;
  wire        buffer_auto_in_a_bits_user_amba_prot_fetch;
  wire        buffer_auto_in_a_bits_user_amba_prot_secure;
  wire        buffer_auto_in_a_bits_user_amba_prot_privileged;
  wire        buffer_auto_in_a_bits_user_amba_prot_writealloc;
  wire        buffer_auto_in_a_bits_user_amba_prot_readalloc;
  wire        buffer_auto_in_a_bits_user_amba_prot_modifiable;
  wire        buffer_auto_in_a_bits_user_amba_prot_bufferable;
  wire [31:0] buffer_auto_in_a_bits_address;
  wire [1:0]  buffer_auto_in_a_bits_source;
  wire [3:0]  buffer_auto_in_a_bits_size;
  wire [2:0]  buffer_auto_in_a_bits_param;
  wire [2:0]  buffer_auto_in_a_bits_opcode;
  wire        buffer_auto_in_a_valid;
  wire        buffer_auto_in_a_ready;
  wire        widget_1_auto_in_d_ready;
  wire        widget_1_auto_in_a_bits_corrupt;
  wire [63:0] widget_1_auto_in_a_bits_data;
  wire [7:0]  widget_1_auto_in_a_bits_mask;
  wire        widget_1_auto_in_a_bits_user_amba_prot_fetch;
  wire        widget_1_auto_in_a_bits_user_amba_prot_secure;
  wire        widget_1_auto_in_a_bits_user_amba_prot_privileged;
  wire        widget_1_auto_in_a_bits_user_amba_prot_writealloc;
  wire        widget_1_auto_in_a_bits_user_amba_prot_readalloc;
  wire        widget_1_auto_in_a_bits_user_amba_prot_modifiable;
  wire        widget_1_auto_in_a_bits_user_amba_prot_bufferable;
  wire [31:0] widget_1_auto_in_a_bits_address;
  wire        widget_1_auto_in_a_bits_source;
  wire [3:0]  widget_1_auto_in_a_bits_size;
  wire [2:0]  widget_1_auto_in_a_bits_param;
  wire [2:0]  widget_1_auto_in_a_bits_opcode;
  wire        widget_1_auto_in_a_valid;
  wire [1:0]  widget_auto_in_e_bits_sink;
  wire        widget_auto_in_e_valid;
  wire        widget_auto_in_d_ready;
  wire        widget_auto_in_c_bits_corrupt;
  wire [63:0] widget_auto_in_c_bits_data;
  wire        widget_auto_in_c_bits_user_amba_prot_fetch;
  wire        widget_auto_in_c_bits_user_amba_prot_secure;
  wire        widget_auto_in_c_bits_user_amba_prot_privileged;
  wire        widget_auto_in_c_bits_user_amba_prot_writealloc;
  wire        widget_auto_in_c_bits_user_amba_prot_readalloc;
  wire        widget_auto_in_c_bits_user_amba_prot_modifiable;
  wire        widget_auto_in_c_bits_user_amba_prot_bufferable;
  wire [31:0] widget_auto_in_c_bits_address;
  wire        widget_auto_in_c_bits_source;
  wire [3:0]  widget_auto_in_c_bits_size;
  wire [2:0]  widget_auto_in_c_bits_param;
  wire [2:0]  widget_auto_in_c_bits_opcode;
  wire        widget_auto_in_c_valid;
  wire        widget_auto_in_b_ready;
  wire        widget_auto_in_a_bits_corrupt;
  wire [63:0] widget_auto_in_a_bits_data;
  wire [7:0]  widget_auto_in_a_bits_mask;
  wire        widget_auto_in_a_bits_user_amba_prot_fetch;
  wire        widget_auto_in_a_bits_user_amba_prot_secure;
  wire        widget_auto_in_a_bits_user_amba_prot_privileged;
  wire        widget_auto_in_a_bits_user_amba_prot_writealloc;
  wire        widget_auto_in_a_bits_user_amba_prot_readalloc;
  wire        widget_auto_in_a_bits_user_amba_prot_modifiable;
  wire        widget_auto_in_a_bits_user_amba_prot_bufferable;
  wire [31:0] widget_auto_in_a_bits_address;
  wire        widget_auto_in_a_bits_source;
  wire [3:0]  widget_auto_in_a_bits_size;
  wire [2:0]  widget_auto_in_a_bits_param;
  wire [2:0]  widget_auto_in_a_bits_opcode;
  wire        widget_auto_in_a_valid;
  wire [2:0]  broadcast_4_auto_in_0_action;
  wire        broadcast_4_auto_in_0_ivalid_0;
  wire        broadcast_4_auto_in_0_wvalid_0;
  wire        broadcast_4_auto_in_0_rvalid_0;
  wire        broadcast_4_auto_in_0_valid_0;
  wire        nexus_1_auto_out_stall;
  wire        nexus_1_auto_out_enable;
  wire [63:0] broadcast_3_auto_in_time;
  wire [33:0] broadcast_3_auto_in_insns_0_tval;
  wire [63:0] broadcast_3_auto_in_insns_0_cause;
  wire        broadcast_3_auto_in_insns_0_interrupt;
  wire        broadcast_3_auto_in_insns_0_exception;
  wire [2:0]  broadcast_3_auto_in_insns_0_priv;
  wire [31:0] broadcast_3_auto_in_insns_0_insn;
  wire [33:0] broadcast_3_auto_in_insns_0_iaddr;
  wire        broadcast_3_auto_in_insns_0_valid;
  wire [31:0] broadcast_2_auto_out_rnmi_exception_vector;
  wire [31:0] broadcast_2_auto_out_rnmi_interrupt_vector;
  wire        broadcast_2_auto_out_rnmi;
  wire [31:0] broadcast_2_auto_in_rnmi_exception_vector;
  wire [31:0] broadcast_2_auto_in_rnmi_interrupt_vector;
  wire        broadcast_2_auto_in_rnmi;
  wire [31:0] broadcast_1_auto_out_0;
  wire [31:0] broadcast_1_auto_in;
  wire        broadcast_auto_out;
  wire        broadcast_auto_in;
  wire        intSinkNodeIn_3;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_2;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_1;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        intSinkNodeIn_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeIn_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeIn_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeIn_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  tlOtherMastersNodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_auto_out_d_bits_corrupt;
  wire [63:0] widget_1_auto_out_d_bits_data;
  wire        widget_1_auto_out_d_bits_denied;
  wire [1:0]  widget_1_auto_out_d_bits_sink;
  wire        widget_1_auto_out_d_bits_source;
  wire [3:0]  widget_1_auto_out_d_bits_size;
  wire [1:0]  widget_1_auto_out_d_bits_param;
  wire [2:0]  widget_1_auto_out_d_bits_opcode;
  wire        widget_1_auto_out_d_valid;
  wire        widget_1_auto_out_a_ready;
  wire        widget_auto_out_e_ready;
  wire        widget_auto_out_d_bits_corrupt;
  wire [63:0] widget_auto_out_d_bits_data;
  wire        widget_auto_out_d_bits_denied;
  wire [1:0]  widget_auto_out_d_bits_sink;
  wire        widget_auto_out_d_bits_source;
  wire [3:0]  widget_auto_out_d_bits_size;
  wire [1:0]  widget_auto_out_d_bits_param;
  wire [2:0]  widget_auto_out_d_bits_opcode;
  wire        widget_auto_out_d_valid;
  wire        widget_auto_out_c_ready;
  wire        widget_auto_out_b_bits_corrupt;
  wire [63:0] widget_auto_out_b_bits_data;
  wire [7:0]  widget_auto_out_b_bits_mask;
  wire [31:0] widget_auto_out_b_bits_address;
  wire        widget_auto_out_b_bits_source;
  wire [3:0]  widget_auto_out_b_bits_size;
  wire [1:0]  widget_auto_out_b_bits_param;
  wire [2:0]  widget_auto_out_b_bits_opcode;
  wire        widget_auto_out_b_valid;
  wire        widget_auto_out_a_ready;
  wire        _core_io_imem_might_request;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_req_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [33:0] _core_io_imem_req_bits_pc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_req_bits_speculative;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_bits_rs1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_bits_rs2;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_sfence_bits_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_bits_asid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_bits_hv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_sfence_bits_hg;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_resp_ready;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_imem_btb_update_bits_prediction_cfiType;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_prediction_taken;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_imem_btb_update_bits_prediction_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_prediction_bridx;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_btb_update_bits_prediction_target;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_prediction_entry;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_imem_btb_update_bits_prediction_bht_history;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_prediction_bht_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_btb_update_bits_pc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_btb_update_bits_target;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_taken;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_btb_update_bits_isValid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_btb_update_bits_br_pc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_imem_btb_update_bits_cfiType;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_imem_bht_update_bits_prediction_history;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_bits_prediction_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_bht_update_bits_pc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_bits_branch;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_bits_taken;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_bht_update_bits_mispredict;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_ras_update_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_imem_ras_update_bits_cfiType;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_imem_ras_update_bits_returnAddr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_flush_icache;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_imem_progress;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [33:0] _core_io_dmem_req_bits_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [5:0]  _core_io_dmem_req_bits_tag;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [4:0]  _core_io_dmem_req_bits_cmd;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_dmem_req_bits_size;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_signed;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_dmem_req_bits_dprv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_dv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_phys;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_no_alloc;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_req_bits_no_xcpt;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_dmem_req_bits_data;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_dmem_req_bits_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_s1_kill;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_dmem_s1_data_data;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_dmem_s1_data_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_s2_kill;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_dmem_keep_clock_enabled;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [3:0]  _core_io_ptw_ptbr_mode;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [15:0] _core_io_ptw_ptbr_asid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [43:0] _core_io_ptw_ptbr_ppn;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [3:0]  _core_io_ptw_hgatp_mode;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [15:0] _core_io_ptw_hgatp_asid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [43:0] _core_io_ptw_hgatp_ppn;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [3:0]  _core_io_ptw_vsatp_mode;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [15:0] _core_io_ptw_vsatp_asid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [43:0] _core_io_ptw_vsatp_ppn;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_valid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_rs1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_rs2;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [32:0] _core_io_ptw_sfence_bits_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_asid;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_hv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_sfence_bits_hg;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_debug;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_cease;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_wfi;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_status_isa;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_dprv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_dv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_prv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_v;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_sd;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [22:0] _core_io_ptw_status_zero2;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mpv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_gva;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mbe;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_sbe;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_sxl;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_uxl;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_sd_rv32;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_ptw_status_zero1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_tsr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_tw;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_tvm;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mxr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_sum;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mprv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_xs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_fs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_mpp;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_status_vs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_spp;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mpie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_ube;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_spie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_upie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_mie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_hie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_sie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_status_uie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_hstatus_zero6;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_hstatus_vsxl;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [8:0]  _core_io_ptw_hstatus_zero5;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_vtsr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_vtw;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_vtvm;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_hstatus_zero3;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [5:0]  _core_io_ptw_hstatus_vgein;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_hstatus_zero2;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_hu;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_spvp;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_spv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_gva;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_hstatus_vsbe;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [4:0]  _core_io_ptw_hstatus_zero1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_debug;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_cease;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_wfi;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_gstatus_isa;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_dprv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_dv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_prv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_v;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_sd;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [22:0] _core_io_ptw_gstatus_zero2;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mpv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_gva;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mbe;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_sbe;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_sxl;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_uxl;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_sd_rv32;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [7:0]  _core_io_ptw_gstatus_zero1;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_tsr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_tw;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_tvm;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mxr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_sum;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mprv;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_xs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_fs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_mpp;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_gstatus_vs;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_spp;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mpie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_ube;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_spie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_upie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_mie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_hie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_sie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_gstatus_uie;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_0_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_0_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_0_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_0_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_0_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_1_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_1_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_1_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_1_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_1_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_2_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_2_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_2_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_2_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_2_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_3_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_3_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_3_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_3_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_3_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_4_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_4_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_4_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_4_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_4_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_5_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_5_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_5_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_5_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_5_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_6_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_6_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_6_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_6_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_6_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_l;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_7_cfg_res;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [1:0]  _core_io_ptw_pmp_7_cfg_a;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_x;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_w;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_pmp_7_cfg_r;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [29:0] _core_io_ptw_pmp_7_addr;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [31:0] _core_io_ptw_pmp_7_mask;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_0_ren;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_0_wen;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_0_wdata;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_0_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_1_ren;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_1_wen;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_1_wdata;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_1_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_2_ren;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_2_wen;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_2_wdata;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_2_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_3_ren;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_ptw_customCSRs_csrs_3_wen;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_3_wdata;	// src/main/scala/tile/RocketTile.scala:127:20
  wire [63:0] _core_io_ptw_customCSRs_csrs_3_value;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _core_io_wfi;	// src/main/scala/tile/RocketTile.scala:127:20
  wire        _ptw_io_requestor_0_req_ready;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_valid;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_ae_ptw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_ae_final;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_gf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_hx;	// src/main/scala/rocket/PTW.scala:801:19
  wire [9:0]  _ptw_io_requestor_0_resp_bits_pte_reserved_for_future;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_0_resp_bits_pte_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_resp_bits_pte_reserved_for_software;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_d;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_g;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_u;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_pte_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_resp_bits_level;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_fragmented_superpage;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_homogeneous;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_gpa_valid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [32:0] _ptw_io_requestor_0_resp_bits_gpa_bits;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_resp_bits_gpa_is_pte;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_0_ptbr_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_0_ptbr_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_0_ptbr_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_0_hgatp_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_0_hgatp_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_0_hgatp_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_0_vsatp_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_0_vsatp_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_0_vsatp_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_cease;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_wfi;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_status_isa;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_dprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_dv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_prv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_sd;	// src/main/scala/rocket/PTW.scala:801:19
  wire [22:0] _ptw_io_requestor_0_status_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mpv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_sbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_sxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_uxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_sd_rv32;	// src/main/scala/rocket/PTW.scala:801:19
  wire [7:0]  _ptw_io_requestor_0_status_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_tsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_tw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_tvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mxr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_sum;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_xs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_fs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_mpp;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_status_vs;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_spp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mpie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_ube;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_spie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_upie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_mie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_hie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_sie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_status_uie;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_hstatus_zero6;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_hstatus_vsxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [8:0]  _ptw_io_requestor_0_hstatus_zero5;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_vtsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_vtw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_vtvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_hstatus_zero3;	// src/main/scala/rocket/PTW.scala:801:19
  wire [5:0]  _ptw_io_requestor_0_hstatus_vgein;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_hstatus_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_hu;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_spvp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_spv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_hstatus_vsbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [4:0]  _ptw_io_requestor_0_hstatus_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_cease;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_wfi;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_gstatus_isa;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_dprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_dv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_prv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_sd;	// src/main/scala/rocket/PTW.scala:801:19
  wire [22:0] _ptw_io_requestor_0_gstatus_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mpv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_sbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_sxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_uxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_sd_rv32;	// src/main/scala/rocket/PTW.scala:801:19
  wire [7:0]  _ptw_io_requestor_0_gstatus_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_tsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_tw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_tvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mxr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_sum;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_xs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_fs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_mpp;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_gstatus_vs;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_spp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mpie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_ube;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_spie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_upie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_mie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_hie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_sie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_gstatus_uie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_0_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_0_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_0_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_0_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_0_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_1_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_1_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_1_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_1_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_1_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_2_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_2_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_2_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_2_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_2_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_3_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_3_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_3_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_3_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_3_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_4_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_4_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_4_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_4_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_4_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_5_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_5_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_5_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_5_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_5_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_6_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_6_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_6_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_6_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_6_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_7_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_0_pmp_7_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_pmp_7_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_0_pmp_7_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_0_pmp_7_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_0_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_0_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_0_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_0_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_1_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_1_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_1_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_1_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_2_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_2_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_2_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_2_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_3_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_0_customCSRs_csrs_3_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_3_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_0_customCSRs_csrs_3_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_req_ready;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_valid;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_ae_ptw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_ae_final;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_gf;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_hx;	// src/main/scala/rocket/PTW.scala:801:19
  wire [9:0]  _ptw_io_requestor_1_resp_bits_pte_reserved_for_future;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_1_resp_bits_pte_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_resp_bits_pte_reserved_for_software;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_d;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_g;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_u;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_pte_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_resp_bits_level;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_fragmented_superpage;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_homogeneous;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_gpa_valid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [32:0] _ptw_io_requestor_1_resp_bits_gpa_bits;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_resp_bits_gpa_is_pte;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_1_ptbr_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_1_ptbr_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_1_ptbr_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_1_hgatp_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_1_hgatp_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_1_hgatp_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire [3:0]  _ptw_io_requestor_1_vsatp_mode;	// src/main/scala/rocket/PTW.scala:801:19
  wire [15:0] _ptw_io_requestor_1_vsatp_asid;	// src/main/scala/rocket/PTW.scala:801:19
  wire [43:0] _ptw_io_requestor_1_vsatp_ppn;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_cease;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_wfi;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_status_isa;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_dprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_dv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_prv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_sd;	// src/main/scala/rocket/PTW.scala:801:19
  wire [22:0] _ptw_io_requestor_1_status_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mpv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_sbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_sxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_uxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_sd_rv32;	// src/main/scala/rocket/PTW.scala:801:19
  wire [7:0]  _ptw_io_requestor_1_status_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_tsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_tw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_tvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mxr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_sum;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_xs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_fs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_mpp;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_status_vs;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_spp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mpie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_ube;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_spie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_upie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_mie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_hie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_sie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_status_uie;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_hstatus_zero6;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_hstatus_vsxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [8:0]  _ptw_io_requestor_1_hstatus_zero5;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_vtsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_vtw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_vtvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_hstatus_zero3;	// src/main/scala/rocket/PTW.scala:801:19
  wire [5:0]  _ptw_io_requestor_1_hstatus_vgein;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_hstatus_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_hu;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_spvp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_spv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_hstatus_vsbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [4:0]  _ptw_io_requestor_1_hstatus_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_debug;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_cease;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_wfi;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_gstatus_isa;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_dprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_dv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_prv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_v;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_sd;	// src/main/scala/rocket/PTW.scala:801:19
  wire [22:0] _ptw_io_requestor_1_gstatus_zero2;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mpv;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_gva;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_sbe;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_sxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_uxl;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_sd_rv32;	// src/main/scala/rocket/PTW.scala:801:19
  wire [7:0]  _ptw_io_requestor_1_gstatus_zero1;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_tsr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_tw;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_tvm;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mxr;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_sum;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mprv;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_xs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_fs;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_mpp;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_gstatus_vs;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_spp;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mpie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_ube;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_spie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_upie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_mie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_hie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_sie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_gstatus_uie;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_0_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_0_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_0_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_0_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_0_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_1_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_1_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_1_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_1_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_1_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_2_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_2_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_2_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_2_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_2_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_3_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_3_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_3_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_3_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_3_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_4_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_4_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_4_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_4_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_4_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_5_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_5_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_5_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_5_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_5_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_6_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_6_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_6_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_6_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_6_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_l;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_7_cfg_res;	// src/main/scala/rocket/PTW.scala:801:19
  wire [1:0]  _ptw_io_requestor_1_pmp_7_cfg_a;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_x;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_w;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_pmp_7_cfg_r;	// src/main/scala/rocket/PTW.scala:801:19
  wire [29:0] _ptw_io_requestor_1_pmp_7_addr;	// src/main/scala/rocket/PTW.scala:801:19
  wire [31:0] _ptw_io_requestor_1_pmp_7_mask;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_0_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_0_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_0_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_0_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_1_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_1_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_1_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_1_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_2_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_2_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_2_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_2_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_3_ren;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_requestor_1_customCSRs_csrs_3_wen;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_3_wdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_requestor_1_customCSRs_csrs_3_value;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_perf_l2miss;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_perf_l2hit;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_perf_pte_miss;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_perf_pte_hit;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_0_stall;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_0_set;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_dpath_customCSRs_csrs_0_sdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_1_stall;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_1_set;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_dpath_customCSRs_csrs_1_sdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_2_stall;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_2_set;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_dpath_customCSRs_csrs_2_sdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_3_stall;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_customCSRs_csrs_3_set;	// src/main/scala/rocket/PTW.scala:801:19
  wire [63:0] _ptw_io_dpath_customCSRs_csrs_3_sdata;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _ptw_io_dpath_clock_enabled;	// src/main/scala/rocket/PTW.scala:801:19
  wire        _dcacheArb_io_requestor_0_req_ready;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_nack;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_nack_cause_raw;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_uncached;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [31:0] _dcacheArb_io_requestor_0_s2_paddr;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_valid;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [33:0] _dcacheArb_io_requestor_0_resp_bits_addr;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [5:0]  _dcacheArb_io_requestor_0_resp_bits_tag;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [4:0]  _dcacheArb_io_requestor_0_resp_bits_cmd;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_requestor_0_resp_bits_size;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_signed;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_requestor_0_resp_bits_dprv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_dv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_requestor_0_resp_bits_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [7:0]  _dcacheArb_io_requestor_0_resp_bits_mask;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_replay;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_resp_bits_has_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_requestor_0_resp_bits_data_word_bypass;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_requestor_0_resp_bits_data_raw;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_requestor_0_resp_bits_store_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_replay_next;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ma_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ma_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_pf_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_pf_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_gf_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_gf_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ae_ld;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_xcpt_ae_st;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [33:0] _dcacheArb_io_requestor_0_s2_gpa;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_s2_gpa_is_pte;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_ordered;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_acquire;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_release;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_grant;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_tlbMiss;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_blocked;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_requestor_0_clock_enabled;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_valid;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [33:0] _dcacheArb_io_mem_req_bits_addr;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [5:0]  _dcacheArb_io_mem_req_bits_tag;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [4:0]  _dcacheArb_io_mem_req_bits_cmd;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_mem_req_bits_size;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_signed;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [1:0]  _dcacheArb_io_mem_req_bits_dprv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_dv;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_phys;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_no_alloc;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_req_bits_no_xcpt;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_mem_req_bits_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [7:0]  _dcacheArb_io_mem_req_bits_mask;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_s1_kill;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [63:0] _dcacheArb_io_mem_s1_data_data;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire [7:0]  _dcacheArb_io_mem_s1_data_mask;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_s2_kill;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _dcacheArb_io_mem_keep_clock_enabled;	// src/main/scala/rocket/HellaCache.scala:286:25
  wire        _frontend_io_cpu_clock_enabled;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_btb_cfiType;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_taken;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_btb_mask;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_bridx;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [32:0] _frontend_io_cpu_resp_bits_btb_target;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_entry;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [7:0]  _frontend_io_cpu_resp_bits_btb_bht_history;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_btb_bht_value;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [33:0] _frontend_io_cpu_resp_bits_pc;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [31:0] _frontend_io_cpu_resp_bits_data;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [1:0]  _frontend_io_cpu_resp_bits_mask;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_pf_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_gf_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_xcpt_ae_inst;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_resp_bits_replay;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_gpa_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [33:0] _frontend_io_cpu_gpa_bits;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [33:0] _frontend_io_cpu_npc;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_perf_acquire;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_cpu_perf_tlbMiss;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_valid;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [20:0] _frontend_io_ptw_req_bits_bits_addr;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_need_gpa;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_vstage1;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_req_bits_bits_stage2;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_0_stall;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_0_set;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [63:0] _frontend_io_ptw_customCSRs_csrs_0_sdata;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_1_stall;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_1_set;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [63:0] _frontend_io_ptw_customCSRs_csrs_1_sdata;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_2_stall;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_2_set;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [63:0] _frontend_io_ptw_customCSRs_csrs_2_sdata;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_3_stall;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _frontend_io_ptw_customCSRs_csrs_3_set;	// src/main/scala/rocket/Frontend.scala:386:28
  wire [63:0] _frontend_io_ptw_customCSRs_csrs_3_sdata;	// src/main/scala/rocket/Frontend.scala:386:28
  wire        _dcache_io_cpu_req_ready;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_nack;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_nack_cause_raw;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_uncached;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [31:0] _dcache_io_cpu_s2_paddr;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_valid;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [33:0] _dcache_io_cpu_resp_bits_addr;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [5:0]  _dcache_io_cpu_resp_bits_tag;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [4:0]  _dcache_io_cpu_resp_bits_cmd;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [1:0]  _dcache_io_cpu_resp_bits_size;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_signed;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [1:0]  _dcache_io_cpu_resp_bits_dprv;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_dv;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_cpu_resp_bits_data;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [7:0]  _dcache_io_cpu_resp_bits_mask;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_replay;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_resp_bits_has_data;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_cpu_resp_bits_data_word_bypass;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_cpu_resp_bits_data_raw;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_cpu_resp_bits_store_data;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_replay_next;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ma_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ma_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_pf_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_pf_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_gf_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_gf_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ae_ld;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_xcpt_ae_st;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [33:0] _dcache_io_cpu_s2_gpa;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_s2_gpa_is_pte;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_ordered;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_acquire;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_release;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_grant;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_tlbMiss;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_blocked;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_canAcceptStoreThenLoad;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_canAcceptStoreThenRMW;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_canAcceptLoadThenLoad;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_storeBufferEmptyAfterLoad;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_perf_storeBufferEmptyAfterStore;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_cpu_clock_enabled;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_valid;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_valid;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [20:0] _dcache_io_ptw_req_bits_bits_addr;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_need_gpa;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_vstage1;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_req_bits_bits_stage2;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_0_stall;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_0_set;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_ptw_customCSRs_csrs_0_sdata;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_1_stall;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_1_set;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_ptw_customCSRs_csrs_1_sdata;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_2_stall;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_2_set;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_ptw_customCSRs_csrs_2_sdata;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_3_stall;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        _dcache_io_ptw_customCSRs_csrs_3_set;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire [63:0] _dcache_io_ptw_customCSRs_csrs_3_sdata;	// src/main/scala/rocket/HellaCache.scala:269:43
  wire        broadcast_clock = clock;
  wire        broadcast_reset = reset;
  wire        broadcast_1_clock = clock;
  wire        broadcast_1_reset = reset;
  wire        broadcast_2_clock = clock;
  wire        broadcast_2_reset = reset;
  wire        nexus_clock = clock;
  wire        nexus_reset = reset;
  wire        broadcast_3_clock = clock;
  wire        broadcast_3_reset = reset;
  wire        nexus_1_clock = clock;
  wire        nexus_1_reset = reset;
  wire        broadcast_4_clock = clock;
  wire        broadcast_4_reset = reset;
  wire        widget_clock = clock;
  wire        widget_reset = reset;
  wire        widget_1_clock = clock;
  wire        widget_1_reset = reset;
  wire        fragmenter_clock = clock;
  wire        fragmenter_reset = reset;
  wire        widget_2_clock = clock;
  wire        widget_2_reset = reset;
  wire        buffer_clock = clock;
  wire        buffer_reset = reset;
  wire        buffer_auto_out_a_ready = auto_buffer_out_a_ready;
  wire        buffer_auto_out_b_valid = auto_buffer_out_b_valid;
  wire [2:0]  buffer_auto_out_b_bits_opcode = auto_buffer_out_b_bits_opcode;
  wire [1:0]  buffer_auto_out_b_bits_param = auto_buffer_out_b_bits_param;
  wire [3:0]  buffer_auto_out_b_bits_size = auto_buffer_out_b_bits_size;
  wire [1:0]  buffer_auto_out_b_bits_source = auto_buffer_out_b_bits_source;
  wire [31:0] buffer_auto_out_b_bits_address = auto_buffer_out_b_bits_address;
  wire [7:0]  buffer_auto_out_b_bits_mask = auto_buffer_out_b_bits_mask;
  wire [63:0] buffer_auto_out_b_bits_data = auto_buffer_out_b_bits_data;
  wire        buffer_auto_out_b_bits_corrupt = auto_buffer_out_b_bits_corrupt;
  wire        buffer_auto_out_c_ready = auto_buffer_out_c_ready;
  wire        buffer_auto_out_d_valid = auto_buffer_out_d_valid;
  wire [2:0]  buffer_auto_out_d_bits_opcode = auto_buffer_out_d_bits_opcode;
  wire [1:0]  buffer_auto_out_d_bits_param = auto_buffer_out_d_bits_param;
  wire [3:0]  buffer_auto_out_d_bits_size = auto_buffer_out_d_bits_size;
  wire [1:0]  buffer_auto_out_d_bits_source = auto_buffer_out_d_bits_source;
  wire [1:0]  buffer_auto_out_d_bits_sink = auto_buffer_out_d_bits_sink;
  wire        buffer_auto_out_d_bits_denied = auto_buffer_out_d_bits_denied;
  wire [63:0] buffer_auto_out_d_bits_data = auto_buffer_out_d_bits_data;
  wire        buffer_auto_out_d_bits_corrupt = auto_buffer_out_d_bits_corrupt;
  wire        buffer_auto_out_e_ready = auto_buffer_out_e_ready;
  wire        buffer_1_clock = clock;
  wire        buffer_1_reset = reset;
  wire        hartidIn = auto_hartid_in;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] reset_vectorIn = auto_reset_vector_in;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        nmiIn_rnmi = auto_nmi_in_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] nmiIn_rnmi_interrupt_vector = auto_nmi_in_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] nmiIn_rnmi_exception_vector = auto_nmi_in_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        int_localIn_0 = auto_int_local_in_0_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_0 = auto_int_local_in_1_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_1 = auto_int_local_in_1_1;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        x1_int_localIn_1_0 = auto_int_local_in_2_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_ = 1'h1;	// src/main/scala/tilelink/Bundles.scala:260:61, src/main/scala/tilelink/WidthWidget.scala:206:20
  wire        widget_1__0 = 1'h1;	// src/main/scala/tilelink/Bundles.scala:262:61, src/main/scala/tilelink/WidthWidget.scala:206:20
  wire        widget_1__1 = 1'h1;	// src/main/scala/tilelink/Bundles.scala:259:61, src/main/scala/tilelink/WidthWidget.scala:206:20
  wire [2:0]  widget_1__2 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [2:0]  widget_1__3 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [2:0]  widget_1__4 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [2:0]  widget_1__5 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [2:0]  widget_1__6 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [2:0]  widget_1__7 = 3'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [1:0]  widget_1__8 = 2'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [1:0]  widget_1__9 = 2'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :262:74
  wire [1:0]  widget_1__10 = 2'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [1:0]  widget_1__11 = 2'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :262:74
  wire [3:0]  widget_1__12 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [3:0]  widget_1__13 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [3:0]  widget_1__14 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [3:0]  widget_1__15 = 4'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [3:0]  traceCoreSourceNodeOut_group_0_itype = 4'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [3:0]  traceCoreSourceNodeOut_priv = 4'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [31:0] widget_1__16 = 32'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [31:0] widget_1__17 = 32'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [31:0] widget_1__18 = 32'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [31:0] widget_1__19 = 32'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [31:0] traceCoreSourceNodeOut_group_0_iaddr = 32'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [31:0] traceCoreSourceNodeOut_tval = 32'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [31:0] traceCoreSourceNodeOut_cause = 32'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tilelink/Bundles.scala:259:74
  wire [7:0]  widget_1__20 = 8'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [7:0]  widget_1__21 = 8'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [63:0] widget_1__22 = 64'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [63:0] widget_1__23 = 64'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire [63:0] widget_1__24 = 64'h0;	// src/main/scala/tilelink/Bundles.scala:259:74
  wire [63:0] widget_1__25 = 64'h0;	// src/main/scala/tilelink/Bundles.scala:259:74, :260:74
  wire        nexus_1_x1_bundleOut_x_sourceOpt_enable = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        nexus_1_x1_bundleOut_x_sourceOpt_stall = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        nexus_1_defaultWireOpt_enable = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        nexus_1_defaultWireOpt_stall = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        widget_auto_out_a_valid;
  wire [2:0]  widget_auto_out_a_bits_opcode;
  wire [2:0]  widget_auto_out_a_bits_param;
  wire [3:0]  widget_auto_out_a_bits_size;
  wire        widget_auto_out_a_bits_source;
  wire [31:0] widget_auto_out_a_bits_address;
  wire        widget_auto_out_a_bits_user_amba_prot_bufferable;
  wire        widget_auto_out_a_bits_user_amba_prot_modifiable;
  wire        widget_auto_out_a_bits_user_amba_prot_readalloc;
  wire        widget_auto_out_a_bits_user_amba_prot_writealloc;
  wire        widget_auto_out_a_bits_user_amba_prot_privileged;
  wire        widget_auto_out_a_bits_user_amba_prot_secure;
  wire        widget_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0]  widget_auto_out_a_bits_mask;
  wire [63:0] widget_auto_out_a_bits_data;
  wire        widget_auto_out_a_bits_corrupt;
  wire        widget_auto_out_b_ready;
  wire        widget_auto_out_c_valid;
  wire [2:0]  widget_auto_out_c_bits_opcode;
  wire [2:0]  widget_auto_out_c_bits_param;
  wire [3:0]  widget_auto_out_c_bits_size;
  wire        widget_auto_out_c_bits_source;
  wire [31:0] widget_auto_out_c_bits_address;
  wire        widget_auto_out_c_bits_user_amba_prot_bufferable;
  wire        widget_auto_out_c_bits_user_amba_prot_modifiable;
  wire        widget_auto_out_c_bits_user_amba_prot_readalloc;
  wire        widget_auto_out_c_bits_user_amba_prot_writealloc;
  wire        widget_auto_out_c_bits_user_amba_prot_privileged;
  wire        widget_auto_out_c_bits_user_amba_prot_secure;
  wire        widget_auto_out_c_bits_user_amba_prot_fetch;
  wire [63:0] widget_auto_out_c_bits_data;
  wire        widget_auto_out_c_bits_corrupt;
  wire        widget_auto_out_d_ready;
  wire        widget_auto_out_e_valid;
  wire [1:0]  widget_auto_out_e_bits_sink;
  wire        widget_1_auto_out_a_valid;
  wire [2:0]  widget_1_auto_out_a_bits_opcode;
  wire [2:0]  widget_1_auto_out_a_bits_param;
  wire [3:0]  widget_1_auto_out_a_bits_size;
  wire        widget_1_auto_out_a_bits_source;
  wire [31:0] widget_1_auto_out_a_bits_address;
  wire        widget_1_auto_out_a_bits_user_amba_prot_bufferable;
  wire        widget_1_auto_out_a_bits_user_amba_prot_modifiable;
  wire        widget_1_auto_out_a_bits_user_amba_prot_readalloc;
  wire        widget_1_auto_out_a_bits_user_amba_prot_writealloc;
  wire        widget_1_auto_out_a_bits_user_amba_prot_privileged;
  wire        widget_1_auto_out_a_bits_user_amba_prot_secure;
  wire        widget_1_auto_out_a_bits_user_amba_prot_fetch;
  wire [7:0]  widget_1_auto_out_a_bits_mask;
  wire [63:0] widget_1_auto_out_a_bits_data;
  wire        widget_1_auto_out_a_bits_corrupt;
  wire        widget_1_auto_out_d_ready;
  wire        widget_1__26 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__27 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__28 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__29 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__30 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:61
  wire        widget_1__31 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__32 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__33 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__34 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__35 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__36 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__37 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__38 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__39 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__40 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__41 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__42 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:262:74
  wire        widget_1__43 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:262:74
  wire        widget_1__44 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__45 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__46 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__47 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:259:74
  wire        widget_1__48 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__49 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__50 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__51 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__52 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__53 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__54 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__55 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__56 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__57 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__58 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:74
  wire        widget_1__59 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:260:61
  wire        widget_1__60 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:262:74
  wire        widget_1__61 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:262:74
  wire        widget_1__62 = 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tilelink/Bundles.scala:262:61
  wire        tlOtherMastersNodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeIn_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeIn_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  tlOtherMastersNodeIn_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeIn_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeIn_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        traceCoreSourceNodeOut_group_0_iretire = 1'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:295:16
  wire        traceCoreSourceNodeOut_group_0_ilastsize = 1'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:295:16
  wire        bundleIn_x_sourceOpt_enable = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        bundleIn_x_sourceOpt_stall = 1'h0;	// src/main/scala/tile/BaseTile.scala:294:19, :295:16
  wire        haltNodeOut_0 = 1'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:295:16
  wire        ceaseNodeOut_0 = 1'h0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:295:16
  wire tlMasterXbar_clock;
    wire tlMasterXbar_reset;
    wire tlMasterXbar_auto_in_1_a_ready;
    wire tlMasterXbar_auto_in_1_a_valid;
    wire[2:0] tlMasterXbar_auto_in_1_a_bits_opcode;
    wire[2:0] tlMasterXbar_auto_in_1_a_bits_param;
    wire[3:0] tlMasterXbar_auto_in_1_a_bits_size;
    wire tlMasterXbar_auto_in_1_a_bits_source;
    wire[31:0] tlMasterXbar_auto_in_1_a_bits_address;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_privileged;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_secure;
    wire tlMasterXbar_auto_in_1_a_bits_user_amba_prot_fetch;
    wire[7:0] tlMasterXbar_auto_in_1_a_bits_mask;
    wire[63:0] tlMasterXbar_auto_in_1_a_bits_data;
    wire tlMasterXbar_auto_in_1_a_bits_corrupt;
    wire tlMasterXbar_auto_in_1_d_ready;
    wire tlMasterXbar_auto_in_1_d_valid;
    wire[2:0] tlMasterXbar_auto_in_1_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_in_1_d_bits_param;
    wire[3:0] tlMasterXbar_auto_in_1_d_bits_size;
    wire tlMasterXbar_auto_in_1_d_bits_source;
    wire[1:0] tlMasterXbar_auto_in_1_d_bits_sink;
    wire tlMasterXbar_auto_in_1_d_bits_denied;
    wire[63:0] tlMasterXbar_auto_in_1_d_bits_data;
    wire tlMasterXbar_auto_in_1_d_bits_corrupt;
    wire tlMasterXbar_auto_in_0_a_ready;
    wire tlMasterXbar_auto_in_0_a_valid;
    wire[2:0] tlMasterXbar_auto_in_0_a_bits_opcode;
    wire[2:0] tlMasterXbar_auto_in_0_a_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_a_bits_size;
    wire tlMasterXbar_auto_in_0_a_bits_source;
    wire[31:0] tlMasterXbar_auto_in_0_a_bits_address;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_secure;
    wire tlMasterXbar_auto_in_0_a_bits_user_amba_prot_fetch;
    wire[7:0] tlMasterXbar_auto_in_0_a_bits_mask;
    wire[63:0] tlMasterXbar_auto_in_0_a_bits_data;
    wire tlMasterXbar_auto_in_0_a_bits_corrupt;
    wire tlMasterXbar_auto_in_0_b_ready;
    wire tlMasterXbar_auto_in_0_b_valid;
    wire[2:0] tlMasterXbar_auto_in_0_b_bits_opcode;
    wire[1:0] tlMasterXbar_auto_in_0_b_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_b_bits_size;
    wire tlMasterXbar_auto_in_0_b_bits_source;
    wire[31:0] tlMasterXbar_auto_in_0_b_bits_address;
    wire[7:0] tlMasterXbar_auto_in_0_b_bits_mask;
    wire[63:0] tlMasterXbar_auto_in_0_b_bits_data;
    wire tlMasterXbar_auto_in_0_b_bits_corrupt;
    wire tlMasterXbar_auto_in_0_c_ready;
    wire tlMasterXbar_auto_in_0_c_valid;
    wire[2:0] tlMasterXbar_auto_in_0_c_bits_opcode;
    wire[2:0] tlMasterXbar_auto_in_0_c_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_c_bits_size;
    wire tlMasterXbar_auto_in_0_c_bits_source;
    wire[31:0] tlMasterXbar_auto_in_0_c_bits_address;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_privileged;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_secure;
    wire tlMasterXbar_auto_in_0_c_bits_user_amba_prot_fetch;
    wire[63:0] tlMasterXbar_auto_in_0_c_bits_data;
    wire tlMasterXbar_auto_in_0_c_bits_corrupt;
    wire tlMasterXbar_auto_in_0_d_ready;
    wire tlMasterXbar_auto_in_0_d_valid;
    wire[2:0] tlMasterXbar_auto_in_0_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_in_0_d_bits_param;
    wire[3:0] tlMasterXbar_auto_in_0_d_bits_size;
    wire tlMasterXbar_auto_in_0_d_bits_source;
    wire[1:0] tlMasterXbar_auto_in_0_d_bits_sink;
    wire tlMasterXbar_auto_in_0_d_bits_denied;
    wire[63:0] tlMasterXbar_auto_in_0_d_bits_data;
    wire tlMasterXbar_auto_in_0_d_bits_corrupt;
    wire tlMasterXbar_auto_in_0_e_ready;
    wire tlMasterXbar_auto_in_0_e_valid;
    wire[1:0] tlMasterXbar_auto_in_0_e_bits_sink;
    wire tlMasterXbar_auto_out_a_ready;
    wire tlMasterXbar_auto_out_a_valid;
    wire[2:0] tlMasterXbar_auto_out_a_bits_opcode;
    wire[2:0] tlMasterXbar_auto_out_a_bits_param;
    wire[3:0] tlMasterXbar_auto_out_a_bits_size;
    wire[1:0] tlMasterXbar_auto_out_a_bits_source;
    wire[31:0] tlMasterXbar_auto_out_a_bits_address;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_secure;
    wire tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch;
    wire[7:0] tlMasterXbar_auto_out_a_bits_mask;
    wire[63:0] tlMasterXbar_auto_out_a_bits_data;
    wire tlMasterXbar_auto_out_a_bits_corrupt;
    wire tlMasterXbar_auto_out_b_ready;
    wire tlMasterXbar_auto_out_b_valid;
    wire[2:0] tlMasterXbar_auto_out_b_bits_opcode;
    wire[1:0] tlMasterXbar_auto_out_b_bits_param;
    wire[3:0] tlMasterXbar_auto_out_b_bits_size;
    wire[1:0] tlMasterXbar_auto_out_b_bits_source;
    wire[31:0] tlMasterXbar_auto_out_b_bits_address;
    wire[7:0] tlMasterXbar_auto_out_b_bits_mask;
    wire[63:0] tlMasterXbar_auto_out_b_bits_data;
    wire tlMasterXbar_auto_out_b_bits_corrupt;
    wire tlMasterXbar_auto_out_c_ready;
    wire tlMasterXbar_auto_out_c_valid;
    wire[2:0] tlMasterXbar_auto_out_c_bits_opcode;
    wire[2:0] tlMasterXbar_auto_out_c_bits_param;
    wire[3:0] tlMasterXbar_auto_out_c_bits_size;
    wire[1:0] tlMasterXbar_auto_out_c_bits_source;
    wire[31:0] tlMasterXbar_auto_out_c_bits_address;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_privileged;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_secure;
    wire tlMasterXbar_auto_out_c_bits_user_amba_prot_fetch;
    wire[63:0] tlMasterXbar_auto_out_c_bits_data;
    wire tlMasterXbar_auto_out_c_bits_corrupt;
    wire tlMasterXbar_auto_out_d_ready;
    wire tlMasterXbar_auto_out_d_valid;
    wire[2:0] tlMasterXbar_auto_out_d_bits_opcode;
    wire[1:0] tlMasterXbar_auto_out_d_bits_param;
    wire[3:0] tlMasterXbar_auto_out_d_bits_size;
    wire[1:0] tlMasterXbar_auto_out_d_bits_source;
    wire[1:0] tlMasterXbar_auto_out_d_bits_sink;
    wire tlMasterXbar_auto_out_d_bits_denied;
    wire[63:0] tlMasterXbar_auto_out_d_bits_data;
    wire tlMasterXbar_auto_out_d_bits_corrupt;
    wire tlMasterXbar_auto_out_e_ready;
    wire tlMasterXbar_auto_out_e_valid;
    wire[1:0] tlMasterXbar_auto_out_e_bits_sink;

    wire[1:0] tlMasterXbar_in_1_a_bits_source ; 
    wire[1:0] tlMasterXbar_in_0_c_bits_source ; 
    wire[1:0] tlMasterXbar_in_0_a_bits_source ; 
    wire tlMasterXbar_nodeIn_a_valid = tlMasterXbar_auto_in_0_a_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_a_bits_opcode = tlMasterXbar_auto_in_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_a_bits_param = tlMasterXbar_auto_in_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_a_bits_size = tlMasterXbar_auto_in_0_a_bits_size ; 
    wire tlMasterXbar_nodeIn_a_bits_source = tlMasterXbar_auto_in_0_a_bits_source ; 
    wire[31:0] tlMasterXbar_nodeIn_a_bits_address = tlMasterXbar_auto_in_0_a_bits_address ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_bufferable = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_modifiable = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_privileged = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_secure = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_nodeIn_a_bits_user_amba_prot_fetch = tlMasterXbar_auto_in_0_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar_nodeIn_a_bits_mask = tlMasterXbar_auto_in_0_a_bits_mask ; 
    wire[63:0] tlMasterXbar_nodeIn_a_bits_data = tlMasterXbar_auto_in_0_a_bits_data ; 
    wire tlMasterXbar_nodeIn_a_bits_corrupt = tlMasterXbar_auto_in_0_a_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_b_ready = tlMasterXbar_auto_in_0_b_ready ; 
    wire tlMasterXbar_nodeIn_c_valid = tlMasterXbar_auto_in_0_c_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_c_bits_opcode = tlMasterXbar_auto_in_0_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_c_bits_param = tlMasterXbar_auto_in_0_c_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_c_bits_size = tlMasterXbar_auto_in_0_c_bits_size ; 
    wire tlMasterXbar_nodeIn_c_bits_source = tlMasterXbar_auto_in_0_c_bits_source ; 
    wire[31:0] tlMasterXbar_nodeIn_c_bits_address = tlMasterXbar_auto_in_0_c_bits_address ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_bufferable = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_modifiable = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_privileged = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_secure = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_nodeIn_c_bits_user_amba_prot_fetch = tlMasterXbar_auto_in_0_c_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_nodeIn_c_bits_data = tlMasterXbar_auto_in_0_c_bits_data ; 
    wire tlMasterXbar_nodeIn_c_bits_corrupt = tlMasterXbar_auto_in_0_c_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_d_ready = tlMasterXbar_auto_in_0_d_ready ; 
    wire tlMasterXbar_nodeIn_e_valid = tlMasterXbar_auto_in_0_e_valid ; 
    wire[1:0] tlMasterXbar_nodeIn_e_bits_sink = tlMasterXbar_auto_in_0_e_bits_sink ; 
    wire tlMasterXbar_nodeIn_1_a_valid = tlMasterXbar_auto_in_1_a_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_1_a_bits_opcode = tlMasterXbar_auto_in_1_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeIn_1_a_bits_param = tlMasterXbar_auto_in_1_a_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_1_a_bits_size = tlMasterXbar_auto_in_1_a_bits_size ; 
    wire tlMasterXbar_nodeIn_1_a_bits_source = tlMasterXbar_auto_in_1_a_bits_source ; 
    wire[31:0] tlMasterXbar_nodeIn_1_a_bits_address = tlMasterXbar_auto_in_1_a_bits_address ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_bufferable = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_modifiable = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_privileged = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_secure = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_fetch = tlMasterXbar_auto_in_1_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar_nodeIn_1_a_bits_mask = tlMasterXbar_auto_in_1_a_bits_mask ; 
    wire[63:0] tlMasterXbar_nodeIn_1_a_bits_data = tlMasterXbar_auto_in_1_a_bits_data ; 
    wire tlMasterXbar_nodeIn_1_a_bits_corrupt = tlMasterXbar_auto_in_1_a_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_1_d_ready = tlMasterXbar_auto_in_1_d_ready ; 
    wire tlMasterXbar_nodeOut_a_ready = tlMasterXbar_auto_out_a_ready ; 
    wire tlMasterXbar_nodeOut_b_valid = tlMasterXbar_auto_out_b_valid ; 
    wire[2:0] tlMasterXbar_nodeOut_b_bits_opcode = tlMasterXbar_auto_out_b_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeOut_b_bits_param = tlMasterXbar_auto_out_b_bits_param ; 
    wire[3:0] tlMasterXbar_nodeOut_b_bits_size = tlMasterXbar_auto_out_b_bits_size ; 
    wire[1:0] tlMasterXbar_nodeOut_b_bits_source = tlMasterXbar_auto_out_b_bits_source ; 
    wire[31:0] tlMasterXbar_nodeOut_b_bits_address = tlMasterXbar_auto_out_b_bits_address ; 
    wire[7:0] tlMasterXbar_nodeOut_b_bits_mask = tlMasterXbar_auto_out_b_bits_mask ; 
    wire[63:0] tlMasterXbar_nodeOut_b_bits_data = tlMasterXbar_auto_out_b_bits_data ; 
    wire tlMasterXbar_nodeOut_b_bits_corrupt = tlMasterXbar_auto_out_b_bits_corrupt ; 
    wire tlMasterXbar_nodeOut_c_ready = tlMasterXbar_auto_out_c_ready ; 
    wire tlMasterXbar_nodeOut_d_valid = tlMasterXbar_auto_out_d_valid ; 
    wire[2:0] tlMasterXbar_nodeOut_d_bits_opcode = tlMasterXbar_auto_out_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeOut_d_bits_param = tlMasterXbar_auto_out_d_bits_param ; 
    wire[3:0] tlMasterXbar_nodeOut_d_bits_size = tlMasterXbar_auto_out_d_bits_size ; 
    wire[1:0] tlMasterXbar_nodeOut_d_bits_source = tlMasterXbar_auto_out_d_bits_source ; 
    wire[1:0] tlMasterXbar_nodeOut_d_bits_sink = tlMasterXbar_auto_out_d_bits_sink ; 
    wire tlMasterXbar_nodeOut_d_bits_denied = tlMasterXbar_auto_out_d_bits_denied ; 
    wire[63:0] tlMasterXbar_nodeOut_d_bits_data = tlMasterXbar_auto_out_d_bits_data ; 
    wire tlMasterXbar_nodeOut_d_bits_corrupt = tlMasterXbar_auto_out_d_bits_corrupt ; 
    wire tlMasterXbar_nodeOut_e_ready = tlMasterXbar_auto_out_e_ready ; 
    wire[8:0] tlMasterXbar_beatsBO_0 =9'h0; 
    wire[8:0] tlMasterXbar_beatsCI_1 =9'h0; 
    wire tlMasterXbar_in_1_b_ready =1'h1; 
    wire tlMasterXbar__GEN =1'h1; 
    wire tlMasterXbar__GEN_0 =1'h1; 
    wire tlMasterXbar_requestAIO_0_0 =1'h1; 
    wire tlMasterXbar_requestAIO_1_0 =1'h1; 
    wire tlMasterXbar_requestCIO_0_0 =1'h1; 
    wire tlMasterXbar_requestCIO_1_0 =1'h1; 
    wire[2:0] tlMasterXbar_in_1_b_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_in_1_c_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_in_1_c_bits_param =3'h0; 
    wire[2:0] tlMasterXbar__GEN_1 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_2 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_3 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_4 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_5 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_6 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_7 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_8 =3'h0; 
    wire[2:0] tlMasterXbar__GEN_9 =3'h0; 
    wire[1:0] tlMasterXbar_in_1_b_bits_param =2'h0; 
    wire[1:0] tlMasterXbar_in_1_b_bits_source =2'h0; 
    wire[1:0] tlMasterXbar_in_1_c_bits_source =2'h0; 
    wire[1:0] tlMasterXbar_in_1_e_bits_sink =2'h0; 
    wire[1:0] tlMasterXbar__GEN_10 =2'h0; 
    wire[1:0] tlMasterXbar__GEN_11 =2'h0; 
    wire[1:0] tlMasterXbar__GEN_12 =2'h0; 
    wire[1:0] tlMasterXbar__GEN_13 =2'h0; 
    wire[1:0] tlMasterXbar__GEN_14 =2'h0; 
    wire[1:0] tlMasterXbar__GEN_15 =2'h0; 
    wire[3:0] tlMasterXbar_in_1_b_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_in_1_c_bits_size =4'h0; 
    wire[3:0] tlMasterXbar__GEN_16 =4'h0; 
    wire[3:0] tlMasterXbar__GEN_17 =4'h0; 
    wire[3:0] tlMasterXbar__GEN_18 =4'h0; 
    wire[3:0] tlMasterXbar__GEN_19 =4'h0; 
    wire[3:0] tlMasterXbar__GEN_20 =4'h0; 
    wire[3:0] tlMasterXbar__GEN_21 =4'h0; 
    wire[31:0] tlMasterXbar_in_1_b_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_in_1_c_bits_address =32'h0; 
    wire[31:0] tlMasterXbar__GEN_22 =32'h0; 
    wire[31:0] tlMasterXbar__GEN_23 =32'h0; 
    wire[31:0] tlMasterXbar__GEN_24 =32'h0; 
    wire[31:0] tlMasterXbar__GEN_25 =32'h0; 
    wire[31:0] tlMasterXbar__GEN_26 =32'h0; 
    wire[31:0] tlMasterXbar__GEN_27 =32'h0; 
    wire[7:0] tlMasterXbar_in_1_b_bits_mask =8'h0; 
    wire[7:0] tlMasterXbar__GEN_28 =8'h0; 
    wire[7:0] tlMasterXbar__GEN_29 =8'h0; 
    wire[7:0] tlMasterXbar__GEN_30 =8'h0; 
    wire[63:0] tlMasterXbar_in_1_b_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_in_1_c_bits_data =64'h0; 
    wire[63:0] tlMasterXbar__GEN_31 =64'h0; 
    wire[63:0] tlMasterXbar__GEN_32 =64'h0; 
    wire[63:0] tlMasterXbar__GEN_33 =64'h0; 
    wire[63:0] tlMasterXbar__GEN_34 =64'h0; 
    wire[63:0] tlMasterXbar__GEN_35 =64'h0; 
    wire[63:0] tlMasterXbar__GEN_36 =64'h0; 
    wire tlMasterXbar_nodeIn_1_d_bits_source =1'h0; 
    wire tlMasterXbar_in_0_a_ready ; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_0_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_0_c_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_1_a_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_1_b_valid =1'h0; 
    wire tlMasterXbar_in_1_b_bits_corrupt =1'h0; 
    wire tlMasterXbar_in_1_c_valid =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_in_1_c_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_in_1_c_bits_corrupt =1'h0; 
    wire tlMasterXbar_in_1_e_valid =1'h0; 
    wire tlMasterXbar__GEN_37 =1'h0; 
    wire tlMasterXbar__GEN_38 =1'h0; 
    wire tlMasterXbar__GEN_39 =1'h0; 
    wire tlMasterXbar__GEN_40 =1'h0; 
    wire tlMasterXbar__GEN_41 =1'h0; 
    wire tlMasterXbar__GEN_42 =1'h0; 
    wire tlMasterXbar__GEN_43 =1'h0; 
    wire tlMasterXbar__GEN_44 =1'h0; 
    wire tlMasterXbar__GEN_45 =1'h0; 
    wire tlMasterXbar__GEN_46 =1'h0; 
    wire tlMasterXbar__GEN_47 =1'h0; 
    wire tlMasterXbar__GEN_48 =1'h0; 
    wire tlMasterXbar__GEN_49 =1'h0; 
    wire tlMasterXbar__GEN_50 =1'h0; 
    wire tlMasterXbar__GEN_51 =1'h0; 
    wire tlMasterXbar__GEN_52 =1'h0; 
    wire tlMasterXbar__GEN_53 =1'h0; 
    wire tlMasterXbar__GEN_54 =1'h0; 
    wire tlMasterXbar__GEN_55 =1'h0; 
    wire tlMasterXbar__GEN_56 =1'h0; 
    wire tlMasterXbar__GEN_57 =1'h0; 
    wire tlMasterXbar__GEN_58 =1'h0; 
    wire tlMasterXbar__GEN_59 =1'h0; 
    wire tlMasterXbar__GEN_60 =1'h0; 
    wire tlMasterXbar__GEN_61 =1'h0; 
    wire tlMasterXbar__GEN_62 =1'h0; 
    wire tlMasterXbar__GEN_63 =1'h0; 
    wire tlMasterXbar__GEN_64 =1'h0; 
    wire tlMasterXbar__GEN_65 =1'h0; 
    wire tlMasterXbar__GEN_66 =1'h0; 
    wire tlMasterXbar__GEN_67 =1'h0; 
    wire tlMasterXbar__GEN_68 =1'h0; 
    wire tlMasterXbar__GEN_69 =1'h0; 
    wire tlMasterXbar__GEN_70 =1'h0; 
    wire tlMasterXbar__GEN_71 =1'h0; 
    wire tlMasterXbar__GEN_72 =1'h0; 
    wire tlMasterXbar__GEN_73 =1'h0; 
    wire tlMasterXbar__GEN_74 =1'h0; 
    wire tlMasterXbar__GEN_75 =1'h0; 
    wire tlMasterXbar__GEN_76 =1'h0; 
    wire tlMasterXbar__GEN_77 =1'h0; 
    wire tlMasterXbar__GEN_78 =1'h0; 
    wire tlMasterXbar__GEN_79 =1'h0; 
    wire tlMasterXbar__GEN_80 =1'h0; 
    wire tlMasterXbar__GEN_81 =1'h0; 
    wire tlMasterXbar__GEN_82 =1'h0; 
    wire tlMasterXbar__GEN_83 =1'h0; 
    wire tlMasterXbar__GEN_84 =1'h0; 
    wire tlMasterXbar__GEN_85 =1'h0; 
    wire tlMasterXbar__GEN_86 =1'h0; 
    wire tlMasterXbar__GEN_87 =1'h0; 
    wire tlMasterXbar__GEN_88 =1'h0; 
    wire tlMasterXbar_portsBIO_filtered_1_ready =1'h0; 
    wire tlMasterXbar_portsCOI_filtered_1_0_ready =1'h0; 
    wire tlMasterXbar_portsEOI_filtered_1_0_ready =1'h0; 
    wire tlMasterXbar__state_WIRE_0 =1'h0; 
    wire tlMasterXbar__state_WIRE_1 =1'h0; 
    wire tlMasterXbar_in_0_a_valid = tlMasterXbar_nodeIn_a_valid ; 
    wire[2:0] tlMasterXbar_in_0_a_bits_opcode = tlMasterXbar_nodeIn_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_in_0_a_bits_param = tlMasterXbar_nodeIn_a_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_a_bits_size = tlMasterXbar_nodeIn_a_bits_size ; 
    wire[31:0] tlMasterXbar_in_0_a_bits_address = tlMasterXbar_nodeIn_a_bits_address ; 
    wire[7:0] tlMasterXbar_in_0_a_bits_mask = tlMasterXbar_nodeIn_a_bits_mask ; 
    wire[63:0] tlMasterXbar_in_0_a_bits_data = tlMasterXbar_nodeIn_a_bits_data ; 
    wire tlMasterXbar_in_0_a_bits_corrupt = tlMasterXbar_nodeIn_a_bits_corrupt ; 
    wire tlMasterXbar_in_0_b_ready = tlMasterXbar_nodeIn_b_ready ; 
    wire tlMasterXbar_in_0_b_valid ; 
    wire[2:0] tlMasterXbar_in_0_b_bits_opcode ; 
    wire[1:0] tlMasterXbar_in_0_b_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_b_bits_size ; 
    wire[31:0] tlMasterXbar_in_0_b_bits_address ; 
    wire[7:0] tlMasterXbar_in_0_b_bits_mask ; 
    wire[63:0] tlMasterXbar_in_0_b_bits_data ; 
    wire tlMasterXbar_in_0_b_bits_corrupt ; 
    wire tlMasterXbar_in_0_c_ready ; 
    wire tlMasterXbar_in_0_c_valid = tlMasterXbar_nodeIn_c_valid ; 
    wire[2:0] tlMasterXbar_in_0_c_bits_opcode = tlMasterXbar_nodeIn_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_in_0_c_bits_param = tlMasterXbar_nodeIn_c_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_c_bits_size = tlMasterXbar_nodeIn_c_bits_size ; 
    wire[31:0] tlMasterXbar_in_0_c_bits_address = tlMasterXbar_nodeIn_c_bits_address ; 
    wire[63:0] tlMasterXbar_in_0_c_bits_data = tlMasterXbar_nodeIn_c_bits_data ; 
    wire tlMasterXbar_in_0_c_bits_corrupt = tlMasterXbar_nodeIn_c_bits_corrupt ; 
    wire tlMasterXbar_in_0_d_ready = tlMasterXbar_nodeIn_d_ready ; 
    wire tlMasterXbar_in_0_d_valid ; 
    wire[2:0] tlMasterXbar_in_0_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_in_0_d_bits_param ; 
    wire[3:0] tlMasterXbar_in_0_d_bits_size ; 
    wire[1:0] tlMasterXbar_in_0_d_bits_sink ; 
    wire tlMasterXbar_in_0_d_bits_denied ; 
    wire[63:0] tlMasterXbar_in_0_d_bits_data ; 
    wire tlMasterXbar_in_0_d_bits_corrupt ; 
    wire tlMasterXbar_in_0_e_ready ; 
    wire tlMasterXbar_in_0_e_valid = tlMasterXbar_nodeIn_e_valid ; 
    wire[1:0] tlMasterXbar_in_0_e_bits_sink = tlMasterXbar_nodeIn_e_bits_sink ; 
    wire tlMasterXbar_in_1_a_ready ; 
    wire tlMasterXbar_in_1_a_valid = tlMasterXbar_nodeIn_1_a_valid ; 
    wire[2:0] tlMasterXbar_in_1_a_bits_opcode = tlMasterXbar_nodeIn_1_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_in_1_a_bits_param = tlMasterXbar_nodeIn_1_a_bits_param ; 
    wire[3:0] tlMasterXbar_in_1_a_bits_size = tlMasterXbar_nodeIn_1_a_bits_size ; 
    wire[31:0] tlMasterXbar_in_1_a_bits_address = tlMasterXbar_nodeIn_1_a_bits_address ; 
    wire[7:0] tlMasterXbar_in_1_a_bits_mask = tlMasterXbar_nodeIn_1_a_bits_mask ; 
    wire[63:0] tlMasterXbar_in_1_a_bits_data = tlMasterXbar_nodeIn_1_a_bits_data ; 
    wire tlMasterXbar_in_1_a_bits_corrupt = tlMasterXbar_nodeIn_1_a_bits_corrupt ; 
    wire tlMasterXbar_in_1_d_ready = tlMasterXbar_nodeIn_1_d_ready ; 
    wire tlMasterXbar_in_1_d_valid ; 
    wire[2:0] tlMasterXbar_in_1_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_in_1_d_bits_param ; 
    wire[3:0] tlMasterXbar_in_1_d_bits_size ; 
    wire[1:0] tlMasterXbar_in_1_d_bits_sink ; 
    wire tlMasterXbar_in_1_d_bits_denied ; 
    wire[63:0] tlMasterXbar_in_1_d_bits_data ; 
    wire tlMasterXbar_in_1_d_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_a_ready ; 
    wire tlMasterXbar_nodeIn_b_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_b_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeIn_b_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_b_bits_size ; 
    wire tlMasterXbar_nodeIn_b_bits_source ; 
    wire[31:0] tlMasterXbar_nodeIn_b_bits_address ; 
    wire[7:0] tlMasterXbar_nodeIn_b_bits_mask ; 
    wire[63:0] tlMasterXbar_nodeIn_b_bits_data ; 
    wire tlMasterXbar_nodeIn_b_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_c_ready ; 
    wire tlMasterXbar_nodeIn_d_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeIn_d_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_d_bits_size ; 
    wire tlMasterXbar_nodeIn_d_bits_source ; 
    wire[1:0] tlMasterXbar_nodeIn_d_bits_sink ; 
    wire tlMasterXbar_nodeIn_d_bits_denied ; 
    wire[63:0] tlMasterXbar_nodeIn_d_bits_data ; 
    wire tlMasterXbar_nodeIn_d_bits_corrupt ; 
    wire tlMasterXbar_nodeIn_e_ready ;  
    wire tlMasterXbar_monitor_clock;
    wire tlMasterXbar_monitor_reset;
    wire tlMasterXbar_monitor_io_in_a_ready;
    wire tlMasterXbar_monitor_io_in_a_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_a_bits_opcode;
    wire[2:0] tlMasterXbar_monitor_io_in_a_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_a_bits_size;
    wire tlMasterXbar_monitor_io_in_a_bits_source;
    wire[31:0] tlMasterXbar_monitor_io_in_a_bits_address;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_privileged;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_secure;
    wire tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_fetch;
    wire[7:0] tlMasterXbar_monitor_io_in_a_bits_mask;
    wire[63:0] tlMasterXbar_monitor_io_in_a_bits_data;
    wire tlMasterXbar_monitor_io_in_a_bits_corrupt;
    wire tlMasterXbar_monitor_io_in_b_ready;
    wire tlMasterXbar_monitor_io_in_b_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_b_bits_opcode;
    wire[1:0] tlMasterXbar_monitor_io_in_b_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_b_bits_size;
    wire tlMasterXbar_monitor_io_in_b_bits_source;
    wire[31:0] tlMasterXbar_monitor_io_in_b_bits_address;
    wire[7:0] tlMasterXbar_monitor_io_in_b_bits_mask;
    wire[63:0] tlMasterXbar_monitor_io_in_b_bits_data;
    wire tlMasterXbar_monitor_io_in_b_bits_corrupt;
    wire tlMasterXbar_monitor_io_in_c_ready;
    wire tlMasterXbar_monitor_io_in_c_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_c_bits_opcode;
    wire[2:0] tlMasterXbar_monitor_io_in_c_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_c_bits_size;
    wire tlMasterXbar_monitor_io_in_c_bits_source;
    wire[31:0] tlMasterXbar_monitor_io_in_c_bits_address;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_privileged;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_secure;
    wire tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_fetch;
    wire[63:0] tlMasterXbar_monitor_io_in_c_bits_data;
    wire tlMasterXbar_monitor_io_in_c_bits_corrupt;
    wire tlMasterXbar_monitor_io_in_d_ready;
    wire tlMasterXbar_monitor_io_in_d_valid;
    wire[2:0] tlMasterXbar_monitor_io_in_d_bits_opcode;
    wire[1:0] tlMasterXbar_monitor_io_in_d_bits_param;
    wire[3:0] tlMasterXbar_monitor_io_in_d_bits_size;
    wire tlMasterXbar_monitor_io_in_d_bits_source;
    wire[1:0] tlMasterXbar_monitor_io_in_d_bits_sink;
    wire tlMasterXbar_monitor_io_in_d_bits_denied;
    wire[63:0] tlMasterXbar_monitor_io_in_d_bits_data;
    wire tlMasterXbar_monitor_io_in_d_bits_corrupt;
    wire tlMasterXbar_monitor_io_in_e_ready;
    wire tlMasterXbar_monitor_io_in_e_valid;
    wire[1:0] tlMasterXbar_monitor_io_in_e_bits_sink;

    wire[31:0] tlMasterXbar_monitor__plusarg_reader_1_out ; 
    wire[31:0] tlMasterXbar_monitor__plusarg_reader_out ; 
    wire[8:0] tlMasterXbar_monitor_b_first_beats1 =9'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_6 =3'h5; 
    wire[2:0] tlMasterXbar_monitor_responseMap_6 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_responseMap_7 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_7 =3'h4; 
    wire tlMasterXbar_monitor__GEN = tlMasterXbar_monitor_io_in_a_bits_opcode <=3'h7==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_0 = tlMasterXbar_monitor_io_in_a_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_1 =& tlMasterXbar_monitor_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor_source_ok = tlMasterXbar_monitor__source_ok_WIRE_0 | tlMasterXbar_monitor__source_ok_WIRE_1 ; 
    wire[26:0] tlMasterXbar_monitor__GEN_0 =27'hFFF<< tlMasterXbar_monitor_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_is_aligned_mask =~( tlMasterXbar_monitor__GEN_0 [11:0]); 
    wire tlMasterXbar_monitor_is_aligned =( tlMasterXbar_monitor_io_in_a_bits_address &{20'h0, tlMasterXbar_monitor_is_aligned_mask })==32'h0; 
    wire[1:0] tlMasterXbar_monitor_mask_sizeOH_shiftAmount = tlMasterXbar_monitor_io_in_a_bits_size [1:0]; 
    wire[3:0] tlMasterXbar_monitor__GEN_1 =4'h1<< tlMasterXbar_monitor_mask_sizeOH_shiftAmount ; 
    wire[2:0] tlMasterXbar_monitor_mask_sizeOH = tlMasterXbar_monitor__GEN_1 [2:0]|3'h1; 
    wire tlMasterXbar_monitor__GEN_2 = tlMasterXbar_monitor_io_in_a_bits_size >=4'h3; 
    wire tlMasterXbar_monitor_mask_size = tlMasterXbar_monitor_mask_sizeOH [2]; 
    wire tlMasterXbar_monitor_mask_bit = tlMasterXbar_monitor_io_in_a_bits_address [2]; 
    wire tlMasterXbar_monitor_mask_nbit = tlMasterXbar_monitor_mask_bit ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq = tlMasterXbar_monitor_mask_nbit &1'h1; 
    wire tlMasterXbar_monitor_mask_acc = tlMasterXbar_monitor__GEN_2 | tlMasterXbar_monitor_mask_size & tlMasterXbar_monitor_mask_eq ; 
    wire tlMasterXbar_monitor_mask_eq_1 = tlMasterXbar_monitor_mask_bit &1'h1; 
    wire tlMasterXbar_monitor_mask_acc_1 = tlMasterXbar_monitor__GEN_2 | tlMasterXbar_monitor_mask_size & tlMasterXbar_monitor_mask_eq_1 ; 
    wire tlMasterXbar_monitor_mask_size_1 = tlMasterXbar_monitor_mask_sizeOH [1]; 
    wire tlMasterXbar_monitor_mask_bit_1 = tlMasterXbar_monitor_io_in_a_bits_address [1]; 
    wire tlMasterXbar_monitor_mask_nbit_1 = tlMasterXbar_monitor_mask_bit_1 ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq_2 = tlMasterXbar_monitor_mask_eq & tlMasterXbar_monitor_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_2 = tlMasterXbar_monitor_mask_acc | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_2 ; 
    wire tlMasterXbar_monitor_mask_eq_3 = tlMasterXbar_monitor_mask_eq & tlMasterXbar_monitor_mask_bit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_3 = tlMasterXbar_monitor_mask_acc | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_3 ; 
    wire tlMasterXbar_monitor_mask_eq_4 = tlMasterXbar_monitor_mask_eq_1 & tlMasterXbar_monitor_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_4 = tlMasterXbar_monitor_mask_acc_1 | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_4 ; 
    wire tlMasterXbar_monitor_mask_eq_5 = tlMasterXbar_monitor_mask_eq_1 & tlMasterXbar_monitor_mask_bit_1 ; 
    wire tlMasterXbar_monitor_mask_acc_5 = tlMasterXbar_monitor_mask_acc_1 | tlMasterXbar_monitor_mask_size_1 & tlMasterXbar_monitor_mask_eq_5 ; 
    wire tlMasterXbar_monitor_mask_size_2 = tlMasterXbar_monitor_mask_sizeOH [0]; 
    wire tlMasterXbar_monitor_mask_bit_2 = tlMasterXbar_monitor_io_in_a_bits_address [0]; 
    wire tlMasterXbar_monitor_mask_nbit_2 = tlMasterXbar_monitor_mask_bit_2 ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq_6 = tlMasterXbar_monitor_mask_eq_2 & tlMasterXbar_monitor_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_6 = tlMasterXbar_monitor_mask_acc_2 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_6 ; 
    wire tlMasterXbar_monitor_mask_eq_7 = tlMasterXbar_monitor_mask_eq_2 & tlMasterXbar_monitor_mask_bit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_7 = tlMasterXbar_monitor_mask_acc_2 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_7 ; 
    wire tlMasterXbar_monitor_mask_eq_8 = tlMasterXbar_monitor_mask_eq_3 & tlMasterXbar_monitor_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_8 = tlMasterXbar_monitor_mask_acc_3 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_8 ; 
    wire tlMasterXbar_monitor_mask_eq_9 = tlMasterXbar_monitor_mask_eq_3 & tlMasterXbar_monitor_mask_bit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_9 = tlMasterXbar_monitor_mask_acc_3 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_9 ; 
    wire tlMasterXbar_monitor_mask_eq_10 = tlMasterXbar_monitor_mask_eq_4 & tlMasterXbar_monitor_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_10 = tlMasterXbar_monitor_mask_acc_4 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_10 ; 
    wire tlMasterXbar_monitor_mask_eq_11 = tlMasterXbar_monitor_mask_eq_4 & tlMasterXbar_monitor_mask_bit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_11 = tlMasterXbar_monitor_mask_acc_4 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_11 ; 
    wire tlMasterXbar_monitor_mask_eq_12 = tlMasterXbar_monitor_mask_eq_5 & tlMasterXbar_monitor_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_12 = tlMasterXbar_monitor_mask_acc_5 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_12 ; 
    wire tlMasterXbar_monitor_mask_eq_13 = tlMasterXbar_monitor_mask_eq_5 & tlMasterXbar_monitor_mask_bit_2 ; 
    wire tlMasterXbar_monitor_mask_acc_13 = tlMasterXbar_monitor_mask_acc_5 | tlMasterXbar_monitor_mask_size_2 & tlMasterXbar_monitor_mask_eq_13 ; 
    wire[1:0] tlMasterXbar_monitor_mask_lo_lo ={ tlMasterXbar_monitor_mask_acc_7 , tlMasterXbar_monitor_mask_acc_6 }; 
    wire[1:0] tlMasterXbar_monitor_mask_lo_hi ={ tlMasterXbar_monitor_mask_acc_9 , tlMasterXbar_monitor_mask_acc_8 }; 
    wire[3:0] tlMasterXbar_monitor_mask_lo ={ tlMasterXbar_monitor_mask_lo_hi , tlMasterXbar_monitor_mask_lo_lo }; 
    wire[1:0] tlMasterXbar_monitor_mask_hi_lo ={ tlMasterXbar_monitor_mask_acc_11 , tlMasterXbar_monitor_mask_acc_10 }; 
    wire[1:0] tlMasterXbar_monitor_mask_hi_hi ={ tlMasterXbar_monitor_mask_acc_13 , tlMasterXbar_monitor_mask_acc_12 }; 
    wire[3:0] tlMasterXbar_monitor_mask_hi ={ tlMasterXbar_monitor_mask_hi_hi , tlMasterXbar_monitor_mask_hi_lo }; 
    wire[7:0] tlMasterXbar_monitor_mask ={ tlMasterXbar_monitor_mask_hi , tlMasterXbar_monitor_mask_lo }; 
    wire tlMasterXbar_monitor__GEN_3 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor__GEN_4 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_5 = tlMasterXbar_monitor_io_in_a_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_6 =& tlMasterXbar_monitor_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor__GEN_7 = tlMasterXbar_monitor__GEN_5  ? 4'h6== tlMasterXbar_monitor_io_in_a_bits_size :1'h0; 
    wire tlMasterXbar_monitor__GEN_8 =( tlMasterXbar_monitor__GEN_7 &((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_9 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_10 = tlMasterXbar_monitor_io_in_a_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_11 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_12 = tlMasterXbar_monitor_io_in_a_bits_param <=3'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_13 =~ tlMasterXbar_monitor_io_in_a_bits_mask ==8'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_14 = tlMasterXbar_monitor_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_15 = tlMasterXbar_monitor_io_in_a_valid &(& tlMasterXbar_monitor_io_in_a_bits_opcode ); 
    wire tlMasterXbar_monitor__GEN_16 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_17 = tlMasterXbar_monitor_io_in_a_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_18 =& tlMasterXbar_monitor_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor__GEN_19 = tlMasterXbar_monitor__GEN_17  ? 4'h6== tlMasterXbar_monitor_io_in_a_bits_size :1'h0; 
    wire tlMasterXbar_monitor__GEN_20 =( tlMasterXbar_monitor__GEN_19 &((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_21 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_22 = tlMasterXbar_monitor_io_in_a_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_23 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_24 = tlMasterXbar_monitor_io_in_a_bits_param <=3'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_25 =(| tlMasterXbar_monitor_io_in_a_bits_param )==1'h0; 
    wire tlMasterXbar_monitor__GEN_26 =~ tlMasterXbar_monitor_io_in_a_bits_mask ==8'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_27 = tlMasterXbar_monitor_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_28 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor__GEN_29 =(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)==1'h0; 
    wire tlMasterXbar_monitor__GEN_30 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_31 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_32 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_33 = tlMasterXbar_monitor_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_34 = tlMasterXbar_monitor_io_in_a_bits_mask == tlMasterXbar_monitor_mask ==1'h0; 
    wire tlMasterXbar_monitor__GEN_35 = tlMasterXbar_monitor_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_36 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor__GEN_37 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h8|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_38 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_39 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_40 = tlMasterXbar_monitor_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_41 = tlMasterXbar_monitor_io_in_a_bits_mask == tlMasterXbar_monitor_mask ==1'h0; 
    wire tlMasterXbar_monitor__GEN_42 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor__GEN_43 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|(4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h8|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_44 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_45 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_46 = tlMasterXbar_monitor_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_47 =( tlMasterXbar_monitor_io_in_a_bits_mask &~ tlMasterXbar_monitor_mask )==8'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_48 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor__GEN_49 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h3|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_50 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_51 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_52 = tlMasterXbar_monitor_io_in_a_bits_param <=3'h4==1'h0; 
    wire tlMasterXbar_monitor__GEN_53 = tlMasterXbar_monitor_io_in_a_bits_mask == tlMasterXbar_monitor_mask ==1'h0; 
    wire tlMasterXbar_monitor__GEN_54 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h3; 
    wire tlMasterXbar_monitor__GEN_55 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'h3|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_56 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_57 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_58 = tlMasterXbar_monitor_io_in_a_bits_param <=3'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_59 = tlMasterXbar_monitor_io_in_a_bits_mask == tlMasterXbar_monitor_mask ==1'h0; 
    wire tlMasterXbar_monitor__GEN_60 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor__GEN_61 =((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_a_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_a_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_a_bits_size & tlMasterXbar_monitor_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_62 = tlMasterXbar_monitor_source_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_63 = tlMasterXbar_monitor_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor__GEN_64 = tlMasterXbar_monitor_io_in_a_bits_param <=3'h1==1'h0; 
    wire tlMasterXbar_monitor__GEN_65 = tlMasterXbar_monitor_io_in_a_bits_mask == tlMasterXbar_monitor_mask ==1'h0; 
    wire tlMasterXbar_monitor__GEN_66 = tlMasterXbar_monitor_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_67 = tlMasterXbar_monitor_io_in_d_bits_opcode <=3'h6==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_1_0 = tlMasterXbar_monitor_io_in_d_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_1_1 =& tlMasterXbar_monitor_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_source_ok_1 = tlMasterXbar_monitor__source_ok_WIRE_1_0 | tlMasterXbar_monitor__source_ok_WIRE_1_1 ; 
    wire tlMasterXbar_monitor_sink_ok ={1'h0, tlMasterXbar_monitor_io_in_d_bits_sink }<3'h4; 
    wire tlMasterXbar_monitor__GEN_68 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor__GEN_69 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_70 = tlMasterXbar_monitor_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_71 = tlMasterXbar_monitor_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_72 = tlMasterXbar_monitor_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_73 = tlMasterXbar_monitor_io_in_d_bits_denied ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_74 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor__GEN_75 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_76 = tlMasterXbar_monitor_sink_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_77 = tlMasterXbar_monitor_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_78 = tlMasterXbar_monitor_io_in_d_bits_param <=2'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_79 = tlMasterXbar_monitor_io_in_d_bits_param !=2'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_80 = tlMasterXbar_monitor_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_81 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor__GEN_82 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_83 = tlMasterXbar_monitor_sink_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_84 = tlMasterXbar_monitor_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_85 = tlMasterXbar_monitor_io_in_d_bits_param <=2'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_86 = tlMasterXbar_monitor_io_in_d_bits_param !=2'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_87 =( tlMasterXbar_monitor_io_in_d_bits_denied ==1'h0| tlMasterXbar_monitor_io_in_d_bits_corrupt )==1'h0; 
    wire tlMasterXbar_monitor__GEN_88 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor__GEN_89 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_90 = tlMasterXbar_monitor_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_91 = tlMasterXbar_monitor_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_92 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor__GEN_93 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_94 = tlMasterXbar_monitor_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_95 =( tlMasterXbar_monitor_io_in_d_bits_denied ==1'h0| tlMasterXbar_monitor_io_in_d_bits_corrupt )==1'h0; 
    wire tlMasterXbar_monitor__GEN_96 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor__GEN_97 = tlMasterXbar_monitor_source_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_98 = tlMasterXbar_monitor_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_99 = tlMasterXbar_monitor_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_100 = tlMasterXbar_monitor_io_in_b_bits_opcode <=3'h6==1'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_0 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'hC000000}&33'h1FC000000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_2 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_3 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address }&33'h1FFFFF000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_4 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_5 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h80000000}&33'h1F0000000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_6 =({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h60000000}&33'h1E0000000)==33'h0; 
    wire tlMasterXbar_monitor_address_ok = tlMasterXbar_monitor__address_ok_WIRE_0 | tlMasterXbar_monitor__address_ok_WIRE_1 | tlMasterXbar_monitor__address_ok_WIRE_2 | tlMasterXbar_monitor__address_ok_WIRE_3 | tlMasterXbar_monitor__address_ok_WIRE_4 | tlMasterXbar_monitor__address_ok_WIRE_5 | tlMasterXbar_monitor__address_ok_WIRE_6 ; 
    wire[26:0] tlMasterXbar_monitor__GEN_101 =27'hFFF<< tlMasterXbar_monitor_io_in_b_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_is_aligned_mask_1 =~( tlMasterXbar_monitor__GEN_101 [11:0]); 
    wire tlMasterXbar_monitor_is_aligned_1 =( tlMasterXbar_monitor_io_in_b_bits_address &{20'h0, tlMasterXbar_monitor_is_aligned_mask_1 })==32'h0; 
    wire[1:0] tlMasterXbar_monitor_mask_sizeOH_shiftAmount_1 = tlMasterXbar_monitor_io_in_b_bits_size [1:0]; 
    wire[3:0] tlMasterXbar_monitor__GEN_102 =4'h1<< tlMasterXbar_monitor_mask_sizeOH_shiftAmount_1 ; 
    wire[2:0] tlMasterXbar_monitor_mask_sizeOH_1 = tlMasterXbar_monitor__GEN_102 [2:0]|3'h1; 
    wire tlMasterXbar_monitor__GEN_103 = tlMasterXbar_monitor_io_in_b_bits_size >=4'h3; 
    wire tlMasterXbar_monitor_mask_size_3 = tlMasterXbar_monitor_mask_sizeOH_1 [2]; 
    wire tlMasterXbar_monitor_mask_bit_3 = tlMasterXbar_monitor_io_in_b_bits_address [2]; 
    wire tlMasterXbar_monitor_mask_nbit_3 = tlMasterXbar_monitor_mask_bit_3 ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq_14 = tlMasterXbar_monitor_mask_nbit_3 &1'h1; 
    wire tlMasterXbar_monitor_mask_acc_14 = tlMasterXbar_monitor__GEN_103 | tlMasterXbar_monitor_mask_size_3 & tlMasterXbar_monitor_mask_eq_14 ; 
    wire tlMasterXbar_monitor_mask_eq_15 = tlMasterXbar_monitor_mask_bit_3 &1'h1; 
    wire tlMasterXbar_monitor_mask_acc_15 = tlMasterXbar_monitor__GEN_103 | tlMasterXbar_monitor_mask_size_3 & tlMasterXbar_monitor_mask_eq_15 ; 
    wire tlMasterXbar_monitor_mask_size_4 = tlMasterXbar_monitor_mask_sizeOH_1 [1]; 
    wire tlMasterXbar_monitor_mask_bit_4 = tlMasterXbar_monitor_io_in_b_bits_address [1]; 
    wire tlMasterXbar_monitor_mask_nbit_4 = tlMasterXbar_monitor_mask_bit_4 ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq_16 = tlMasterXbar_monitor_mask_eq_14 & tlMasterXbar_monitor_mask_nbit_4 ; 
    wire tlMasterXbar_monitor_mask_acc_16 = tlMasterXbar_monitor_mask_acc_14 | tlMasterXbar_monitor_mask_size_4 & tlMasterXbar_monitor_mask_eq_16 ; 
    wire tlMasterXbar_monitor_mask_eq_17 = tlMasterXbar_monitor_mask_eq_14 & tlMasterXbar_monitor_mask_bit_4 ; 
    wire tlMasterXbar_monitor_mask_acc_17 = tlMasterXbar_monitor_mask_acc_14 | tlMasterXbar_monitor_mask_size_4 & tlMasterXbar_monitor_mask_eq_17 ; 
    wire tlMasterXbar_monitor_mask_eq_18 = tlMasterXbar_monitor_mask_eq_15 & tlMasterXbar_monitor_mask_nbit_4 ; 
    wire tlMasterXbar_monitor_mask_acc_18 = tlMasterXbar_monitor_mask_acc_15 | tlMasterXbar_monitor_mask_size_4 & tlMasterXbar_monitor_mask_eq_18 ; 
    wire tlMasterXbar_monitor_mask_eq_19 = tlMasterXbar_monitor_mask_eq_15 & tlMasterXbar_monitor_mask_bit_4 ; 
    wire tlMasterXbar_monitor_mask_acc_19 = tlMasterXbar_monitor_mask_acc_15 | tlMasterXbar_monitor_mask_size_4 & tlMasterXbar_monitor_mask_eq_19 ; 
    wire tlMasterXbar_monitor_mask_size_5 = tlMasterXbar_monitor_mask_sizeOH_1 [0]; 
    wire tlMasterXbar_monitor_mask_bit_5 = tlMasterXbar_monitor_io_in_b_bits_address [0]; 
    wire tlMasterXbar_monitor_mask_nbit_5 = tlMasterXbar_monitor_mask_bit_5 ==1'h0; 
    wire tlMasterXbar_monitor_mask_eq_20 = tlMasterXbar_monitor_mask_eq_16 & tlMasterXbar_monitor_mask_nbit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_20 = tlMasterXbar_monitor_mask_acc_16 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_20 ; 
    wire tlMasterXbar_monitor_mask_eq_21 = tlMasterXbar_monitor_mask_eq_16 & tlMasterXbar_monitor_mask_bit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_21 = tlMasterXbar_monitor_mask_acc_16 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_21 ; 
    wire tlMasterXbar_monitor_mask_eq_22 = tlMasterXbar_monitor_mask_eq_17 & tlMasterXbar_monitor_mask_nbit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_22 = tlMasterXbar_monitor_mask_acc_17 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_22 ; 
    wire tlMasterXbar_monitor_mask_eq_23 = tlMasterXbar_monitor_mask_eq_17 & tlMasterXbar_monitor_mask_bit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_23 = tlMasterXbar_monitor_mask_acc_17 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_23 ; 
    wire tlMasterXbar_monitor_mask_eq_24 = tlMasterXbar_monitor_mask_eq_18 & tlMasterXbar_monitor_mask_nbit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_24 = tlMasterXbar_monitor_mask_acc_18 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_24 ; 
    wire tlMasterXbar_monitor_mask_eq_25 = tlMasterXbar_monitor_mask_eq_18 & tlMasterXbar_monitor_mask_bit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_25 = tlMasterXbar_monitor_mask_acc_18 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_25 ; 
    wire tlMasterXbar_monitor_mask_eq_26 = tlMasterXbar_monitor_mask_eq_19 & tlMasterXbar_monitor_mask_nbit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_26 = tlMasterXbar_monitor_mask_acc_19 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_26 ; 
    wire tlMasterXbar_monitor_mask_eq_27 = tlMasterXbar_monitor_mask_eq_19 & tlMasterXbar_monitor_mask_bit_5 ; 
    wire tlMasterXbar_monitor_mask_acc_27 = tlMasterXbar_monitor_mask_acc_19 | tlMasterXbar_monitor_mask_size_5 & tlMasterXbar_monitor_mask_eq_27 ; 
    wire[1:0] tlMasterXbar_monitor_mask_lo_lo_1 ={ tlMasterXbar_monitor_mask_acc_21 , tlMasterXbar_monitor_mask_acc_20 }; 
    wire[1:0] tlMasterXbar_monitor_mask_lo_hi_1 ={ tlMasterXbar_monitor_mask_acc_23 , tlMasterXbar_monitor_mask_acc_22 }; 
    wire[3:0] tlMasterXbar_monitor_mask_lo_1 ={ tlMasterXbar_monitor_mask_lo_hi_1 , tlMasterXbar_monitor_mask_lo_lo_1 }; 
    wire[1:0] tlMasterXbar_monitor_mask_hi_lo_1 ={ tlMasterXbar_monitor_mask_acc_25 , tlMasterXbar_monitor_mask_acc_24 }; 
    wire[1:0] tlMasterXbar_monitor_mask_hi_hi_1 ={ tlMasterXbar_monitor_mask_acc_27 , tlMasterXbar_monitor_mask_acc_26 }; 
    wire[3:0] tlMasterXbar_monitor_mask_hi_1 ={ tlMasterXbar_monitor_mask_hi_hi_1 , tlMasterXbar_monitor_mask_hi_lo_1 }; 
    wire[7:0] tlMasterXbar_monitor_mask_1 ={ tlMasterXbar_monitor_mask_hi_1 , tlMasterXbar_monitor_mask_lo_1 }; 
    wire tlMasterXbar_monitor__legal_source_WIRE_0 = tlMasterXbar_monitor_io_in_b_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__legal_source_WIRE_1 =& tlMasterXbar_monitor_io_in_b_bits_source ; 
    wire tlMasterXbar_monitor__legal_source_WIRE_1_0 = tlMasterXbar_monitor__legal_source_WIRE_1 |1'h0; 
    wire tlMasterXbar_monitor_legal_source = tlMasterXbar_monitor__legal_source_WIRE_1_0 == tlMasterXbar_monitor_io_in_b_bits_source ; 
    wire tlMasterXbar_monitor__GEN_104 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor__GEN_105 = tlMasterXbar_monitor_io_in_b_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_106 =& tlMasterXbar_monitor_io_in_b_bits_source ; 
    wire tlMasterXbar_monitor__GEN_107 = tlMasterXbar_monitor__GEN_105  ? 4'h6== tlMasterXbar_monitor_io_in_b_bits_size :1'h0; 
    wire tlMasterXbar_monitor__GEN_108 =( tlMasterXbar_monitor__GEN_107 &((4'h0<= tlMasterXbar_monitor_io_in_b_bits_size & tlMasterXbar_monitor_io_in_b_bits_size <=4'hC|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_b_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_b_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_109 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_110 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_111 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_112 = tlMasterXbar_monitor_io_in_b_bits_param <=2'h2==1'h0; 
    wire tlMasterXbar_monitor__GEN_113 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_114 = tlMasterXbar_monitor_io_in_b_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_115 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor__GEN_116 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_117 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_118 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_119 = tlMasterXbar_monitor_io_in_b_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_120 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_121 = tlMasterXbar_monitor_io_in_b_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_122 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor__GEN_123 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_124 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_125 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_126 = tlMasterXbar_monitor_io_in_b_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_127 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_128 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor__GEN_129 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_130 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_131 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_132 = tlMasterXbar_monitor_io_in_b_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_133 =( tlMasterXbar_monitor_io_in_b_bits_mask &~ tlMasterXbar_monitor_mask_1 )==8'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_134 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor__GEN_135 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_136 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_137 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_138 ={1'h0, tlMasterXbar_monitor_io_in_b_bits_param }<=3'h4==1'h0; 
    wire tlMasterXbar_monitor__GEN_139 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_140 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h3; 
    wire tlMasterXbar_monitor__GEN_141 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_142 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_143 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_144 ={1'h0, tlMasterXbar_monitor_io_in_b_bits_param }<=3'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_145 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_146 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_io_in_b_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor__GEN_147 = tlMasterXbar_monitor_address_ok ==1'h0; 
    wire tlMasterXbar_monitor__GEN_148 = tlMasterXbar_monitor_legal_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_149 = tlMasterXbar_monitor_is_aligned_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_150 = tlMasterXbar_monitor_io_in_b_bits_mask == tlMasterXbar_monitor_mask_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_151 = tlMasterXbar_monitor_io_in_b_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_152 = tlMasterXbar_monitor_io_in_c_bits_opcode <=3'h7==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_2_0 = tlMasterXbar_monitor_io_in_c_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__source_ok_WIRE_2_1 =& tlMasterXbar_monitor_io_in_c_bits_source ; 
    wire tlMasterXbar_monitor_source_ok_2 = tlMasterXbar_monitor__source_ok_WIRE_2_0 | tlMasterXbar_monitor__source_ok_WIRE_2_1 ; 
    wire[26:0] tlMasterXbar_monitor__GEN_153 =27'hFFF<< tlMasterXbar_monitor_io_in_c_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_is_aligned_mask_2 =~( tlMasterXbar_monitor__GEN_153 [11:0]); 
    wire tlMasterXbar_monitor_is_aligned_2 =( tlMasterXbar_monitor_io_in_c_bits_address &{20'h0, tlMasterXbar_monitor_is_aligned_mask_2 })==32'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_0 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_1 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'hC000000}&33'h1FC000000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_2 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_3 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address }&33'h1FFFFF000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_4 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_5 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h80000000}&33'h1F0000000)==33'h0; 
    wire tlMasterXbar_monitor__address_ok_WIRE_1_6 =({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h60000000}&33'h1E0000000)==33'h0; 
    wire tlMasterXbar_monitor_address_ok_1 = tlMasterXbar_monitor__address_ok_WIRE_1_0 | tlMasterXbar_monitor__address_ok_WIRE_1_1 | tlMasterXbar_monitor__address_ok_WIRE_1_2 | tlMasterXbar_monitor__address_ok_WIRE_1_3 | tlMasterXbar_monitor__address_ok_WIRE_1_4 | tlMasterXbar_monitor__address_ok_WIRE_1_5 | tlMasterXbar_monitor__address_ok_WIRE_1_6 ; 
    wire tlMasterXbar_monitor__GEN_154 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor__GEN_155 = tlMasterXbar_monitor_address_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_156 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_157 = tlMasterXbar_monitor_io_in_c_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_158 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_159 = tlMasterXbar_monitor_io_in_c_bits_param <=3'h5==1'h0; 
    wire tlMasterXbar_monitor__GEN_160 = tlMasterXbar_monitor_io_in_c_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_161 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor__GEN_162 = tlMasterXbar_monitor_address_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_163 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_164 = tlMasterXbar_monitor_io_in_c_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_165 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_166 = tlMasterXbar_monitor_io_in_c_bits_param <=3'h5==1'h0; 
    wire tlMasterXbar_monitor__GEN_167 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor__GEN_168 =((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_c_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_c_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_169 = tlMasterXbar_monitor_io_in_c_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_170 =& tlMasterXbar_monitor_io_in_c_bits_source ; 
    wire tlMasterXbar_monitor__GEN_171 = tlMasterXbar_monitor__GEN_169  ? 4'h6== tlMasterXbar_monitor_io_in_c_bits_size :1'h0; 
    wire tlMasterXbar_monitor__GEN_172 =( tlMasterXbar_monitor__GEN_171 &((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'hC|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_c_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_173 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_174 = tlMasterXbar_monitor_io_in_c_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_175 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_176 = tlMasterXbar_monitor_io_in_c_bits_param <=3'h5==1'h0; 
    wire tlMasterXbar_monitor__GEN_177 = tlMasterXbar_monitor_io_in_c_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_178 = tlMasterXbar_monitor_io_in_c_valid &(& tlMasterXbar_monitor_io_in_c_bits_opcode ); 
    wire tlMasterXbar_monitor__GEN_179 =((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'hC&( tlMasterXbar_monitor_io_in_c_bits_source ==1'h0|(& tlMasterXbar_monitor_io_in_c_bits_source ))|1'h0)&((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_180 = tlMasterXbar_monitor_io_in_c_bits_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_181 =& tlMasterXbar_monitor_io_in_c_bits_source ; 
    wire tlMasterXbar_monitor__GEN_182 = tlMasterXbar_monitor__GEN_180  ? 4'h6== tlMasterXbar_monitor_io_in_c_bits_size :1'h0; 
    wire tlMasterXbar_monitor__GEN_183 =( tlMasterXbar_monitor__GEN_182 &((4'h0<= tlMasterXbar_monitor_io_in_c_bits_size & tlMasterXbar_monitor_io_in_c_bits_size <=4'hC|1'h0)&(({1'h0, tlMasterXbar_monitor_io_in_c_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_io_in_c_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor__GEN_184 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_185 = tlMasterXbar_monitor_io_in_c_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor__GEN_186 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_187 = tlMasterXbar_monitor_io_in_c_bits_param <=3'h5==1'h0; 
    wire tlMasterXbar_monitor__GEN_188 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor__GEN_189 = tlMasterXbar_monitor_address_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_190 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_191 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_192 = tlMasterXbar_monitor_io_in_c_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_193 = tlMasterXbar_monitor_io_in_c_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_194 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor__GEN_195 = tlMasterXbar_monitor_address_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_196 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_197 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_198 = tlMasterXbar_monitor_io_in_c_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_199 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor__GEN_200 = tlMasterXbar_monitor_address_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_201 = tlMasterXbar_monitor_source_ok_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_202 = tlMasterXbar_monitor_is_aligned_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_203 = tlMasterXbar_monitor_io_in_c_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_204 = tlMasterXbar_monitor_io_in_c_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_sink_ok_1 ={1'h0, tlMasterXbar_monitor_io_in_e_bits_sink }<3'h4; 
    wire tlMasterXbar_monitor__GEN_205 = tlMasterXbar_monitor_sink_ok_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_206 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_207 =27'hFFF<< tlMasterXbar_monitor_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_208 =~( tlMasterXbar_monitor__GEN_207 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_a_first_beats1_decode = tlMasterXbar_monitor__GEN_208 [11:3]; 
    wire tlMasterXbar_monitor_a_first_beats1_opdata = tlMasterXbar_monitor_io_in_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_monitor_a_first_beats1 = tlMasterXbar_monitor_a_first_beats1_opdata  ?  tlMasterXbar_monitor_a_first_beats1_decode :9'h0; reg[8:0] tlMasterXbar_monitor_a_first_counter ; 
    wire[9:0] tlMasterXbar_monitor__GEN_209 ={1'h0, tlMasterXbar_monitor_a_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_a_first_counter1 = tlMasterXbar_monitor__GEN_209 [8:0]; 
    wire tlMasterXbar_monitor_a_first = tlMasterXbar_monitor_a_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_a_first_last = tlMasterXbar_monitor_a_first_counter ==9'h1| tlMasterXbar_monitor_a_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_a_first_done = tlMasterXbar_monitor_a_first_last & tlMasterXbar_monitor__GEN_206 ; 
    wire[8:0] tlMasterXbar_monitor_a_first_count = tlMasterXbar_monitor_a_first_beats1 &~ tlMasterXbar_monitor_a_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode ; reg[2:0] tlMasterXbar_monitor_param ; reg[3:0] tlMasterXbar_monitor_size ; 
    reg tlMasterXbar_monitor_source ; reg[31:0] tlMasterXbar_monitor_address ; 
    wire tlMasterXbar_monitor__GEN_210 = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first ==1'h0; 
    wire tlMasterXbar_monitor__GEN_211 = tlMasterXbar_monitor_io_in_a_bits_opcode == tlMasterXbar_monitor_opcode ==1'h0; 
    wire tlMasterXbar_monitor__GEN_212 = tlMasterXbar_monitor_io_in_a_bits_param == tlMasterXbar_monitor_param ==1'h0; 
    wire tlMasterXbar_monitor__GEN_213 = tlMasterXbar_monitor_io_in_a_bits_size == tlMasterXbar_monitor_size ==1'h0; 
    wire tlMasterXbar_monitor__GEN_214 = tlMasterXbar_monitor_io_in_a_bits_source == tlMasterXbar_monitor_source ==1'h0; 
    wire tlMasterXbar_monitor__GEN_215 = tlMasterXbar_monitor_io_in_a_bits_address == tlMasterXbar_monitor_address ==1'h0; 
    wire tlMasterXbar_monitor__GEN_216 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first ; 
    wire tlMasterXbar_monitor__GEN_217 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_218 =27'hFFF<< tlMasterXbar_monitor_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_219 =~( tlMasterXbar_monitor__GEN_218 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_decode = tlMasterXbar_monitor__GEN_219 [11:3]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1 = tlMasterXbar_monitor_d_first_beats1_opdata  ?  tlMasterXbar_monitor_d_first_beats1_decode :9'h0; reg[8:0] tlMasterXbar_monitor_d_first_counter ; 
    wire[9:0] tlMasterXbar_monitor__GEN_220 ={1'h0, tlMasterXbar_monitor_d_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_d_first_counter1 = tlMasterXbar_monitor__GEN_220 [8:0]; 
    wire tlMasterXbar_monitor_d_first = tlMasterXbar_monitor_d_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_d_first_last = tlMasterXbar_monitor_d_first_counter ==9'h1| tlMasterXbar_monitor_d_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_done = tlMasterXbar_monitor_d_first_last & tlMasterXbar_monitor__GEN_217 ; 
    wire[8:0] tlMasterXbar_monitor_d_first_count = tlMasterXbar_monitor_d_first_beats1 &~ tlMasterXbar_monitor_d_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode_1 ; reg[1:0] tlMasterXbar_monitor_param_1 ; reg[3:0] tlMasterXbar_monitor_size_1 ; 
    reg tlMasterXbar_monitor_source_1 ; reg[1:0] tlMasterXbar_monitor_sink ; 
    reg tlMasterXbar_monitor_denied ; 
    wire tlMasterXbar_monitor__GEN_221 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first ==1'h0; 
    wire tlMasterXbar_monitor__GEN_222 = tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_opcode_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_223 = tlMasterXbar_monitor_io_in_d_bits_param == tlMasterXbar_monitor_param_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_224 = tlMasterXbar_monitor_io_in_d_bits_size == tlMasterXbar_monitor_size_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_225 = tlMasterXbar_monitor_io_in_d_bits_source == tlMasterXbar_monitor_source_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_226 = tlMasterXbar_monitor_io_in_d_bits_sink == tlMasterXbar_monitor_sink ==1'h0; 
    wire tlMasterXbar_monitor__GEN_227 = tlMasterXbar_monitor_io_in_d_bits_denied == tlMasterXbar_monitor_denied ==1'h0; 
    wire tlMasterXbar_monitor__GEN_228 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first ; 
    wire tlMasterXbar_monitor__GEN_229 = tlMasterXbar_monitor_io_in_b_ready & tlMasterXbar_monitor_io_in_b_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_230 =27'hFFF<< tlMasterXbar_monitor_io_in_b_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_231 =~( tlMasterXbar_monitor__GEN_230 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_b_first_beats1_decode = tlMasterXbar_monitor__GEN_231 [11:3]; 
    wire tlMasterXbar_monitor_b_first_beats1_opdata = tlMasterXbar_monitor_io_in_b_bits_opcode [2]==1'h0; reg[8:0] tlMasterXbar_monitor_b_first_counter ; 
    wire[9:0] tlMasterXbar_monitor__GEN_232 ={1'h0, tlMasterXbar_monitor_b_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_b_first_counter1 = tlMasterXbar_monitor__GEN_232 [8:0]; 
    wire tlMasterXbar_monitor_b_first = tlMasterXbar_monitor_b_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_b_first_last = tlMasterXbar_monitor_b_first_counter ==9'h1| tlMasterXbar_monitor_b_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_b_first_done = tlMasterXbar_monitor_b_first_last & tlMasterXbar_monitor__GEN_229 ; 
    wire[8:0] tlMasterXbar_monitor_b_first_count = tlMasterXbar_monitor_b_first_beats1 &~ tlMasterXbar_monitor_b_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode_2 ; reg[1:0] tlMasterXbar_monitor_param_2 ; reg[3:0] tlMasterXbar_monitor_size_2 ; 
    reg tlMasterXbar_monitor_source_2 ; reg[31:0] tlMasterXbar_monitor_address_1 ; 
    wire tlMasterXbar_monitor__GEN_233 = tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_b_first ==1'h0; 
    wire tlMasterXbar_monitor__GEN_234 = tlMasterXbar_monitor_io_in_b_bits_opcode == tlMasterXbar_monitor_opcode_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_235 = tlMasterXbar_monitor_io_in_b_bits_param == tlMasterXbar_monitor_param_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_236 = tlMasterXbar_monitor_io_in_b_bits_size == tlMasterXbar_monitor_size_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_237 = tlMasterXbar_monitor_io_in_b_bits_source == tlMasterXbar_monitor_source_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_238 = tlMasterXbar_monitor_io_in_b_bits_address == tlMasterXbar_monitor_address_1 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_239 = tlMasterXbar_monitor_io_in_b_ready & tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_b_first ; 
    wire tlMasterXbar_monitor__GEN_240 = tlMasterXbar_monitor_io_in_c_ready & tlMasterXbar_monitor_io_in_c_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_241 =27'hFFF<< tlMasterXbar_monitor_io_in_c_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_242 =~( tlMasterXbar_monitor__GEN_241 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_c_first_beats1_decode = tlMasterXbar_monitor__GEN_242 [11:3]; 
    wire tlMasterXbar_monitor_c_first_beats1_opdata = tlMasterXbar_monitor_io_in_c_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_c_first_beats1 = tlMasterXbar_monitor_c_first_beats1_opdata  ?  tlMasterXbar_monitor_c_first_beats1_decode :9'h0; reg[8:0] tlMasterXbar_monitor_c_first_counter ; 
    wire[9:0] tlMasterXbar_monitor__GEN_243 ={1'h0, tlMasterXbar_monitor_c_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_c_first_counter1 = tlMasterXbar_monitor__GEN_243 [8:0]; 
    wire tlMasterXbar_monitor_c_first = tlMasterXbar_monitor_c_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_c_first_last = tlMasterXbar_monitor_c_first_counter ==9'h1| tlMasterXbar_monitor_c_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_c_first_done = tlMasterXbar_monitor_c_first_last & tlMasterXbar_monitor__GEN_240 ; 
    wire[8:0] tlMasterXbar_monitor_c_first_count = tlMasterXbar_monitor_c_first_beats1 &~ tlMasterXbar_monitor_c_first_counter1 ; reg[2:0] tlMasterXbar_monitor_opcode_3 ; reg[2:0] tlMasterXbar_monitor_param_3 ; reg[3:0] tlMasterXbar_monitor_size_3 ; 
    reg tlMasterXbar_monitor_source_3 ; reg[31:0] tlMasterXbar_monitor_address_2 ; 
    wire tlMasterXbar_monitor__GEN_244 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_c_first ==1'h0; 
    wire tlMasterXbar_monitor__GEN_245 = tlMasterXbar_monitor_io_in_c_bits_opcode == tlMasterXbar_monitor_opcode_3 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_246 = tlMasterXbar_monitor_io_in_c_bits_param == tlMasterXbar_monitor_param_3 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_247 = tlMasterXbar_monitor_io_in_c_bits_size == tlMasterXbar_monitor_size_3 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_248 = tlMasterXbar_monitor_io_in_c_bits_source == tlMasterXbar_monitor_source_3 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_249 = tlMasterXbar_monitor_io_in_c_bits_address == tlMasterXbar_monitor_address_2 ==1'h0; 
    wire tlMasterXbar_monitor__GEN_250 = tlMasterXbar_monitor_io_in_c_ready & tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_c_first ; reg[1:0] tlMasterXbar_monitor_inflight ; reg[7:0] tlMasterXbar_monitor_inflight_opcodes ; reg[15:0] tlMasterXbar_monitor_inflight_sizes ; 
    wire tlMasterXbar_monitor__GEN_251 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_252 =27'hFFF<< tlMasterXbar_monitor_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_253 =~( tlMasterXbar_monitor__GEN_252 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_a_first_beats1_decode_1 = tlMasterXbar_monitor__GEN_253 [11:3]; 
    wire tlMasterXbar_monitor_a_first_beats1_opdata_1 = tlMasterXbar_monitor_io_in_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_monitor_a_first_beats1_1 = tlMasterXbar_monitor_a_first_beats1_opdata_1  ?  tlMasterXbar_monitor_a_first_beats1_decode_1 :9'h0; reg[8:0] tlMasterXbar_monitor_a_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor__GEN_254 ={1'h0, tlMasterXbar_monitor_a_first_counter_1 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_a_first_counter1_1 = tlMasterXbar_monitor__GEN_254 [8:0]; 
    wire tlMasterXbar_monitor_a_first_1 = tlMasterXbar_monitor_a_first_counter_1 ==9'h0; 
    wire tlMasterXbar_monitor_a_first_last_1 = tlMasterXbar_monitor_a_first_counter_1 ==9'h1| tlMasterXbar_monitor_a_first_beats1_1 ==9'h0; 
    wire tlMasterXbar_monitor_a_first_done_1 = tlMasterXbar_monitor_a_first_last_1 & tlMasterXbar_monitor__GEN_251 ; 
    wire[8:0] tlMasterXbar_monitor_a_first_count_1 = tlMasterXbar_monitor_a_first_beats1_1 &~ tlMasterXbar_monitor_a_first_counter1_1 ; 
    wire tlMasterXbar_monitor__GEN_255 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_256 =27'hFFF<< tlMasterXbar_monitor_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_257 =~( tlMasterXbar_monitor__GEN_256 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_decode_1 = tlMasterXbar_monitor__GEN_257 [11:3]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata_1 = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_1 = tlMasterXbar_monitor_d_first_beats1_opdata_1  ?  tlMasterXbar_monitor_d_first_beats1_decode_1 :9'h0; reg[8:0] tlMasterXbar_monitor_d_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor__GEN_258 ={1'h0, tlMasterXbar_monitor_d_first_counter_1 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_d_first_counter1_1 = tlMasterXbar_monitor__GEN_258 [8:0]; 
    wire tlMasterXbar_monitor_d_first_1 = tlMasterXbar_monitor_d_first_counter_1 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_last_1 = tlMasterXbar_monitor_d_first_counter_1 ==9'h1| tlMasterXbar_monitor_d_first_beats1_1 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_done_1 = tlMasterXbar_monitor_d_first_last_1 & tlMasterXbar_monitor__GEN_255 ; 
    wire[8:0] tlMasterXbar_monitor_d_first_count_1 = tlMasterXbar_monitor_d_first_beats1_1 &~ tlMasterXbar_monitor_d_first_counter1_1 ; 
    wire[15:0] tlMasterXbar_monitor__GEN_259 =({8'h0, tlMasterXbar_monitor_inflight_opcodes >>({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h2)}&16'hF)>>16'h1; 
    wire[3:0] tlMasterXbar_monitor_a_opcode_lookup = tlMasterXbar_monitor__GEN_259 [3:0]; 
    wire[15:0] tlMasterXbar_monitor__GEN_260 =( tlMasterXbar_monitor_inflight_sizes >>({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h3)&16'hFF)>>16'h1; 
    wire[7:0] tlMasterXbar_monitor_a_size_lookup = tlMasterXbar_monitor__GEN_260 [7:0]; 
    wire[2:0] tlMasterXbar_monitor_responseMap_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMap_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMap_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMap_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMap_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMap_5 =3'h2; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_responseMapSecondOption_5 =3'h2; 
    wire[1:0] tlMasterXbar_monitor_a_set_wo_ready = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first_1  ? 2'h1<< tlMasterXbar_monitor_io_in_a_bits_source :2'h0; 
    wire tlMasterXbar_monitor__GEN_261 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first_1 ; 
    wire[1:0] tlMasterXbar_monitor_a_set = tlMasterXbar_monitor__GEN_261  ? 2'h1<< tlMasterXbar_monitor_io_in_a_bits_source :2'h0; 
    wire[3:0] tlMasterXbar_monitor_a_opcodes_set_interm = tlMasterXbar_monitor__GEN_261  ? {1'h0, tlMasterXbar_monitor_io_in_a_bits_opcode }<<4'h1|4'h1:4'h0; 
    wire[4:0] tlMasterXbar_monitor_a_sizes_set_interm = tlMasterXbar_monitor__GEN_261  ? {1'h0, tlMasterXbar_monitor_io_in_a_bits_size }<<5'h1|5'h1:5'h0; 
    wire[18:0] tlMasterXbar_monitor__GEN_262 ={15'h0, tlMasterXbar_monitor_a_opcodes_set_interm }<<({3'h0, tlMasterXbar_monitor_io_in_a_bits_source }<<4'h2); 
    wire[7:0] tlMasterXbar_monitor_a_opcodes_set = tlMasterXbar_monitor__GEN_261  ?  tlMasterXbar_monitor__GEN_262 [7:0]:8'h0; 
    wire[19:0] tlMasterXbar_monitor__GEN_263 ={15'h0, tlMasterXbar_monitor_a_sizes_set_interm }<<({3'h0, tlMasterXbar_monitor_io_in_a_bits_source }<<4'h3); 
    wire[15:0] tlMasterXbar_monitor_a_sizes_set = tlMasterXbar_monitor__GEN_261  ?  tlMasterXbar_monitor__GEN_263 [15:0]:16'h0; 
    wire[1:0] tlMasterXbar_monitor__GEN_264 = tlMasterXbar_monitor_inflight >> tlMasterXbar_monitor_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor__GEN_265 = tlMasterXbar_monitor__GEN_264 [0]==1'h0==1'h0; 
    wire tlMasterXbar_monitor_d_release_ack = tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h6; 
    wire[1:0] tlMasterXbar_monitor_d_clr_wo_ready = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_1 & tlMasterXbar_monitor_d_release_ack ==1'h0 ? 2'h1<< tlMasterXbar_monitor_io_in_d_bits_source :2'h0; 
    wire tlMasterXbar_monitor__GEN_266 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_1 & tlMasterXbar_monitor_d_release_ack ==1'h0; 
    wire[1:0] tlMasterXbar_monitor_d_clr = tlMasterXbar_monitor__GEN_266  ? 2'h1<< tlMasterXbar_monitor_io_in_d_bits_source :2'h0; 
    wire[30:0] tlMasterXbar_monitor__GEN_267 =31'hF<<({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h2); 
    wire[7:0] tlMasterXbar_monitor_d_opcodes_clr = tlMasterXbar_monitor__GEN_266  ?  tlMasterXbar_monitor__GEN_267 [7:0]:8'h0; 
    wire[30:0] tlMasterXbar_monitor__GEN_268 =31'hFF<<({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h3); 
    wire[15:0] tlMasterXbar_monitor_d_sizes_clr = tlMasterXbar_monitor__GEN_266  ?  tlMasterXbar_monitor__GEN_268 [15:0]:16'h0; 
    wire tlMasterXbar_monitor__GEN_269 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_1 & tlMasterXbar_monitor_d_release_ack ==1'h0; 
    wire tlMasterXbar_monitor_same_cycle_resp = tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_a_first_1 & tlMasterXbar_monitor_io_in_a_bits_source == tlMasterXbar_monitor_io_in_d_bits_source ; 
    wire[1:0] tlMasterXbar_monitor__GEN_270 = tlMasterXbar_monitor_inflight >> tlMasterXbar_monitor_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor__GEN_271 =( tlMasterXbar_monitor__GEN_270 [0]| tlMasterXbar_monitor_same_cycle_resp )==1'h0; 
    wire tlMasterXbar_monitor__GEN_272 = tlMasterXbar_monitor__GEN_269 & tlMasterXbar_monitor_same_cycle_resp ; reg[2:0] tlMasterXbar_monitor_casez_tmp ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_6 ;
              default : 
                  tlMasterXbar_monitor_casez_tmp  = tlMasterXbar_monitor_responseMap_7 ;endcase
         end
  reg[2:0] tlMasterXbar_monitor_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_6 ;
              default : 
                  tlMasterXbar_monitor_casez_tmp_0  = tlMasterXbar_monitor_responseMapSecondOption_7 ;endcase
         end
    wire tlMasterXbar_monitor__GEN_273 =( tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp | tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_0 )==1'h0; 
    wire tlMasterXbar_monitor__GEN_274 = tlMasterXbar_monitor_io_in_a_bits_size == tlMasterXbar_monitor_io_in_d_bits_size ==1'h0; 
    wire tlMasterXbar_monitor__GEN_275 = tlMasterXbar_monitor__GEN_269 &~ tlMasterXbar_monitor_same_cycle_resp ; reg[2:0] tlMasterXbar_monitor_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_6 ;
              default : 
                  tlMasterXbar_monitor_casez_tmp_1  = tlMasterXbar_monitor_responseMap_7 ;endcase
         end
  reg[2:0] tlMasterXbar_monitor_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_6 ;
              default : 
                  tlMasterXbar_monitor_casez_tmp_2  = tlMasterXbar_monitor_responseMapSecondOption_7 ;endcase
         end
    wire tlMasterXbar_monitor__GEN_276 =( tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_1 | tlMasterXbar_monitor_io_in_d_bits_opcode == tlMasterXbar_monitor_casez_tmp_2 )==1'h0; 
    wire tlMasterXbar_monitor__GEN_277 ={4'h0, tlMasterXbar_monitor_io_in_d_bits_size }== tlMasterXbar_monitor_a_size_lookup ==1'h0; 
    wire tlMasterXbar_monitor__GEN_278 =( tlMasterXbar_monitor_io_in_d_ready ==1'h0| tlMasterXbar_monitor_io_in_a_ready )==1'h0; 
    wire tlMasterXbar_monitor__GEN_279 =( tlMasterXbar_monitor_a_set_wo_ready != tlMasterXbar_monitor_d_clr_wo_ready |(| tlMasterXbar_monitor_a_set_wo_ready )==1'h0)==1'h0; reg[31:0] tlMasterXbar_monitor_watchdog ;  
    wire tlMasterXbar_monitor__GEN_280 =((| tlMasterXbar_monitor_inflight )==1'h0| tlMasterXbar_monitor__plusarg_reader_out ==32'h0| tlMasterXbar_monitor_watchdog < tlMasterXbar_monitor__plusarg_reader_out )==1'h0; 
    wire[32:0] tlMasterXbar_monitor__GEN_281 ={1'h0, tlMasterXbar_monitor_watchdog }+33'h1; 
    wire tlMasterXbar_monitor__GEN_282 = tlMasterXbar_monitor_io_in_a_ready & tlMasterXbar_monitor_io_in_a_valid | tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; reg[1:0] tlMasterXbar_monitor_inflight_1 ; reg[7:0] tlMasterXbar_monitor_inflight_opcodes_1 ; reg[15:0] tlMasterXbar_monitor_inflight_sizes_1 ; 
    wire tlMasterXbar_monitor__GEN_283 = tlMasterXbar_monitor_io_in_c_ready & tlMasterXbar_monitor_io_in_c_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_284 =27'hFFF<< tlMasterXbar_monitor_io_in_c_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_285 =~( tlMasterXbar_monitor__GEN_284 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_c_first_beats1_decode_1 = tlMasterXbar_monitor__GEN_285 [11:3]; 
    wire tlMasterXbar_monitor_c_first_beats1_opdata_1 = tlMasterXbar_monitor_io_in_c_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_c_first_beats1_1 = tlMasterXbar_monitor_c_first_beats1_opdata_1  ?  tlMasterXbar_monitor_c_first_beats1_decode_1 :9'h0; reg[8:0] tlMasterXbar_monitor_c_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor__GEN_286 ={1'h0, tlMasterXbar_monitor_c_first_counter_1 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_c_first_counter1_1 = tlMasterXbar_monitor__GEN_286 [8:0]; 
    wire tlMasterXbar_monitor_c_first_1 = tlMasterXbar_monitor_c_first_counter_1 ==9'h0; 
    wire tlMasterXbar_monitor_c_first_last_1 = tlMasterXbar_monitor_c_first_counter_1 ==9'h1| tlMasterXbar_monitor_c_first_beats1_1 ==9'h0; 
    wire tlMasterXbar_monitor_c_first_done_1 = tlMasterXbar_monitor_c_first_last_1 & tlMasterXbar_monitor__GEN_283 ; 
    wire[8:0] tlMasterXbar_monitor_c_first_count_1 = tlMasterXbar_monitor_c_first_beats1_1 &~ tlMasterXbar_monitor_c_first_counter1_1 ; 
    wire tlMasterXbar_monitor__GEN_287 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_288 =27'hFFF<< tlMasterXbar_monitor_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_289 =~( tlMasterXbar_monitor__GEN_288 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_decode_2 = tlMasterXbar_monitor__GEN_289 [11:3]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata_2 = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_2 = tlMasterXbar_monitor_d_first_beats1_opdata_2  ?  tlMasterXbar_monitor_d_first_beats1_decode_2 :9'h0; reg[8:0] tlMasterXbar_monitor_d_first_counter_2 ; 
    wire[9:0] tlMasterXbar_monitor__GEN_290 ={1'h0, tlMasterXbar_monitor_d_first_counter_2 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_d_first_counter1_2 = tlMasterXbar_monitor__GEN_290 [8:0]; 
    wire tlMasterXbar_monitor_d_first_2 = tlMasterXbar_monitor_d_first_counter_2 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_last_2 = tlMasterXbar_monitor_d_first_counter_2 ==9'h1| tlMasterXbar_monitor_d_first_beats1_2 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_done_2 = tlMasterXbar_monitor_d_first_last_2 & tlMasterXbar_monitor__GEN_287 ; 
    wire[8:0] tlMasterXbar_monitor_d_first_count_2 = tlMasterXbar_monitor_d_first_beats1_2 &~ tlMasterXbar_monitor_d_first_counter1_2 ; 
    wire[15:0] tlMasterXbar_monitor__GEN_291 =({8'h0, tlMasterXbar_monitor_inflight_opcodes_1 >>({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h2)}&16'hF)>>16'h1; 
    wire[3:0] tlMasterXbar_monitor_c_opcode_lookup = tlMasterXbar_monitor__GEN_291 [3:0]; 
    wire[15:0] tlMasterXbar_monitor__GEN_292 =( tlMasterXbar_monitor_inflight_sizes_1 >>({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h3)&16'hFF)>>16'h1; 
    wire[7:0] tlMasterXbar_monitor_c_size_lookup = tlMasterXbar_monitor__GEN_292 [7:0]; 
    wire[1:0] tlMasterXbar_monitor_c_set_wo_ready = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_c_first_1 & tlMasterXbar_monitor_io_in_c_bits_opcode [2]& tlMasterXbar_monitor_io_in_c_bits_opcode [1] ? 2'h1<< tlMasterXbar_monitor_io_in_c_bits_source :2'h0; 
    wire tlMasterXbar_monitor__GEN_293 = tlMasterXbar_monitor_io_in_c_ready & tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_c_first_1 & tlMasterXbar_monitor_io_in_c_bits_opcode [2]& tlMasterXbar_monitor_io_in_c_bits_opcode [1]; 
    wire[1:0] tlMasterXbar_monitor_c_set = tlMasterXbar_monitor__GEN_293  ? 2'h1<< tlMasterXbar_monitor_io_in_c_bits_source :2'h0; 
    wire[3:0] tlMasterXbar_monitor_c_opcodes_set_interm = tlMasterXbar_monitor__GEN_293  ? {1'h0, tlMasterXbar_monitor_io_in_c_bits_opcode }<<4'h1|4'h1:4'h0; 
    wire[4:0] tlMasterXbar_monitor_c_sizes_set_interm = tlMasterXbar_monitor__GEN_293  ? {1'h0, tlMasterXbar_monitor_io_in_c_bits_size }<<5'h1|5'h1:5'h0; 
    wire[18:0] tlMasterXbar_monitor__GEN_294 ={15'h0, tlMasterXbar_monitor_c_opcodes_set_interm }<<({3'h0, tlMasterXbar_monitor_io_in_c_bits_source }<<4'h2); 
    wire[7:0] tlMasterXbar_monitor_c_opcodes_set = tlMasterXbar_monitor__GEN_293  ?  tlMasterXbar_monitor__GEN_294 [7:0]:8'h0; 
    wire[19:0] tlMasterXbar_monitor__GEN_295 ={15'h0, tlMasterXbar_monitor_c_sizes_set_interm }<<({3'h0, tlMasterXbar_monitor_io_in_c_bits_source }<<4'h3); 
    wire[15:0] tlMasterXbar_monitor_c_sizes_set = tlMasterXbar_monitor__GEN_293  ?  tlMasterXbar_monitor__GEN_295 [15:0]:16'h0; 
    wire[1:0] tlMasterXbar_monitor__GEN_296 = tlMasterXbar_monitor_inflight_1 >> tlMasterXbar_monitor_io_in_c_bits_source ; 
    wire tlMasterXbar_monitor__GEN_297 = tlMasterXbar_monitor__GEN_296 [0]==1'h0==1'h0; 
    wire tlMasterXbar_monitor_c_probe_ack = tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h4| tlMasterXbar_monitor_io_in_c_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor_d_release_ack_1 = tlMasterXbar_monitor_io_in_d_bits_opcode ==3'h6; 
    wire[1:0] tlMasterXbar_monitor_d_clr_wo_ready_1 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_d_release_ack_1  ? 2'h1<< tlMasterXbar_monitor_io_in_d_bits_source :2'h0; 
    wire tlMasterXbar_monitor__GEN_298 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_d_release_ack_1 ; 
    wire[1:0] tlMasterXbar_monitor_d_clr_1 = tlMasterXbar_monitor__GEN_298  ? 2'h1<< tlMasterXbar_monitor_io_in_d_bits_source :2'h0; 
    wire[30:0] tlMasterXbar_monitor__GEN_299 =31'hF<<({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h2); 
    wire[7:0] tlMasterXbar_monitor_d_opcodes_clr_1 = tlMasterXbar_monitor__GEN_298  ?  tlMasterXbar_monitor__GEN_299 [7:0]:8'h0; 
    wire[30:0] tlMasterXbar_monitor__GEN_300 =31'hFF<<({3'h0, tlMasterXbar_monitor_io_in_d_bits_source }<<4'h3); 
    wire[15:0] tlMasterXbar_monitor_d_sizes_clr_1 = tlMasterXbar_monitor__GEN_298  ?  tlMasterXbar_monitor__GEN_300 [15:0]:16'h0; 
    wire tlMasterXbar_monitor__GEN_301 = tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_d_release_ack_1 ; 
    wire tlMasterXbar_monitor_same_cycle_resp_1 = tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_c_first_1 & tlMasterXbar_monitor_io_in_c_bits_opcode [2]& tlMasterXbar_monitor_io_in_c_bits_opcode [1]& tlMasterXbar_monitor_io_in_c_bits_source == tlMasterXbar_monitor_io_in_d_bits_source ; 
    wire[1:0] tlMasterXbar_monitor__GEN_302 = tlMasterXbar_monitor_inflight_1 >> tlMasterXbar_monitor_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor__GEN_303 =( tlMasterXbar_monitor__GEN_302 [0]| tlMasterXbar_monitor_same_cycle_resp_1 )==1'h0; 
    wire tlMasterXbar_monitor__GEN_304 = tlMasterXbar_monitor_io_in_d_bits_size == tlMasterXbar_monitor_io_in_c_bits_size ==1'h0; 
    wire tlMasterXbar_monitor__GEN_305 ={4'h0, tlMasterXbar_monitor_io_in_d_bits_size }== tlMasterXbar_monitor_c_size_lookup ==1'h0; 
    wire tlMasterXbar_monitor__GEN_306 =( tlMasterXbar_monitor_io_in_d_ready ==1'h0| tlMasterXbar_monitor_io_in_c_ready )==1'h0; 
    wire tlMasterXbar_monitor__GEN_307 = tlMasterXbar_monitor_c_set_wo_ready != tlMasterXbar_monitor_d_clr_wo_ready_1 ==1'h0; reg[31:0] tlMasterXbar_monitor_watchdog_1 ;  
    wire tlMasterXbar_monitor__GEN_308 =((| tlMasterXbar_monitor_inflight_1 )==1'h0| tlMasterXbar_monitor__plusarg_reader_1_out ==32'h0| tlMasterXbar_monitor_watchdog_1 < tlMasterXbar_monitor__plusarg_reader_1_out )==1'h0; 
    wire[32:0] tlMasterXbar_monitor__GEN_309 ={1'h0, tlMasterXbar_monitor_watchdog_1 }+33'h1; 
    wire tlMasterXbar_monitor__GEN_310 = tlMasterXbar_monitor_io_in_c_ready & tlMasterXbar_monitor_io_in_c_valid | tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; reg[3:0] tlMasterXbar_monitor_inflight_2 ; 
    wire tlMasterXbar_monitor__GEN_311 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor__GEN_312 =27'hFFF<< tlMasterXbar_monitor_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor__GEN_313 =~( tlMasterXbar_monitor__GEN_312 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_decode_3 = tlMasterXbar_monitor__GEN_313 [11:3]; 
    wire tlMasterXbar_monitor_d_first_beats1_opdata_3 = tlMasterXbar_monitor_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_d_first_beats1_3 = tlMasterXbar_monitor_d_first_beats1_opdata_3  ?  tlMasterXbar_monitor_d_first_beats1_decode_3 :9'h0; reg[8:0] tlMasterXbar_monitor_d_first_counter_3 ; 
    wire[9:0] tlMasterXbar_monitor__GEN_314 ={1'h0, tlMasterXbar_monitor_d_first_counter_3 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_d_first_counter1_3 = tlMasterXbar_monitor__GEN_314 [8:0]; 
    wire tlMasterXbar_monitor_d_first_3 = tlMasterXbar_monitor_d_first_counter_3 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_last_3 = tlMasterXbar_monitor_d_first_counter_3 ==9'h1| tlMasterXbar_monitor_d_first_beats1_3 ==9'h0; 
    wire tlMasterXbar_monitor_d_first_done_3 = tlMasterXbar_monitor_d_first_last_3 & tlMasterXbar_monitor__GEN_311 ; 
    wire[8:0] tlMasterXbar_monitor_d_first_count_3 = tlMasterXbar_monitor_d_first_beats1_3 &~ tlMasterXbar_monitor_d_first_counter1_3 ; 
    wire tlMasterXbar_monitor__GEN_315 = tlMasterXbar_monitor_io_in_d_ready & tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_3 & tlMasterXbar_monitor_io_in_d_bits_opcode [2]& tlMasterXbar_monitor_io_in_d_bits_opcode [1]==1'h0; 
    wire[3:0] tlMasterXbar_monitor_d_set = tlMasterXbar_monitor__GEN_315  ? 4'h1<< tlMasterXbar_monitor_io_in_d_bits_sink :4'h0; 
    wire[3:0] tlMasterXbar_monitor__GEN_316 = tlMasterXbar_monitor_inflight_2 >> tlMasterXbar_monitor_io_in_d_bits_sink ; 
    wire tlMasterXbar_monitor__GEN_317 = tlMasterXbar_monitor__GEN_316 [0]==1'h0==1'h0; 
    wire tlMasterXbar_monitor__GEN_318 = tlMasterXbar_monitor_io_in_e_ready & tlMasterXbar_monitor_io_in_e_valid ; 
    wire[3:0] tlMasterXbar_monitor_e_clr = tlMasterXbar_monitor__GEN_318  ? 4'h1<< tlMasterXbar_monitor_io_in_e_bits_sink :4'h0; 
    wire[3:0] tlMasterXbar_monitor__GEN_319 =( tlMasterXbar_monitor_d_set | tlMasterXbar_monitor_inflight_2 )>> tlMasterXbar_monitor_io_in_e_bits_sink ; 
    wire tlMasterXbar_monitor__GEN_320 = tlMasterXbar_monitor__GEN_319 [0]==1'h0; 
  always @( posedge  tlMasterXbar_monitor_clock )
         begin 
             if ( tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_4 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_8 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_9 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_10 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_11 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_12 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_13 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_3 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_14 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_16 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_20 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_21 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_22 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_23 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_24 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_25 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_26 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_15 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_27 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_29 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_30 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_31 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_32 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_33 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_34 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_28 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_35 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_37 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_38 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_39 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_40 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_36 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_41 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_42 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_43 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_42 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_44 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_42 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_45 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_42 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_46 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_42 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_47 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_48 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_49 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_48 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_50 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_48 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_51 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_48 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_52 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_48 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_53 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_54 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_55 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_54 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_56 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_54 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_57 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_54 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_58 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_54 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_59 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_61 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_62 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_63 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_64 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_65 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_60 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_66 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_67 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_68 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_69 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_68 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_70 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_68 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_71 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_68 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_72 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_68 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_73 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_75 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_76 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_77 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_78 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_79 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_74 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_80 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_82 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_83 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_84 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_85 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_86 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_81 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_87 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_88 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_89 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_88 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_90 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_88 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_91 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_92 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_93 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_92 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_94 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_92 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_95 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_96 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_97 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_96 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_98 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_96 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_99 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is denied (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_b_valid & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_100 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_108 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries Probe type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_109 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_110 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_111 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_112 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe carries invalid cap param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_113 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_104 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_114 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Probe is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries Get type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_116 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_117 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_118 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_119 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_120 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_115 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_121 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Get is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_123 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutFull carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_124 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutFull carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_125 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutFull address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_126 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutFull carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_122 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_127 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutFull contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_129 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutPartial carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_130 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutPartial carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_131 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_132 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutPartial carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_128 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_133 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries Arithmetic type unsupported by master (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_135 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Arithmetic carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_136 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Arithmetic carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_137 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_138 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_134 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_139 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries Logical type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_141 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Logical carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_142 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Logical carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_143 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Logical address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_144 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_140 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_145 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Logical contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'B' channel carries Hint type unsupported by client (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_147 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Hint carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_148 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Hint carries source that is not first source (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_149 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Hint address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_150 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Hint contains invalid mask (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_146 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_151 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel Hint is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_152 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel has invalid opcode (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'C' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_155 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_156 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_157 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_158 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_159 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_154 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_160 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_161 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_162 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_161 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_163 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAckData carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_161 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_164 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAckData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_161 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_165 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_161 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_166 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ProbeAckData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_168 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel carries Release type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_172 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_173 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel Release carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_174 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel Release smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_175 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel Release address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_176 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel Release carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_167 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_177 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel Release is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_179 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel carries ReleaseData type unsupported by manager (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_183 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel carries Release from a client which does not support Probe (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_184 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ReleaseData carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_185 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ReleaseData smaller than a beat (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_186 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ReleaseData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_178 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_187 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel ReleaseData carries invalid report param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_188 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_189 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_188 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_190 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_188 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_191 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_188 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_192 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_188 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_193 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_194 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_195 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAckData carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_194 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_196 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAckData carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_194 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_197 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAckData address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_194 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_198 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_199 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_200 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel HintAck carries unmanaged address (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_199 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_201 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel HintAck carries invalid source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_199 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_202 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel HintAck address not aligned to size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_199 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_203 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel HintAck carries invalid param (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_199 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_204 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel HintAck is corrupt (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_e_valid & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_205 )
                 begin 
                     if (1)$error("Assertion failed: 'E' channels carries invalid sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_210 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_211 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_210 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_212 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_210 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_213 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_210 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_214 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_210 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_215 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_222 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_223 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_224 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_225 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_226 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_221 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_227 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_233 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_234 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_233 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_235 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_233 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_236 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_233 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_237 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_233 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_238 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel addresss changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_244 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_245 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_244 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_246 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel param changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_244 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_247 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel size changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_244 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_248 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel source changed within multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_244 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_249 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel address changed with multibeat operation (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_261 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_265 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_269 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_271 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_272 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_273 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_272 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_274 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_275 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_276 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_275 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_277 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_1 & tlMasterXbar_monitor_a_first_1 & tlMasterXbar_monitor_io_in_a_valid & tlMasterXbar_monitor_io_in_a_bits_source == tlMasterXbar_monitor_io_in_d_bits_source & tlMasterXbar_monitor_d_release_ack ==1'h0& tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_278 )
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_279 )
                 begin 
                     if (1)$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_280 )
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_293 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_297 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_301 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_303 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_301 & tlMasterXbar_monitor_same_cycle_resp_1 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_304 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_301 &~ tlMasterXbar_monitor_same_cycle_resp_1 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_305 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_io_in_d_valid & tlMasterXbar_monitor_d_first_2 & tlMasterXbar_monitor_c_first_1 & tlMasterXbar_monitor_io_in_c_valid & tlMasterXbar_monitor_io_in_c_bits_source == tlMasterXbar_monitor_io_in_d_bits_source & tlMasterXbar_monitor_d_release_ack_1 & tlMasterXbar_monitor_c_probe_ack ==1'h0& tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_306 )
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ((| tlMasterXbar_monitor_c_set_wo_ready )& tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_307 )
                 begin 
                     if (1)$error("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_308 )
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_315 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_317 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel re-used a sink ID (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor__GEN_318 & tlMasterXbar_monitor_reset ==1'h0& tlMasterXbar_monitor__GEN_320 )
                 begin 
                     if (1)$error("Assertion failed: 'E' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/HellaCache.scala:271:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
         end
  always @( posedge  tlMasterXbar_monitor_clock )
         begin 
             if ( tlMasterXbar_monitor_reset )
                 begin  
                     tlMasterXbar_monitor_a_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_d_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_b_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_c_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_inflight  <=2'h0; 
                     tlMasterXbar_monitor_inflight_opcodes  <=8'h0; 
                     tlMasterXbar_monitor_inflight_sizes  <=16'h0; 
                     tlMasterXbar_monitor_a_first_counter_1  <=9'h0; 
                     tlMasterXbar_monitor_d_first_counter_1  <=9'h0; 
                     tlMasterXbar_monitor_watchdog  <=32'h0; 
                     tlMasterXbar_monitor_inflight_1  <=2'h0; 
                     tlMasterXbar_monitor_inflight_opcodes_1  <=8'h0; 
                     tlMasterXbar_monitor_inflight_sizes_1  <=16'h0; 
                     tlMasterXbar_monitor_c_first_counter_1  <=9'h0; 
                     tlMasterXbar_monitor_d_first_counter_2  <=9'h0; 
                     tlMasterXbar_monitor_watchdog_1  <=32'h0; 
                     tlMasterXbar_monitor_inflight_2  <=4'h0; 
                     tlMasterXbar_monitor_d_first_counter_3  <=9'h0;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_monitor__GEN_206 )
                         begin 
                             if ( tlMasterXbar_monitor_a_first ) 
                                 tlMasterXbar_monitor_a_first_counter  <= tlMasterXbar_monitor_a_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_a_first_counter  <= tlMasterXbar_monitor_a_first_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_217 )
                         begin 
                             if ( tlMasterXbar_monitor_d_first ) 
                                 tlMasterXbar_monitor_d_first_counter  <= tlMasterXbar_monitor_d_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter  <= tlMasterXbar_monitor_d_first_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_229 )
                         begin 
                             if ( tlMasterXbar_monitor_b_first ) 
                                 tlMasterXbar_monitor_b_first_counter  <= tlMasterXbar_monitor_b_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_b_first_counter  <= tlMasterXbar_monitor_b_first_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_240 )
                         begin 
                             if ( tlMasterXbar_monitor_c_first ) 
                                 tlMasterXbar_monitor_c_first_counter  <= tlMasterXbar_monitor_c_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_c_first_counter  <= tlMasterXbar_monitor_c_first_counter1 ;
                         end 
                      else 
                         begin 
                         end  
                     tlMasterXbar_monitor_inflight  <=( tlMasterXbar_monitor_inflight | tlMasterXbar_monitor_a_set )&~ tlMasterXbar_monitor_d_clr ; 
                     tlMasterXbar_monitor_inflight_opcodes  <=( tlMasterXbar_monitor_inflight_opcodes | tlMasterXbar_monitor_a_opcodes_set )&~ tlMasterXbar_monitor_d_opcodes_clr ; 
                     tlMasterXbar_monitor_inflight_sizes  <=( tlMasterXbar_monitor_inflight_sizes | tlMasterXbar_monitor_a_sizes_set )&~ tlMasterXbar_monitor_d_sizes_clr ;
                     if ( tlMasterXbar_monitor__GEN_251 )
                         begin 
                             if ( tlMasterXbar_monitor_a_first_1 ) 
                                 tlMasterXbar_monitor_a_first_counter_1  <= tlMasterXbar_monitor_a_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_a_first_counter_1  <= tlMasterXbar_monitor_a_first_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_255 )
                         begin 
                             if ( tlMasterXbar_monitor_d_first_1 ) 
                                 tlMasterXbar_monitor_d_first_counter_1  <= tlMasterXbar_monitor_d_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter_1  <= tlMasterXbar_monitor_d_first_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_282 ) 
                         tlMasterXbar_monitor_watchdog  <=32'h0;
                      else  
                         tlMasterXbar_monitor_watchdog  <= tlMasterXbar_monitor__GEN_281 [31:0]; 
                     tlMasterXbar_monitor_inflight_1  <=( tlMasterXbar_monitor_inflight_1 | tlMasterXbar_monitor_c_set )&~ tlMasterXbar_monitor_d_clr_1 ; 
                     tlMasterXbar_monitor_inflight_opcodes_1  <=( tlMasterXbar_monitor_inflight_opcodes_1 | tlMasterXbar_monitor_c_opcodes_set )&~ tlMasterXbar_monitor_d_opcodes_clr_1 ; 
                     tlMasterXbar_monitor_inflight_sizes_1  <=( tlMasterXbar_monitor_inflight_sizes_1 | tlMasterXbar_monitor_c_sizes_set )&~ tlMasterXbar_monitor_d_sizes_clr_1 ;
                     if ( tlMasterXbar_monitor__GEN_283 )
                         begin 
                             if ( tlMasterXbar_monitor_c_first_1 ) 
                                 tlMasterXbar_monitor_c_first_counter_1  <= tlMasterXbar_monitor_c_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_c_first_counter_1  <= tlMasterXbar_monitor_c_first_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_287 )
                         begin 
                             if ( tlMasterXbar_monitor_d_first_2 ) 
                                 tlMasterXbar_monitor_d_first_counter_2  <= tlMasterXbar_monitor_d_first_beats1_2 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter_2  <= tlMasterXbar_monitor_d_first_counter1_2 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor__GEN_310 ) 
                         tlMasterXbar_monitor_watchdog_1  <=32'h0;
                      else  
                         tlMasterXbar_monitor_watchdog_1  <= tlMasterXbar_monitor__GEN_309 [31:0]; 
                     tlMasterXbar_monitor_inflight_2  <=( tlMasterXbar_monitor_inflight_2 | tlMasterXbar_monitor_d_set )&~ tlMasterXbar_monitor_e_clr ;
                     if ( tlMasterXbar_monitor__GEN_311 )
                         begin 
                             if ( tlMasterXbar_monitor_d_first_3 ) 
                                 tlMasterXbar_monitor_d_first_counter_3  <= tlMasterXbar_monitor_d_first_beats1_3 ;
                              else  
                                 tlMasterXbar_monitor_d_first_counter_3  <= tlMasterXbar_monitor_d_first_counter1_3 ;
                         end 
                      else 
                         begin 
                         end 
                 end 
         end
  always @( posedge  tlMasterXbar_monitor_clock )
         begin 
             if ( tlMasterXbar_monitor__GEN_216 )
                 begin  
                     tlMasterXbar_monitor_opcode  <= tlMasterXbar_monitor_io_in_a_bits_opcode ; 
                     tlMasterXbar_monitor_param  <= tlMasterXbar_monitor_io_in_a_bits_param ; 
                     tlMasterXbar_monitor_size  <= tlMasterXbar_monitor_io_in_a_bits_size ; 
                     tlMasterXbar_monitor_source  <= tlMasterXbar_monitor_io_in_a_bits_source ; 
                     tlMasterXbar_monitor_address  <= tlMasterXbar_monitor_io_in_a_bits_address ;
                 end 
              else 
                 begin 
                 end 
             if ( tlMasterXbar_monitor__GEN_228 )
                 begin  
                     tlMasterXbar_monitor_opcode_1  <= tlMasterXbar_monitor_io_in_d_bits_opcode ; 
                     tlMasterXbar_monitor_param_1  <= tlMasterXbar_monitor_io_in_d_bits_param ; 
                     tlMasterXbar_monitor_size_1  <= tlMasterXbar_monitor_io_in_d_bits_size ; 
                     tlMasterXbar_monitor_source_1  <= tlMasterXbar_monitor_io_in_d_bits_source ; 
                     tlMasterXbar_monitor_sink  <= tlMasterXbar_monitor_io_in_d_bits_sink ; 
                     tlMasterXbar_monitor_denied  <= tlMasterXbar_monitor_io_in_d_bits_denied ;
                 end 
              else 
                 begin 
                 end 
             if ( tlMasterXbar_monitor__GEN_239 )
                 begin  
                     tlMasterXbar_monitor_opcode_2  <= tlMasterXbar_monitor_io_in_b_bits_opcode ; 
                     tlMasterXbar_monitor_param_2  <= tlMasterXbar_monitor_io_in_b_bits_param ; 
                     tlMasterXbar_monitor_size_2  <= tlMasterXbar_monitor_io_in_b_bits_size ; 
                     tlMasterXbar_monitor_source_2  <= tlMasterXbar_monitor_io_in_b_bits_source ; 
                     tlMasterXbar_monitor_address_1  <= tlMasterXbar_monitor_io_in_b_bits_address ;
                 end 
              else 
                 begin 
                 end 
             if ( tlMasterXbar_monitor__GEN_250 )
                 begin  
                     tlMasterXbar_monitor_opcode_3  <= tlMasterXbar_monitor_io_in_c_bits_opcode ; 
                     tlMasterXbar_monitor_param_3  <= tlMasterXbar_monitor_io_in_c_bits_param ; 
                     tlMasterXbar_monitor_size_3  <= tlMasterXbar_monitor_io_in_c_bits_size ; 
                     tlMasterXbar_monitor_source_3  <= tlMasterXbar_monitor_io_in_c_bits_source ; 
                     tlMasterXbar_monitor_address_2  <= tlMasterXbar_monitor_io_in_c_bits_address ;
                 end 
              else 
                 begin 
                 end 
         end
 
    assign tlMasterXbar_monitor_clock = tlMasterXbar_clock;
    assign tlMasterXbar_monitor_reset = tlMasterXbar_reset;
    assign tlMasterXbar_monitor_io_in_a_ready = tlMasterXbar_nodeIn_a_ready;
    assign tlMasterXbar_monitor_io_in_a_valid = tlMasterXbar_nodeIn_a_valid;
    assign tlMasterXbar_monitor_io_in_a_bits_opcode = tlMasterXbar_nodeIn_a_bits_opcode;
    assign tlMasterXbar_monitor_io_in_a_bits_param = tlMasterXbar_nodeIn_a_bits_param;
    assign tlMasterXbar_monitor_io_in_a_bits_size = tlMasterXbar_nodeIn_a_bits_size;
    assign tlMasterXbar_monitor_io_in_a_bits_source = tlMasterXbar_nodeIn_a_bits_source;
    assign tlMasterXbar_monitor_io_in_a_bits_address = tlMasterXbar_nodeIn_a_bits_address;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_bufferable = tlMasterXbar_nodeIn_a_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_modifiable = tlMasterXbar_nodeIn_a_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_readalloc = tlMasterXbar_nodeIn_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_writealloc = tlMasterXbar_nodeIn_a_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_privileged = tlMasterXbar_nodeIn_a_bits_user_amba_prot_privileged;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_secure = tlMasterXbar_nodeIn_a_bits_user_amba_prot_secure;
    assign tlMasterXbar_monitor_io_in_a_bits_user_amba_prot_fetch = tlMasterXbar_nodeIn_a_bits_user_amba_prot_fetch;
    assign tlMasterXbar_monitor_io_in_a_bits_mask = tlMasterXbar_nodeIn_a_bits_mask;
    assign tlMasterXbar_monitor_io_in_a_bits_data = tlMasterXbar_nodeIn_a_bits_data;
    assign tlMasterXbar_monitor_io_in_a_bits_corrupt = tlMasterXbar_nodeIn_a_bits_corrupt;
    assign tlMasterXbar_monitor_io_in_b_ready = tlMasterXbar_nodeIn_b_ready;
    assign tlMasterXbar_monitor_io_in_b_valid = tlMasterXbar_nodeIn_b_valid;
    assign tlMasterXbar_monitor_io_in_b_bits_opcode = tlMasterXbar_nodeIn_b_bits_opcode;
    assign tlMasterXbar_monitor_io_in_b_bits_param = tlMasterXbar_nodeIn_b_bits_param;
    assign tlMasterXbar_monitor_io_in_b_bits_size = tlMasterXbar_nodeIn_b_bits_size;
    assign tlMasterXbar_monitor_io_in_b_bits_source = tlMasterXbar_nodeIn_b_bits_source;
    assign tlMasterXbar_monitor_io_in_b_bits_address = tlMasterXbar_nodeIn_b_bits_address;
    assign tlMasterXbar_monitor_io_in_b_bits_mask = tlMasterXbar_nodeIn_b_bits_mask;
    assign tlMasterXbar_monitor_io_in_b_bits_data = tlMasterXbar_nodeIn_b_bits_data;
    assign tlMasterXbar_monitor_io_in_b_bits_corrupt = tlMasterXbar_nodeIn_b_bits_corrupt;
    assign tlMasterXbar_monitor_io_in_c_ready = tlMasterXbar_nodeIn_c_ready;
    assign tlMasterXbar_monitor_io_in_c_valid = tlMasterXbar_nodeIn_c_valid;
    assign tlMasterXbar_monitor_io_in_c_bits_opcode = tlMasterXbar_nodeIn_c_bits_opcode;
    assign tlMasterXbar_monitor_io_in_c_bits_param = tlMasterXbar_nodeIn_c_bits_param;
    assign tlMasterXbar_monitor_io_in_c_bits_size = tlMasterXbar_nodeIn_c_bits_size;
    assign tlMasterXbar_monitor_io_in_c_bits_source = tlMasterXbar_nodeIn_c_bits_source;
    assign tlMasterXbar_monitor_io_in_c_bits_address = tlMasterXbar_nodeIn_c_bits_address;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_bufferable = tlMasterXbar_nodeIn_c_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_modifiable = tlMasterXbar_nodeIn_c_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_readalloc = tlMasterXbar_nodeIn_c_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_writealloc = tlMasterXbar_nodeIn_c_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_privileged = tlMasterXbar_nodeIn_c_bits_user_amba_prot_privileged;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_secure = tlMasterXbar_nodeIn_c_bits_user_amba_prot_secure;
    assign tlMasterXbar_monitor_io_in_c_bits_user_amba_prot_fetch = tlMasterXbar_nodeIn_c_bits_user_amba_prot_fetch;
    assign tlMasterXbar_monitor_io_in_c_bits_data = tlMasterXbar_nodeIn_c_bits_data;
    assign tlMasterXbar_monitor_io_in_c_bits_corrupt = tlMasterXbar_nodeIn_c_bits_corrupt;
    assign tlMasterXbar_monitor_io_in_d_ready = tlMasterXbar_nodeIn_d_ready;
    assign tlMasterXbar_monitor_io_in_d_valid = tlMasterXbar_nodeIn_d_valid;
    assign tlMasterXbar_monitor_io_in_d_bits_opcode = tlMasterXbar_nodeIn_d_bits_opcode;
    assign tlMasterXbar_monitor_io_in_d_bits_param = tlMasterXbar_nodeIn_d_bits_param;
    assign tlMasterXbar_monitor_io_in_d_bits_size = tlMasterXbar_nodeIn_d_bits_size;
    assign tlMasterXbar_monitor_io_in_d_bits_source = tlMasterXbar_nodeIn_d_bits_source;
    assign tlMasterXbar_monitor_io_in_d_bits_sink = tlMasterXbar_nodeIn_d_bits_sink;
    assign tlMasterXbar_monitor_io_in_d_bits_denied = tlMasterXbar_nodeIn_d_bits_denied;
    assign tlMasterXbar_monitor_io_in_d_bits_data = tlMasterXbar_nodeIn_d_bits_data;
    assign tlMasterXbar_monitor_io_in_d_bits_corrupt = tlMasterXbar_nodeIn_d_bits_corrupt;
    assign tlMasterXbar_monitor_io_in_e_ready = tlMasterXbar_nodeIn_e_ready;
    assign tlMasterXbar_monitor_io_in_e_valid = tlMasterXbar_nodeIn_e_valid;
    assign tlMasterXbar_monitor_io_in_e_bits_sink = tlMasterXbar_nodeIn_e_bits_sink;
     
    wire tlMasterXbar_nodeIn_1_a_ready ; 
    wire tlMasterXbar_nodeIn_1_d_valid ; 
    wire[2:0] tlMasterXbar_nodeIn_1_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_nodeIn_1_d_bits_param ; 
    wire[3:0] tlMasterXbar_nodeIn_1_d_bits_size ; 
    wire[1:0] tlMasterXbar_nodeIn_1_d_bits_sink ; 
    wire tlMasterXbar_nodeIn_1_d_bits_denied ; 
    wire[63:0] tlMasterXbar_nodeIn_1_d_bits_data ; 
    wire tlMasterXbar_nodeIn_1_d_bits_corrupt ;  
    wire tlMasterXbar_monitor_1_clock;
    wire tlMasterXbar_monitor_1_reset;
    wire tlMasterXbar_monitor_1_io_in_a_ready;
    wire tlMasterXbar_monitor_1_io_in_a_valid;
    wire[2:0] tlMasterXbar_monitor_1_io_in_a_bits_opcode;
    wire[2:0] tlMasterXbar_monitor_1_io_in_a_bits_param;
    wire[3:0] tlMasterXbar_monitor_1_io_in_a_bits_size;
    wire tlMasterXbar_monitor_1_io_in_a_bits_source;
    wire[31:0] tlMasterXbar_monitor_1_io_in_a_bits_address;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_bufferable;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_modifiable;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_readalloc;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_writealloc;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_privileged;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_secure;
    wire tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_fetch;
    wire[7:0] tlMasterXbar_monitor_1_io_in_a_bits_mask;
    wire[63:0] tlMasterXbar_monitor_1_io_in_a_bits_data;
    wire tlMasterXbar_monitor_1_io_in_a_bits_corrupt;
    wire tlMasterXbar_monitor_1_io_in_d_ready;
    wire tlMasterXbar_monitor_1_io_in_d_valid;
    wire[2:0] tlMasterXbar_monitor_1_io_in_d_bits_opcode;
    wire[1:0] tlMasterXbar_monitor_1_io_in_d_bits_param;
    wire[3:0] tlMasterXbar_monitor_1_io_in_d_bits_size;
    wire tlMasterXbar_monitor_1_io_in_d_bits_source;
    wire[1:0] tlMasterXbar_monitor_1_io_in_d_bits_sink;
    wire tlMasterXbar_monitor_1_io_in_d_bits_denied;
    wire[63:0] tlMasterXbar_monitor_1_io_in_d_bits_data;
    wire tlMasterXbar_monitor_1_io_in_d_bits_corrupt;

    wire[31:0] tlMasterXbar_monitor_1__plusarg_reader_1_out ; 
    wire[31:0] tlMasterXbar_monitor_1__plusarg_reader_out ; 
    wire[8:0] tlMasterXbar_monitor_1_c_first_beats1 =9'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_0 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_first_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_first_WIRE_2_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_1 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_2 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_3 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_4 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_set_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_5 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_address =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_6 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_7 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_8 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_9 =32'h0; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_10 =32'h0; 
    wire[7:0] tlMasterXbar_monitor_1__GEN_11 =8'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_12 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_13 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_first_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_first_WIRE_2_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_14 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_15 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_16 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_17 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_set_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_18 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_data =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_19 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_20 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_21 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_22 =64'h0; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_23 =64'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_24 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_25 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_first_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_first_WIRE_2_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_26 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_27 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_28 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_29 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_set_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_30 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_size =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_31 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_32 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_33 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_34 =4'h0; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_35 =4'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_6 =3'h5; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_6 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_7 =3'h4; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_7 =3'h4; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_36 =2'h0; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_37 =2'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_38 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_39 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_40 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_2_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_2_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_41 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_42 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_43 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_44 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_45 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_46 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_47 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_48 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_49 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_50 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_opcode =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_param =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_51 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_52 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_53 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_54 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_55 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_56 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_57 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_58 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_59 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_60 =3'h0; 
    wire tlMasterXbar_monitor_1__GEN_61 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_62 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_63 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_64 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_65 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_66 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_67 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_68 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_69 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_70 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_71 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_72 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_73 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_74 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_75 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_76 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_77 =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_2_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_78 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_79 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_80 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_81 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_82 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_83 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_84 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_85 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_86 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_87 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_88 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_89 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_90 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_91 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_92 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_93 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_94 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_95 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_96 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_97 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_98 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_99 =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_100 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_101 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_102 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_103 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_104 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_105 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_106 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_107 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_108 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_109 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_110 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_111 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_112 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_113 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_114 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_115 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_116 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_117 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_118 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_119 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_120 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_121 =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_122 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_123 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_124 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_125 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_126 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_127 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_128 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_129 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_130 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_131 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_132 =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_ready =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_valid =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_ready =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_valid =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_ready =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_valid =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_ready =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_valid =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_source =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_bufferable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_modifiable =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_readalloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_writealloc =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_privileged =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_secure =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_fetch =1'h0; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_corrupt =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_133 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_134 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_135 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_136 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_137 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_138 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_139 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_140 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_141 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_142 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_143 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_144 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_145 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_146 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_147 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_148 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_149 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_150 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_151 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_152 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_153 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_154 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_155 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_156 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_157 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_158 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_159 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_160 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_161 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_162 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_163 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_164 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_165 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_166 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_167 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_168 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_169 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_170 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_171 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_172 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_173 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_174 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_175 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_176 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_177 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_178 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_179 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_180 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_181 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_182 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_183 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_184 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_185 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_186 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_187 =1'h0; 
    wire tlMasterXbar_monitor_1__GEN_188 = tlMasterXbar_monitor_1_io_in_a_bits_opcode <=3'h7==1'h0; 
    wire tlMasterXbar_monitor_1__source_ok_WIRE_0 = tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_189 =27'hFFF<< tlMasterXbar_monitor_1_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1_is_aligned_mask =~( tlMasterXbar_monitor_1__GEN_189 [11:0]); 
    wire tlMasterXbar_monitor_1_is_aligned =( tlMasterXbar_monitor_1_io_in_a_bits_address &{20'h0, tlMasterXbar_monitor_1_is_aligned_mask })==32'h0; 
    wire[1:0] tlMasterXbar_monitor_1_mask_sizeOH_shiftAmount = tlMasterXbar_monitor_1_io_in_a_bits_size [1:0]; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_190 =4'h1<< tlMasterXbar_monitor_1_mask_sizeOH_shiftAmount ; 
    wire[2:0] tlMasterXbar_monitor_1_mask_sizeOH = tlMasterXbar_monitor_1__GEN_190 [2:0]|3'h1; 
    wire tlMasterXbar_monitor_1__GEN_191 = tlMasterXbar_monitor_1_io_in_a_bits_size >=4'h3; 
    wire tlMasterXbar_monitor_1_mask_size = tlMasterXbar_monitor_1_mask_sizeOH [2]; 
    wire tlMasterXbar_monitor_1_mask_bit = tlMasterXbar_monitor_1_io_in_a_bits_address [2]; 
    wire tlMasterXbar_monitor_1_mask_nbit = tlMasterXbar_monitor_1_mask_bit ==1'h0; 
    wire tlMasterXbar_monitor_1_mask_eq = tlMasterXbar_monitor_1_mask_nbit &1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc = tlMasterXbar_monitor_1__GEN_191 | tlMasterXbar_monitor_1_mask_size & tlMasterXbar_monitor_1_mask_eq ; 
    wire tlMasterXbar_monitor_1_mask_eq_1 = tlMasterXbar_monitor_1_mask_bit &1'h1; 
    wire tlMasterXbar_monitor_1_mask_acc_1 = tlMasterXbar_monitor_1__GEN_191 | tlMasterXbar_monitor_1_mask_size & tlMasterXbar_monitor_1_mask_eq_1 ; 
    wire tlMasterXbar_monitor_1_mask_size_1 = tlMasterXbar_monitor_1_mask_sizeOH [1]; 
    wire tlMasterXbar_monitor_1_mask_bit_1 = tlMasterXbar_monitor_1_io_in_a_bits_address [1]; 
    wire tlMasterXbar_monitor_1_mask_nbit_1 = tlMasterXbar_monitor_1_mask_bit_1 ==1'h0; 
    wire tlMasterXbar_monitor_1_mask_eq_2 = tlMasterXbar_monitor_1_mask_eq & tlMasterXbar_monitor_1_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_1_mask_acc_2 = tlMasterXbar_monitor_1_mask_acc | tlMasterXbar_monitor_1_mask_size_1 & tlMasterXbar_monitor_1_mask_eq_2 ; 
    wire tlMasterXbar_monitor_1_mask_eq_3 = tlMasterXbar_monitor_1_mask_eq & tlMasterXbar_monitor_1_mask_bit_1 ; 
    wire tlMasterXbar_monitor_1_mask_acc_3 = tlMasterXbar_monitor_1_mask_acc | tlMasterXbar_monitor_1_mask_size_1 & tlMasterXbar_monitor_1_mask_eq_3 ; 
    wire tlMasterXbar_monitor_1_mask_eq_4 = tlMasterXbar_monitor_1_mask_eq_1 & tlMasterXbar_monitor_1_mask_nbit_1 ; 
    wire tlMasterXbar_monitor_1_mask_acc_4 = tlMasterXbar_monitor_1_mask_acc_1 | tlMasterXbar_monitor_1_mask_size_1 & tlMasterXbar_monitor_1_mask_eq_4 ; 
    wire tlMasterXbar_monitor_1_mask_eq_5 = tlMasterXbar_monitor_1_mask_eq_1 & tlMasterXbar_monitor_1_mask_bit_1 ; 
    wire tlMasterXbar_monitor_1_mask_acc_5 = tlMasterXbar_monitor_1_mask_acc_1 | tlMasterXbar_monitor_1_mask_size_1 & tlMasterXbar_monitor_1_mask_eq_5 ; 
    wire tlMasterXbar_monitor_1_mask_size_2 = tlMasterXbar_monitor_1_mask_sizeOH [0]; 
    wire tlMasterXbar_monitor_1_mask_bit_2 = tlMasterXbar_monitor_1_io_in_a_bits_address [0]; 
    wire tlMasterXbar_monitor_1_mask_nbit_2 = tlMasterXbar_monitor_1_mask_bit_2 ==1'h0; 
    wire tlMasterXbar_monitor_1_mask_eq_6 = tlMasterXbar_monitor_1_mask_eq_2 & tlMasterXbar_monitor_1_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_6 = tlMasterXbar_monitor_1_mask_acc_2 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_6 ; 
    wire tlMasterXbar_monitor_1_mask_eq_7 = tlMasterXbar_monitor_1_mask_eq_2 & tlMasterXbar_monitor_1_mask_bit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_7 = tlMasterXbar_monitor_1_mask_acc_2 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_7 ; 
    wire tlMasterXbar_monitor_1_mask_eq_8 = tlMasterXbar_monitor_1_mask_eq_3 & tlMasterXbar_monitor_1_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_8 = tlMasterXbar_monitor_1_mask_acc_3 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_8 ; 
    wire tlMasterXbar_monitor_1_mask_eq_9 = tlMasterXbar_monitor_1_mask_eq_3 & tlMasterXbar_monitor_1_mask_bit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_9 = tlMasterXbar_monitor_1_mask_acc_3 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_9 ; 
    wire tlMasterXbar_monitor_1_mask_eq_10 = tlMasterXbar_monitor_1_mask_eq_4 & tlMasterXbar_monitor_1_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_10 = tlMasterXbar_monitor_1_mask_acc_4 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_10 ; 
    wire tlMasterXbar_monitor_1_mask_eq_11 = tlMasterXbar_monitor_1_mask_eq_4 & tlMasterXbar_monitor_1_mask_bit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_11 = tlMasterXbar_monitor_1_mask_acc_4 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_11 ; 
    wire tlMasterXbar_monitor_1_mask_eq_12 = tlMasterXbar_monitor_1_mask_eq_5 & tlMasterXbar_monitor_1_mask_nbit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_12 = tlMasterXbar_monitor_1_mask_acc_5 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_12 ; 
    wire tlMasterXbar_monitor_1_mask_eq_13 = tlMasterXbar_monitor_1_mask_eq_5 & tlMasterXbar_monitor_1_mask_bit_2 ; 
    wire tlMasterXbar_monitor_1_mask_acc_13 = tlMasterXbar_monitor_1_mask_acc_5 | tlMasterXbar_monitor_1_mask_size_2 & tlMasterXbar_monitor_1_mask_eq_13 ; 
    wire[1:0] tlMasterXbar_monitor_1_mask_lo_lo ={ tlMasterXbar_monitor_1_mask_acc_7 , tlMasterXbar_monitor_1_mask_acc_6 }; 
    wire[1:0] tlMasterXbar_monitor_1_mask_lo_hi ={ tlMasterXbar_monitor_1_mask_acc_9 , tlMasterXbar_monitor_1_mask_acc_8 }; 
    wire[3:0] tlMasterXbar_monitor_1_mask_lo ={ tlMasterXbar_monitor_1_mask_lo_hi , tlMasterXbar_monitor_1_mask_lo_lo }; 
    wire[1:0] tlMasterXbar_monitor_1_mask_hi_lo ={ tlMasterXbar_monitor_1_mask_acc_11 , tlMasterXbar_monitor_1_mask_acc_10 }; 
    wire[1:0] tlMasterXbar_monitor_1_mask_hi_hi ={ tlMasterXbar_monitor_1_mask_acc_13 , tlMasterXbar_monitor_1_mask_acc_12 }; 
    wire[3:0] tlMasterXbar_monitor_1_mask_hi ={ tlMasterXbar_monitor_1_mask_hi_hi , tlMasterXbar_monitor_1_mask_hi_lo }; 
    wire[7:0] tlMasterXbar_monitor_1_mask ={ tlMasterXbar_monitor_1_mask_hi , tlMasterXbar_monitor_1_mask_lo }; 
    wire tlMasterXbar_monitor_1__GEN_192 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor_1__GEN_193 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_194 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_195 = tlMasterXbar_monitor_1_io_in_a_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_196 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_197 = tlMasterXbar_monitor_1_io_in_a_bits_param <=3'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_198 =~ tlMasterXbar_monitor_1_io_in_a_bits_mask ==8'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_199 = tlMasterXbar_monitor_1_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_200 = tlMasterXbar_monitor_1_io_in_a_valid &(& tlMasterXbar_monitor_1_io_in_a_bits_opcode ); 
    wire tlMasterXbar_monitor_1__GEN_201 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h6|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_202 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_203 = tlMasterXbar_monitor_1_io_in_a_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_204 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_205 = tlMasterXbar_monitor_1_io_in_a_bits_param <=3'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_206 =(| tlMasterXbar_monitor_1_io_in_a_bits_param )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_207 =~ tlMasterXbar_monitor_1_io_in_a_bits_mask ==8'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_208 = tlMasterXbar_monitor_1_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_209 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor_1__GEN_210 =(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_211 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h10000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_212 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_213 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_214 = tlMasterXbar_monitor_1_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_215 = tlMasterXbar_monitor_1_io_in_a_bits_mask == tlMasterXbar_monitor_1_mask ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_216 = tlMasterXbar_monitor_1_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_217 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor_1__GEN_218 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h8|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_219 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_220 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_221 = tlMasterXbar_monitor_1_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_222 = tlMasterXbar_monitor_1_io_in_a_bits_mask == tlMasterXbar_monitor_1_mask ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_223 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor_1__GEN_224 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0|(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h6|1'h0)&(({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h80000000}&33'h1F0000000)==33'h0)|(4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h8|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h60000000}&33'h1E0000000)==33'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_225 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_226 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_227 = tlMasterXbar_monitor_1_io_in_a_bits_param ==3'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_228 =( tlMasterXbar_monitor_1_io_in_a_bits_mask &~ tlMasterXbar_monitor_1_mask )==8'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_229 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor_1__GEN_230 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h3|1'h0)&(({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_231 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_232 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_233 = tlMasterXbar_monitor_1_io_in_a_bits_param <=3'h4==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_234 = tlMasterXbar_monitor_1_io_in_a_bits_mask == tlMasterXbar_monitor_1_mask ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_235 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h3; 
    wire tlMasterXbar_monitor_1__GEN_236 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'h3|1'h0)&(({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address }&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h2000000}&33'h1FFFF0000)==33'h0|({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'hC000000}&33'h1FC000000)==33'h0)|1'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_237 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_238 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_239 = tlMasterXbar_monitor_1_io_in_a_bits_param <=3'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_240 = tlMasterXbar_monitor_1_io_in_a_bits_mask == tlMasterXbar_monitor_1_mask ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_241 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor_1__GEN_242 =((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC& tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0|1'h0)&((4'h0<= tlMasterXbar_monitor_1_io_in_a_bits_size & tlMasterXbar_monitor_1_io_in_a_bits_size <=4'hC|1'h0)&({1'h0, tlMasterXbar_monitor_1_io_in_a_bits_address ^32'h3000}&33'h1FFFFF000)==33'h0|1'h0))==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_243 = tlMasterXbar_monitor_1__source_ok_WIRE_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_244 = tlMasterXbar_monitor_1_is_aligned ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_245 = tlMasterXbar_monitor_1_io_in_a_bits_param <=3'h1==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_246 = tlMasterXbar_monitor_1_io_in_a_bits_mask == tlMasterXbar_monitor_1_mask ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_247 = tlMasterXbar_monitor_1_io_in_a_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_248 = tlMasterXbar_monitor_1_io_in_d_bits_opcode <=3'h6==1'h0; 
    wire tlMasterXbar_monitor_1__source_ok_WIRE_1_0 = tlMasterXbar_monitor_1_io_in_d_bits_source ==1'h0; 
    wire tlMasterXbar_monitor_1_sink_ok ={1'h0, tlMasterXbar_monitor_1_io_in_d_bits_sink }<3'h4; 
    wire tlMasterXbar_monitor_1__GEN_249 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h6; 
    wire tlMasterXbar_monitor_1__GEN_250 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_251 = tlMasterXbar_monitor_1_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_252 = tlMasterXbar_monitor_1_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_253 = tlMasterXbar_monitor_1_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_254 = tlMasterXbar_monitor_1_io_in_d_bits_denied ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_255 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h4; 
    wire tlMasterXbar_monitor_1__GEN_256 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_257 = tlMasterXbar_monitor_1_sink_ok ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_258 = tlMasterXbar_monitor_1_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_259 = tlMasterXbar_monitor_1_io_in_d_bits_param <=2'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_260 = tlMasterXbar_monitor_1_io_in_d_bits_param !=2'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_261 = tlMasterXbar_monitor_1_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_262 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor_1__GEN_263 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_264 = tlMasterXbar_monitor_1_sink_ok ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_265 = tlMasterXbar_monitor_1_io_in_d_bits_size >=4'h3==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_266 = tlMasterXbar_monitor_1_io_in_d_bits_param <=2'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_267 = tlMasterXbar_monitor_1_io_in_d_bits_param !=2'h2==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_268 =( tlMasterXbar_monitor_1_io_in_d_bits_denied ==1'h0| tlMasterXbar_monitor_1_io_in_d_bits_corrupt )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_269 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h0; 
    wire tlMasterXbar_monitor_1__GEN_270 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_271 = tlMasterXbar_monitor_1_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_272 = tlMasterXbar_monitor_1_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_273 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h1; 
    wire tlMasterXbar_monitor_1__GEN_274 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_275 = tlMasterXbar_monitor_1_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_276 =( tlMasterXbar_monitor_1_io_in_d_bits_denied ==1'h0| tlMasterXbar_monitor_1_io_in_d_bits_corrupt )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_277 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h2; 
    wire tlMasterXbar_monitor_1__GEN_278 = tlMasterXbar_monitor_1__source_ok_WIRE_1_0 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_279 = tlMasterXbar_monitor_1_io_in_d_bits_param ==2'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_280 = tlMasterXbar_monitor_1_io_in_d_bits_corrupt ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_281 = tlMasterXbar_monitor_1__GEN_61 ; 
    wire tlMasterXbar_monitor_1__GEN_282 = tlMasterXbar_monitor_1__GEN_62 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_283 = tlMasterXbar_monitor_1__GEN_38 ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_284 = tlMasterXbar_monitor_1__GEN_36 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_285 = tlMasterXbar_monitor_1__GEN_24 ; 
    wire tlMasterXbar_monitor_1__GEN_286 = tlMasterXbar_monitor_1__GEN_63 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_287 = tlMasterXbar_monitor_1__GEN ; 
    wire[7:0] tlMasterXbar_monitor_1__GEN_288 = tlMasterXbar_monitor_1__GEN_11 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_289 = tlMasterXbar_monitor_1__GEN_12 ; 
    wire tlMasterXbar_monitor_1__GEN_290 = tlMasterXbar_monitor_1__GEN_64 ; 
    wire tlMasterXbar_monitor_1__GEN_291 = tlMasterXbar_monitor_1__GEN_282 ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_292 = tlMasterXbar_monitor_1__GEN_65 ; 
    wire tlMasterXbar_monitor_1__GEN_293 = tlMasterXbar_monitor_1__GEN_66 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_294 = tlMasterXbar_monitor_1__GEN_39 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_295 = tlMasterXbar_monitor_1__GEN_40 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_296 = tlMasterXbar_monitor_1__GEN_25 ; 
    wire tlMasterXbar_monitor_1__GEN_297 = tlMasterXbar_monitor_1__GEN_67 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_298 = tlMasterXbar_monitor_1__GEN_0 ; 
    wire tlMasterXbar_monitor_1__GEN_299 = tlMasterXbar_monitor_1__GEN_68 ; 
    wire tlMasterXbar_monitor_1__GEN_300 = tlMasterXbar_monitor_1__GEN_69 ; 
    wire tlMasterXbar_monitor_1__GEN_301 = tlMasterXbar_monitor_1__GEN_70 ; 
    wire tlMasterXbar_monitor_1__GEN_302 = tlMasterXbar_monitor_1__GEN_71 ; 
    wire tlMasterXbar_monitor_1__GEN_303 = tlMasterXbar_monitor_1__GEN_72 ; 
    wire tlMasterXbar_monitor_1__GEN_304 = tlMasterXbar_monitor_1__GEN_73 ; 
    wire tlMasterXbar_monitor_1__GEN_305 = tlMasterXbar_monitor_1__GEN_74 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_306 = tlMasterXbar_monitor_1__GEN_13 ; 
    wire tlMasterXbar_monitor_1__GEN_307 = tlMasterXbar_monitor_1__GEN_75 ; 
    wire tlMasterXbar_monitor_1__GEN_308 = tlMasterXbar_monitor_1__GEN_293 ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_309 = tlMasterXbar_monitor_1__GEN_76 ; 
    wire tlMasterXbar_monitor_1__GEN_310 = tlMasterXbar_monitor_1__GEN_77 ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_311 = tlMasterXbar_monitor_1__GEN_37 ; 
    wire tlMasterXbar_monitor_1__GEN_312 = tlMasterXbar_monitor_1__GEN_310 ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_313 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_314 =27'hFFF<< tlMasterXbar_monitor_1_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_315 =~( tlMasterXbar_monitor_1__GEN_314 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_a_first_beats1_decode = tlMasterXbar_monitor_1__GEN_315 [11:3]; 
    wire tlMasterXbar_monitor_1_a_first_beats1_opdata = tlMasterXbar_monitor_1_io_in_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_beats1 = tlMasterXbar_monitor_1_a_first_beats1_opdata  ?  tlMasterXbar_monitor_1_a_first_beats1_decode :9'h0; reg[8:0] tlMasterXbar_monitor_1_a_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_316 ={1'h0, tlMasterXbar_monitor_1_a_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_counter1 = tlMasterXbar_monitor_1__GEN_316 [8:0]; 
    wire tlMasterXbar_monitor_1_a_first = tlMasterXbar_monitor_1_a_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_1_a_first_last = tlMasterXbar_monitor_1_a_first_counter ==9'h1| tlMasterXbar_monitor_1_a_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_1_a_first_done = tlMasterXbar_monitor_1_a_first_last & tlMasterXbar_monitor_1__GEN_313 ; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_count = tlMasterXbar_monitor_1_a_first_beats1 &~ tlMasterXbar_monitor_1_a_first_counter1 ; reg[2:0] tlMasterXbar_monitor_1_opcode ; reg[2:0] tlMasterXbar_monitor_1_param ; reg[3:0] tlMasterXbar_monitor_1_size ; 
    reg tlMasterXbar_monitor_1_source ; reg[31:0] tlMasterXbar_monitor_1_address ; 
    wire tlMasterXbar_monitor_1__GEN_317 = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_318 = tlMasterXbar_monitor_1_io_in_a_bits_opcode == tlMasterXbar_monitor_1_opcode ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_319 = tlMasterXbar_monitor_1_io_in_a_bits_param == tlMasterXbar_monitor_1_param ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_320 = tlMasterXbar_monitor_1_io_in_a_bits_size == tlMasterXbar_monitor_1_size ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_321 = tlMasterXbar_monitor_1_io_in_a_bits_source == tlMasterXbar_monitor_1_source ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_322 = tlMasterXbar_monitor_1_io_in_a_bits_address == tlMasterXbar_monitor_1_address ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_323 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first ; 
    wire tlMasterXbar_monitor_1__GEN_324 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_325 =27'hFFF<< tlMasterXbar_monitor_1_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_326 =~( tlMasterXbar_monitor_1__GEN_325 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1_decode = tlMasterXbar_monitor_1__GEN_326 [11:3]; 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1 = tlMasterXbar_monitor_1_d_first_beats1_opdata  ?  tlMasterXbar_monitor_1_d_first_beats1_decode :9'h0; reg[8:0] tlMasterXbar_monitor_1_d_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_327 ={1'h0, tlMasterXbar_monitor_1_d_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_counter1 = tlMasterXbar_monitor_1__GEN_327 [8:0]; 
    wire tlMasterXbar_monitor_1_d_first = tlMasterXbar_monitor_1_d_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_last = tlMasterXbar_monitor_1_d_first_counter ==9'h1| tlMasterXbar_monitor_1_d_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_done = tlMasterXbar_monitor_1_d_first_last & tlMasterXbar_monitor_1__GEN_324 ; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_count = tlMasterXbar_monitor_1_d_first_beats1 &~ tlMasterXbar_monitor_1_d_first_counter1 ; reg[2:0] tlMasterXbar_monitor_1_opcode_1 ; reg[1:0] tlMasterXbar_monitor_1_param_1 ; reg[3:0] tlMasterXbar_monitor_1_size_1 ; 
    reg tlMasterXbar_monitor_1_source_1 ; reg[1:0] tlMasterXbar_monitor_1_sink ; 
    reg tlMasterXbar_monitor_1_denied ; 
    wire tlMasterXbar_monitor_1__GEN_328 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_329 = tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_opcode_1 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_330 = tlMasterXbar_monitor_1_io_in_d_bits_param == tlMasterXbar_monitor_1_param_1 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_331 = tlMasterXbar_monitor_1_io_in_d_bits_size == tlMasterXbar_monitor_1_size_1 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_332 = tlMasterXbar_monitor_1_io_in_d_bits_source == tlMasterXbar_monitor_1_source_1 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_333 = tlMasterXbar_monitor_1_io_in_d_bits_sink == tlMasterXbar_monitor_1_sink ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_334 = tlMasterXbar_monitor_1_io_in_d_bits_denied == tlMasterXbar_monitor_1_denied ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_335 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first ; 
    reg tlMasterXbar_monitor_1_inflight ; reg[3:0] tlMasterXbar_monitor_1_inflight_opcodes ; reg[7:0] tlMasterXbar_monitor_1_inflight_sizes ; 
    wire tlMasterXbar_monitor_1__GEN_336 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_337 =27'hFFF<< tlMasterXbar_monitor_1_io_in_a_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_338 =~( tlMasterXbar_monitor_1__GEN_337 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_a_first_beats1_decode_1 = tlMasterXbar_monitor_1__GEN_338 [11:3]; 
    wire tlMasterXbar_monitor_1_a_first_beats1_opdata_1 = tlMasterXbar_monitor_1_io_in_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_beats1_1 = tlMasterXbar_monitor_1_a_first_beats1_opdata_1  ?  tlMasterXbar_monitor_1_a_first_beats1_decode_1 :9'h0; reg[8:0] tlMasterXbar_monitor_1_a_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_339 ={1'h0, tlMasterXbar_monitor_1_a_first_counter_1 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_counter1_1 = tlMasterXbar_monitor_1__GEN_339 [8:0]; 
    wire tlMasterXbar_monitor_1_a_first_1 = tlMasterXbar_monitor_1_a_first_counter_1 ==9'h0; 
    wire tlMasterXbar_monitor_1_a_first_last_1 = tlMasterXbar_monitor_1_a_first_counter_1 ==9'h1| tlMasterXbar_monitor_1_a_first_beats1_1 ==9'h0; 
    wire tlMasterXbar_monitor_1_a_first_done_1 = tlMasterXbar_monitor_1_a_first_last_1 & tlMasterXbar_monitor_1__GEN_336 ; 
    wire[8:0] tlMasterXbar_monitor_1_a_first_count_1 = tlMasterXbar_monitor_1_a_first_beats1_1 &~ tlMasterXbar_monitor_1_a_first_counter1_1 ; 
    wire tlMasterXbar_monitor_1__GEN_340 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_341 =27'hFFF<< tlMasterXbar_monitor_1_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_342 =~( tlMasterXbar_monitor_1__GEN_341 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1_decode_1 = tlMasterXbar_monitor_1__GEN_342 [11:3]; 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata_1 = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1_1 = tlMasterXbar_monitor_1_d_first_beats1_opdata_1  ?  tlMasterXbar_monitor_1_d_first_beats1_decode_1 :9'h0; reg[8:0] tlMasterXbar_monitor_1_d_first_counter_1 ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_343 ={1'h0, tlMasterXbar_monitor_1_d_first_counter_1 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_counter1_1 = tlMasterXbar_monitor_1__GEN_343 [8:0]; 
    wire tlMasterXbar_monitor_1_d_first_1 = tlMasterXbar_monitor_1_d_first_counter_1 ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_last_1 = tlMasterXbar_monitor_1_d_first_counter_1 ==9'h1| tlMasterXbar_monitor_1_d_first_beats1_1 ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_done_1 = tlMasterXbar_monitor_1_d_first_last_1 & tlMasterXbar_monitor_1__GEN_340 ; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_count_1 = tlMasterXbar_monitor_1_d_first_beats1_1 &~ tlMasterXbar_monitor_1_d_first_counter1_1 ; 
    wire[15:0] tlMasterXbar_monitor_1__GEN_344 =({12'h0, tlMasterXbar_monitor_1_inflight_opcodes >>({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h2)}&16'hF)>>16'h1; 
    wire[3:0] tlMasterXbar_monitor_1_a_opcode_lookup = tlMasterXbar_monitor_1__GEN_344 [3:0]; 
    wire[15:0] tlMasterXbar_monitor_1__GEN_345 =({8'h0, tlMasterXbar_monitor_1_inflight_sizes >>({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h3)}&16'hFF)>>16'h1; 
    wire[7:0] tlMasterXbar_monitor_1_a_size_lookup = tlMasterXbar_monitor_1__GEN_345 [7:0]; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMap_5 =3'h2; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_0 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_1 =3'h0; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_2 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_3 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_4 =3'h1; 
    wire[2:0] tlMasterXbar_monitor_1_responseMapSecondOption_5 =3'h2; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_346 =2'h1<< tlMasterXbar_monitor_1_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor_1_a_set_wo_ready = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first_1  ?  tlMasterXbar_monitor_1__GEN_346 [0]:1'h0; 
    wire tlMasterXbar_monitor_1__GEN_347 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first_1 ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_348 =2'h1<< tlMasterXbar_monitor_1_io_in_a_bits_source ; 
    wire tlMasterXbar_monitor_1_a_set = tlMasterXbar_monitor_1__GEN_347  ?  tlMasterXbar_monitor_1__GEN_348 [0]:1'h0; 
    wire[3:0] tlMasterXbar_monitor_1_a_opcodes_set_interm = tlMasterXbar_monitor_1__GEN_347  ? {1'h0, tlMasterXbar_monitor_1_io_in_a_bits_opcode }<<4'h1|4'h1:4'h0; 
    wire[4:0] tlMasterXbar_monitor_1_a_sizes_set_interm = tlMasterXbar_monitor_1__GEN_347  ? {1'h0, tlMasterXbar_monitor_1_io_in_a_bits_size }<<5'h1|5'h1:5'h0; 
    wire[18:0] tlMasterXbar_monitor_1__GEN_349 ={15'h0, tlMasterXbar_monitor_1_a_opcodes_set_interm }<<({3'h0, tlMasterXbar_monitor_1_io_in_a_bits_source }<<4'h2); 
    wire[3:0] tlMasterXbar_monitor_1_a_opcodes_set = tlMasterXbar_monitor_1__GEN_347  ?  tlMasterXbar_monitor_1__GEN_349 [3:0]:4'h0; 
    wire[19:0] tlMasterXbar_monitor_1__GEN_350 ={15'h0, tlMasterXbar_monitor_1_a_sizes_set_interm }<<({3'h0, tlMasterXbar_monitor_1_io_in_a_bits_source }<<4'h3); 
    wire[7:0] tlMasterXbar_monitor_1_a_sizes_set = tlMasterXbar_monitor_1__GEN_347  ?  tlMasterXbar_monitor_1__GEN_350 [7:0]:8'h0; 
    wire tlMasterXbar_monitor_1__GEN_351 = tlMasterXbar_monitor_1_inflight >> tlMasterXbar_monitor_1_io_in_a_bits_source ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1_d_release_ack = tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h6; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_352 =2'h1<< tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1_d_clr_wo_ready = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_1 & tlMasterXbar_monitor_1_d_release_ack ==1'h0 ?  tlMasterXbar_monitor_1__GEN_352 [0]:1'h0; 
    wire tlMasterXbar_monitor_1__GEN_353 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_1 & tlMasterXbar_monitor_1_d_release_ack ==1'h0; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_354 =2'h1<< tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1_d_clr = tlMasterXbar_monitor_1__GEN_353  ?  tlMasterXbar_monitor_1__GEN_354 [0]:1'h0; 
    wire[30:0] tlMasterXbar_monitor_1__GEN_355 =31'hF<<({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h2); 
    wire[3:0] tlMasterXbar_monitor_1_d_opcodes_clr = tlMasterXbar_monitor_1__GEN_353  ?  tlMasterXbar_monitor_1__GEN_355 [3:0]:4'h0; 
    wire[30:0] tlMasterXbar_monitor_1__GEN_356 =31'hFF<<({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h3); 
    wire[7:0] tlMasterXbar_monitor_1_d_sizes_clr = tlMasterXbar_monitor_1__GEN_353  ?  tlMasterXbar_monitor_1__GEN_356 [7:0]:8'h0; 
    wire tlMasterXbar_monitor_1__GEN_357 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_1 & tlMasterXbar_monitor_1_d_release_ack ==1'h0; 
    wire tlMasterXbar_monitor_1_same_cycle_resp = tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_a_first_1 & tlMasterXbar_monitor_1_io_in_a_bits_source == tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1__GEN_358 =( tlMasterXbar_monitor_1_inflight >> tlMasterXbar_monitor_1_io_in_d_bits_source | tlMasterXbar_monitor_1_same_cycle_resp )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_359 = tlMasterXbar_monitor_1__GEN_357 & tlMasterXbar_monitor_1_same_cycle_resp ; reg[2:0] tlMasterXbar_monitor_1_casez_tmp ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_6 ;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp  = tlMasterXbar_monitor_1_responseMap_7 ;endcase
         end
  reg[2:0] tlMasterXbar_monitor_1_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_io_in_a_bits_opcode )
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_6 ;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp_0  = tlMasterXbar_monitor_1_responseMapSecondOption_7 ;endcase
         end
    wire tlMasterXbar_monitor_1__GEN_360 =( tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp | tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp_0 )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_361 = tlMasterXbar_monitor_1_io_in_a_bits_size == tlMasterXbar_monitor_1_io_in_d_bits_size ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_362 = tlMasterXbar_monitor_1__GEN_357 &~ tlMasterXbar_monitor_1_same_cycle_resp ; reg[2:0] tlMasterXbar_monitor_1_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_6 ;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp_1  = tlMasterXbar_monitor_1_responseMap_7 ;endcase
         end
  reg[2:0] tlMasterXbar_monitor_1_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( tlMasterXbar_monitor_1_a_opcode_lookup [2:0])
              3 'b000: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_0 ;
              3 'b001: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_1 ;
              3 'b010: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_2 ;
              3 'b011: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_3 ;
              3 'b100: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_4 ;
              3 'b101: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_5 ;
              3 'b110: 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_6 ;
              default : 
                  tlMasterXbar_monitor_1_casez_tmp_2  = tlMasterXbar_monitor_1_responseMapSecondOption_7 ;endcase
         end
    wire tlMasterXbar_monitor_1__GEN_363 =( tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp_1 | tlMasterXbar_monitor_1_io_in_d_bits_opcode == tlMasterXbar_monitor_1_casez_tmp_2 )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_364 ={4'h0, tlMasterXbar_monitor_1_io_in_d_bits_size }== tlMasterXbar_monitor_1_a_size_lookup ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_365 =( tlMasterXbar_monitor_1_io_in_d_ready ==1'h0| tlMasterXbar_monitor_1_io_in_a_ready )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_366 =( tlMasterXbar_monitor_1_a_set_wo_ready != tlMasterXbar_monitor_1_d_clr_wo_ready |(| tlMasterXbar_monitor_1_a_set_wo_ready )==1'h0)==1'h0; reg[31:0] tlMasterXbar_monitor_1_watchdog ;  
    wire tlMasterXbar_monitor_1__GEN_367 =((| tlMasterXbar_monitor_1_inflight )==1'h0| tlMasterXbar_monitor_1__plusarg_reader_out ==32'h0| tlMasterXbar_monitor_1_watchdog < tlMasterXbar_monitor_1__plusarg_reader_out )==1'h0; 
    wire[32:0] tlMasterXbar_monitor_1__GEN_368 ={1'h0, tlMasterXbar_monitor_1_watchdog }+33'h1; 
    wire tlMasterXbar_monitor_1__GEN_369 = tlMasterXbar_monitor_1_io_in_a_ready & tlMasterXbar_monitor_1_io_in_a_valid | tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid ; 
    reg tlMasterXbar_monitor_1_inflight_1 ; reg[3:0] tlMasterXbar_monitor_1_inflight_opcodes_1 ; reg[7:0] tlMasterXbar_monitor_1_inflight_sizes_1 ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_ready = tlMasterXbar_monitor_1__c_first_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_valid = tlMasterXbar_monitor_1__c_first_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_first_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_first_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_first_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_first_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_first_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_first_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_first_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_first_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_first_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_first_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_first_WIRE_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_ready = tlMasterXbar_monitor_1__c_first_WIRE_2_ready ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_valid = tlMasterXbar_monitor_1__c_first_WIRE_2_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_3_bits_opcode = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_first_WIRE_3_bits_param = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_first_WIRE_3_bits_size = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_size ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_source = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_first_WIRE_3_bits_address = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_address ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_first_WIRE_3_bits_data = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_data ; 
    wire tlMasterXbar_monitor_1__c_first_WIRE_3_bits_corrupt = tlMasterXbar_monitor_1__c_first_WIRE_2_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__GEN_370 = tlMasterXbar_monitor_1__c_first_WIRE_3_ready & tlMasterXbar_monitor_1__c_first_WIRE_3_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_371 =27'hFFF<< tlMasterXbar_monitor_1__c_first_WIRE_1_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_372 =~( tlMasterXbar_monitor_1__GEN_371 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_c_first_beats1_decode = tlMasterXbar_monitor_1__GEN_372 [11:3]; 
    wire tlMasterXbar_monitor_1_c_first_beats1_opdata = tlMasterXbar_monitor_1__c_first_WIRE_1_bits_opcode [0]; reg[8:0] tlMasterXbar_monitor_1_c_first_counter ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_373 ={1'h0, tlMasterXbar_monitor_1_c_first_counter }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_c_first_counter1 = tlMasterXbar_monitor_1__GEN_373 [8:0]; 
    wire tlMasterXbar_monitor_1_c_first = tlMasterXbar_monitor_1_c_first_counter ==9'h0; 
    wire tlMasterXbar_monitor_1_c_first_last = tlMasterXbar_monitor_1_c_first_counter ==9'h1| tlMasterXbar_monitor_1_c_first_beats1 ==9'h0; 
    wire tlMasterXbar_monitor_1_c_first_done = tlMasterXbar_monitor_1_c_first_last & tlMasterXbar_monitor_1__GEN_370 ; 
    wire[8:0] tlMasterXbar_monitor_1_c_first_count = tlMasterXbar_monitor_1_c_first_beats1 &~ tlMasterXbar_monitor_1_c_first_counter1 ; 
    wire tlMasterXbar_monitor_1__GEN_374 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid ; 
    wire[26:0] tlMasterXbar_monitor_1__GEN_375 =27'hFFF<< tlMasterXbar_monitor_1_io_in_d_bits_size ; 
    wire[11:0] tlMasterXbar_monitor_1__GEN_376 =~( tlMasterXbar_monitor_1__GEN_375 [11:0]); 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1_decode_2 = tlMasterXbar_monitor_1__GEN_376 [11:3]; 
    wire tlMasterXbar_monitor_1_d_first_beats1_opdata_2 = tlMasterXbar_monitor_1_io_in_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_beats1_2 = tlMasterXbar_monitor_1_d_first_beats1_opdata_2  ?  tlMasterXbar_monitor_1_d_first_beats1_decode_2 :9'h0; reg[8:0] tlMasterXbar_monitor_1_d_first_counter_2 ; 
    wire[9:0] tlMasterXbar_monitor_1__GEN_377 ={1'h0, tlMasterXbar_monitor_1_d_first_counter_2 }-10'h1; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_counter1_2 = tlMasterXbar_monitor_1__GEN_377 [8:0]; 
    wire tlMasterXbar_monitor_1_d_first_2 = tlMasterXbar_monitor_1_d_first_counter_2 ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_last_2 = tlMasterXbar_monitor_1_d_first_counter_2 ==9'h1| tlMasterXbar_monitor_1_d_first_beats1_2 ==9'h0; 
    wire tlMasterXbar_monitor_1_d_first_done_2 = tlMasterXbar_monitor_1_d_first_last_2 & tlMasterXbar_monitor_1__GEN_374 ; 
    wire[8:0] tlMasterXbar_monitor_1_d_first_count_2 = tlMasterXbar_monitor_1_d_first_beats1_2 &~ tlMasterXbar_monitor_1_d_first_counter1_2 ; 
    wire[15:0] tlMasterXbar_monitor_1__GEN_378 =({12'h0, tlMasterXbar_monitor_1_inflight_opcodes_1 >>({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h2)}&16'hF)>>16'h1; 
    wire[3:0] tlMasterXbar_monitor_1_c_opcode_lookup = tlMasterXbar_monitor_1__GEN_378 [3:0]; 
    wire[15:0] tlMasterXbar_monitor_1__GEN_379 =({8'h0, tlMasterXbar_monitor_1_inflight_sizes_1 >>({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h3)}&16'hFF)>>16'h1; 
    wire[7:0] tlMasterXbar_monitor_1_c_size_lookup = tlMasterXbar_monitor_1__GEN_379 [7:0]; 
    wire tlMasterXbar_monitor_1__GEN_380 = tlMasterXbar_monitor_1__GEN_78 ; 
    wire tlMasterXbar_monitor_1__GEN_381 = tlMasterXbar_monitor_1__GEN_79 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_382 = tlMasterXbar_monitor_1__GEN_41 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_383 = tlMasterXbar_monitor_1__GEN_42 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_384 = tlMasterXbar_monitor_1__GEN_26 ; 
    wire tlMasterXbar_monitor_1__GEN_385 = tlMasterXbar_monitor_1__GEN_80 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_386 = tlMasterXbar_monitor_1__GEN_1 ; 
    wire tlMasterXbar_monitor_1__GEN_387 = tlMasterXbar_monitor_1__GEN_81 ; 
    wire tlMasterXbar_monitor_1__GEN_388 = tlMasterXbar_monitor_1__GEN_82 ; 
    wire tlMasterXbar_monitor_1__GEN_389 = tlMasterXbar_monitor_1__GEN_83 ; 
    wire tlMasterXbar_monitor_1__GEN_390 = tlMasterXbar_monitor_1__GEN_84 ; 
    wire tlMasterXbar_monitor_1__GEN_391 = tlMasterXbar_monitor_1__GEN_85 ; 
    wire tlMasterXbar_monitor_1__GEN_392 = tlMasterXbar_monitor_1__GEN_86 ; 
    wire tlMasterXbar_monitor_1__GEN_393 = tlMasterXbar_monitor_1__GEN_87 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_394 = tlMasterXbar_monitor_1__GEN_14 ; 
    wire tlMasterXbar_monitor_1__GEN_395 = tlMasterXbar_monitor_1__GEN_88 ; 
    wire tlMasterXbar_monitor_1__GEN_396 = tlMasterXbar_monitor_1__GEN_89 ; 
    wire tlMasterXbar_monitor_1__GEN_397 = tlMasterXbar_monitor_1__GEN_90 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_398 = tlMasterXbar_monitor_1__GEN_43 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_399 = tlMasterXbar_monitor_1__GEN_44 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_400 = tlMasterXbar_monitor_1__GEN_27 ; 
    wire tlMasterXbar_monitor_1__GEN_401 = tlMasterXbar_monitor_1__GEN_91 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_402 = tlMasterXbar_monitor_1__GEN_2 ; 
    wire tlMasterXbar_monitor_1__GEN_403 = tlMasterXbar_monitor_1__GEN_92 ; 
    wire tlMasterXbar_monitor_1__GEN_404 = tlMasterXbar_monitor_1__GEN_93 ; 
    wire tlMasterXbar_monitor_1__GEN_405 = tlMasterXbar_monitor_1__GEN_94 ; 
    wire tlMasterXbar_monitor_1__GEN_406 = tlMasterXbar_monitor_1__GEN_95 ; 
    wire tlMasterXbar_monitor_1__GEN_407 = tlMasterXbar_monitor_1__GEN_96 ; 
    wire tlMasterXbar_monitor_1__GEN_408 = tlMasterXbar_monitor_1__GEN_97 ; 
    wire tlMasterXbar_monitor_1__GEN_409 = tlMasterXbar_monitor_1__GEN_98 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_410 = tlMasterXbar_monitor_1__GEN_15 ; 
    wire tlMasterXbar_monitor_1__GEN_411 = tlMasterXbar_monitor_1__GEN_99 ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_ready = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_valid = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_bits_corrupt ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_412 =2'h1<< tlMasterXbar_monitor_1__c_set_wo_ready_WIRE_1_bits_source ; 
    wire tlMasterXbar_monitor_1_c_set_wo_ready = tlMasterXbar_monitor_1__GEN_381 & tlMasterXbar_monitor_1_c_first & tlMasterXbar_monitor_1__GEN_398 [2]& tlMasterXbar_monitor_1__GEN_398 [1] ?  tlMasterXbar_monitor_1__GEN_412 [0]:1'h0; 
    wire tlMasterXbar_monitor_1__GEN_413 = tlMasterXbar_monitor_1__GEN_100 ; 
    wire tlMasterXbar_monitor_1__GEN_414 = tlMasterXbar_monitor_1__GEN_101 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_415 = tlMasterXbar_monitor_1__GEN_45 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_416 = tlMasterXbar_monitor_1__GEN_46 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_417 = tlMasterXbar_monitor_1__GEN_28 ; 
    wire tlMasterXbar_monitor_1__GEN_418 = tlMasterXbar_monitor_1__GEN_102 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_419 = tlMasterXbar_monitor_1__GEN_3 ; 
    wire tlMasterXbar_monitor_1__GEN_420 = tlMasterXbar_monitor_1__GEN_103 ; 
    wire tlMasterXbar_monitor_1__GEN_421 = tlMasterXbar_monitor_1__GEN_104 ; 
    wire tlMasterXbar_monitor_1__GEN_422 = tlMasterXbar_monitor_1__GEN_105 ; 
    wire tlMasterXbar_monitor_1__GEN_423 = tlMasterXbar_monitor_1__GEN_106 ; 
    wire tlMasterXbar_monitor_1__GEN_424 = tlMasterXbar_monitor_1__GEN_107 ; 
    wire tlMasterXbar_monitor_1__GEN_425 = tlMasterXbar_monitor_1__GEN_108 ; 
    wire tlMasterXbar_monitor_1__GEN_426 = tlMasterXbar_monitor_1__GEN_109 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_427 = tlMasterXbar_monitor_1__GEN_16 ; 
    wire tlMasterXbar_monitor_1__GEN_428 = tlMasterXbar_monitor_1__GEN_110 ; 
    wire tlMasterXbar_monitor_1__GEN_429 = tlMasterXbar_monitor_1__GEN_111 ; 
    wire tlMasterXbar_monitor_1__GEN_430 = tlMasterXbar_monitor_1__GEN_112 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_431 = tlMasterXbar_monitor_1__GEN_47 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_432 = tlMasterXbar_monitor_1__GEN_48 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_433 = tlMasterXbar_monitor_1__GEN_29 ; 
    wire tlMasterXbar_monitor_1__GEN_434 = tlMasterXbar_monitor_1__GEN_113 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_435 = tlMasterXbar_monitor_1__GEN_4 ; 
    wire tlMasterXbar_monitor_1__GEN_436 = tlMasterXbar_monitor_1__GEN_114 ; 
    wire tlMasterXbar_monitor_1__GEN_437 = tlMasterXbar_monitor_1__GEN_115 ; 
    wire tlMasterXbar_monitor_1__GEN_438 = tlMasterXbar_monitor_1__GEN_116 ; 
    wire tlMasterXbar_monitor_1__GEN_439 = tlMasterXbar_monitor_1__GEN_117 ; 
    wire tlMasterXbar_monitor_1__GEN_440 = tlMasterXbar_monitor_1__GEN_118 ; 
    wire tlMasterXbar_monitor_1__GEN_441 = tlMasterXbar_monitor_1__GEN_119 ; 
    wire tlMasterXbar_monitor_1__GEN_442 = tlMasterXbar_monitor_1__GEN_120 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_443 = tlMasterXbar_monitor_1__GEN_17 ; 
    wire tlMasterXbar_monitor_1__GEN_444 = tlMasterXbar_monitor_1__GEN_121 ; 
    wire tlMasterXbar_monitor_1__GEN_445 = tlMasterXbar_monitor_1__GEN_413 & tlMasterXbar_monitor_1__GEN_414 & tlMasterXbar_monitor_1_c_first & tlMasterXbar_monitor_1__GEN_431 [2]& tlMasterXbar_monitor_1__GEN_431 [1]; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_ready = tlMasterXbar_monitor_1__c_set_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_valid = tlMasterXbar_monitor_1__c_set_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_set_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_set_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_set_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_set_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_set_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_set_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_set_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_set_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_set_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_set_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_set_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_set_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_set_WIRE_bits_corrupt ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_446 =2'h1<< tlMasterXbar_monitor_1__c_set_WIRE_1_bits_source ; 
    wire tlMasterXbar_monitor_1_c_set = tlMasterXbar_monitor_1__GEN_445  ?  tlMasterXbar_monitor_1__GEN_446 [0]:1'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_ready = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_valid = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_bits_corrupt ; 
    wire[3:0] tlMasterXbar_monitor_1_c_opcodes_set_interm = tlMasterXbar_monitor_1__GEN_445  ? {1'h0, tlMasterXbar_monitor_1__c_opcodes_set_interm_WIRE_1_bits_opcode }<<4'h1|4'h1:4'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_ready = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_valid = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_bits_corrupt ; 
    wire[4:0] tlMasterXbar_monitor_1_c_sizes_set_interm = tlMasterXbar_monitor_1__GEN_445  ? {1'h0, tlMasterXbar_monitor_1__c_sizes_set_interm_WIRE_1_bits_size }<<5'h1|5'h1:5'h0; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_ready = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_valid = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_opcodes_set_WIRE_bits_corrupt ; 
    wire[18:0] tlMasterXbar_monitor_1__GEN_447 ={15'h0, tlMasterXbar_monitor_1_c_opcodes_set_interm }<<({3'h0, tlMasterXbar_monitor_1__c_opcodes_set_WIRE_1_bits_source }<<4'h2); 
    wire[3:0] tlMasterXbar_monitor_1_c_opcodes_set = tlMasterXbar_monitor_1__GEN_445  ?  tlMasterXbar_monitor_1__GEN_447 [3:0]:4'h0; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_ready = tlMasterXbar_monitor_1__c_sizes_set_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_valid = tlMasterXbar_monitor_1__c_sizes_set_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_sizes_set_WIRE_bits_corrupt ; 
    wire[19:0] tlMasterXbar_monitor_1__GEN_448 ={15'h0, tlMasterXbar_monitor_1_c_sizes_set_interm }<<({3'h0, tlMasterXbar_monitor_1__c_sizes_set_WIRE_1_bits_source }<<4'h3); 
    wire[7:0] tlMasterXbar_monitor_1_c_sizes_set = tlMasterXbar_monitor_1__GEN_445  ?  tlMasterXbar_monitor_1__GEN_448 [7:0]:8'h0; 
    wire tlMasterXbar_monitor_1__GEN_449 = tlMasterXbar_monitor_1__GEN_122 ; 
    wire tlMasterXbar_monitor_1__GEN_450 = tlMasterXbar_monitor_1__GEN_123 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_451 = tlMasterXbar_monitor_1__GEN_49 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_452 = tlMasterXbar_monitor_1__GEN_50 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_453 = tlMasterXbar_monitor_1__GEN_30 ; 
    wire tlMasterXbar_monitor_1__GEN_454 = tlMasterXbar_monitor_1__GEN_124 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_455 = tlMasterXbar_monitor_1__GEN_5 ; 
    wire tlMasterXbar_monitor_1__GEN_456 = tlMasterXbar_monitor_1__GEN_125 ; 
    wire tlMasterXbar_monitor_1__GEN_457 = tlMasterXbar_monitor_1__GEN_126 ; 
    wire tlMasterXbar_monitor_1__GEN_458 = tlMasterXbar_monitor_1__GEN_127 ; 
    wire tlMasterXbar_monitor_1__GEN_459 = tlMasterXbar_monitor_1__GEN_128 ; 
    wire tlMasterXbar_monitor_1__GEN_460 = tlMasterXbar_monitor_1__GEN_129 ; 
    wire tlMasterXbar_monitor_1__GEN_461 = tlMasterXbar_monitor_1__GEN_130 ; 
    wire tlMasterXbar_monitor_1__GEN_462 = tlMasterXbar_monitor_1__GEN_131 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_463 = tlMasterXbar_monitor_1__GEN_18 ; 
    wire tlMasterXbar_monitor_1__GEN_464 = tlMasterXbar_monitor_1__GEN_132 ; 
    wire tlMasterXbar_monitor_1__GEN_465 = tlMasterXbar_monitor_1_inflight_1 >> tlMasterXbar_monitor_1__GEN_454 ==1'h0==1'h0; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_ready = tlMasterXbar_monitor_1__c_probe_ack_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_valid = tlMasterXbar_monitor_1__c_probe_ack_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_param = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_size = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_source = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_address = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_data = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__c_probe_ack_WIRE_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_ready = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_ready ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_valid = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_opcode = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_param = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_size = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_size ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_source = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_address = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_address ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_data = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_data ; 
    wire tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_corrupt = tlMasterXbar_monitor_1__c_probe_ack_WIRE_2_bits_corrupt ; 
    wire tlMasterXbar_monitor_1_c_probe_ack = tlMasterXbar_monitor_1__c_probe_ack_WIRE_1_bits_opcode ==3'h4| tlMasterXbar_monitor_1__c_probe_ack_WIRE_3_bits_opcode ==3'h5; 
    wire tlMasterXbar_monitor_1_d_release_ack_1 = tlMasterXbar_monitor_1_io_in_d_bits_opcode ==3'h6; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_466 =2'h1<< tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1_d_clr_wo_ready_1 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_2 & tlMasterXbar_monitor_1_d_release_ack_1  ?  tlMasterXbar_monitor_1__GEN_466 [0]:1'h0; 
    wire tlMasterXbar_monitor_1__GEN_467 = tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_2 & tlMasterXbar_monitor_1_d_release_ack_1 ; 
    wire[1:0] tlMasterXbar_monitor_1__GEN_468 =2'h1<< tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1_d_clr_1 = tlMasterXbar_monitor_1__GEN_467  ?  tlMasterXbar_monitor_1__GEN_468 [0]:1'h0; 
    wire[30:0] tlMasterXbar_monitor_1__GEN_469 =31'hF<<({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h2); 
    wire[3:0] tlMasterXbar_monitor_1_d_opcodes_clr_1 = tlMasterXbar_monitor_1__GEN_467  ?  tlMasterXbar_monitor_1__GEN_469 [3:0]:4'h0; 
    wire[30:0] tlMasterXbar_monitor_1__GEN_470 =31'hFF<<({3'h0, tlMasterXbar_monitor_1_io_in_d_bits_source }<<4'h3); 
    wire[7:0] tlMasterXbar_monitor_1_d_sizes_clr_1 = tlMasterXbar_monitor_1__GEN_467  ?  tlMasterXbar_monitor_1__GEN_470 [7:0]:8'h0; 
    wire tlMasterXbar_monitor_1__GEN_471 = tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_2 & tlMasterXbar_monitor_1_d_release_ack_1 ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_ready = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_ready ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_valid = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_opcode = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_param = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_size = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_size ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_source = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_address = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_address ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_data = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_data ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_bits_corrupt = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_ready = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_ready ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_valid = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_opcode = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_param = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_size = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_size ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_source = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_address = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_address ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_data = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_data ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_corrupt = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_2_bits_corrupt ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_ready = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_ready ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_valid = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_valid ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_opcode = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_opcode ; 
    wire[2:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_param = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_param ; 
    wire[3:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_size = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_size ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_source = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_source ; 
    wire[31:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_address = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_address ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_bufferable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_modifiable = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_readalloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_writealloc = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_privileged = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_secure = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_user_amba_prot_fetch = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_data = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_data ; 
    wire tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_corrupt = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_4_bits_corrupt ; 
    wire tlMasterXbar_monitor_1_same_cycle_resp_1 = tlMasterXbar_monitor_1__same_cycle_resp_WIRE_1_valid & tlMasterXbar_monitor_1_c_first & tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_opcode [2]& tlMasterXbar_monitor_1__same_cycle_resp_WIRE_3_bits_opcode [1]& tlMasterXbar_monitor_1__same_cycle_resp_WIRE_5_bits_source == tlMasterXbar_monitor_1_io_in_d_bits_source ; 
    wire tlMasterXbar_monitor_1__GEN_472 =( tlMasterXbar_monitor_1_inflight_1 >> tlMasterXbar_monitor_1_io_in_d_bits_source | tlMasterXbar_monitor_1_same_cycle_resp_1 )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_473 = tlMasterXbar_monitor_1__GEN_133 ; 
    wire tlMasterXbar_monitor_1__GEN_474 = tlMasterXbar_monitor_1__GEN_134 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_475 = tlMasterXbar_monitor_1__GEN_51 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_476 = tlMasterXbar_monitor_1__GEN_52 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_477 = tlMasterXbar_monitor_1__GEN_31 ; 
    wire tlMasterXbar_monitor_1__GEN_478 = tlMasterXbar_monitor_1__GEN_135 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_479 = tlMasterXbar_monitor_1__GEN_6 ; 
    wire tlMasterXbar_monitor_1__GEN_480 = tlMasterXbar_monitor_1__GEN_136 ; 
    wire tlMasterXbar_monitor_1__GEN_481 = tlMasterXbar_monitor_1__GEN_137 ; 
    wire tlMasterXbar_monitor_1__GEN_482 = tlMasterXbar_monitor_1__GEN_138 ; 
    wire tlMasterXbar_monitor_1__GEN_483 = tlMasterXbar_monitor_1__GEN_139 ; 
    wire tlMasterXbar_monitor_1__GEN_484 = tlMasterXbar_monitor_1__GEN_140 ; 
    wire tlMasterXbar_monitor_1__GEN_485 = tlMasterXbar_monitor_1__GEN_141 ; 
    wire tlMasterXbar_monitor_1__GEN_486 = tlMasterXbar_monitor_1__GEN_142 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_487 = tlMasterXbar_monitor_1__GEN_19 ; 
    wire tlMasterXbar_monitor_1__GEN_488 = tlMasterXbar_monitor_1__GEN_143 ; 
    wire tlMasterXbar_monitor_1__GEN_489 = tlMasterXbar_monitor_1_io_in_d_bits_size == tlMasterXbar_monitor_1__GEN_477 ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_490 ={4'h0, tlMasterXbar_monitor_1_io_in_d_bits_size }== tlMasterXbar_monitor_1_c_size_lookup ==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_491 = tlMasterXbar_monitor_1__GEN_144 ; 
    wire tlMasterXbar_monitor_1__GEN_492 = tlMasterXbar_monitor_1__GEN_145 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_493 = tlMasterXbar_monitor_1__GEN_53 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_494 = tlMasterXbar_monitor_1__GEN_54 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_495 = tlMasterXbar_monitor_1__GEN_32 ; 
    wire tlMasterXbar_monitor_1__GEN_496 = tlMasterXbar_monitor_1__GEN_146 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_497 = tlMasterXbar_monitor_1__GEN_7 ; 
    wire tlMasterXbar_monitor_1__GEN_498 = tlMasterXbar_monitor_1__GEN_147 ; 
    wire tlMasterXbar_monitor_1__GEN_499 = tlMasterXbar_monitor_1__GEN_148 ; 
    wire tlMasterXbar_monitor_1__GEN_500 = tlMasterXbar_monitor_1__GEN_149 ; 
    wire tlMasterXbar_monitor_1__GEN_501 = tlMasterXbar_monitor_1__GEN_150 ; 
    wire tlMasterXbar_monitor_1__GEN_502 = tlMasterXbar_monitor_1__GEN_151 ; 
    wire tlMasterXbar_monitor_1__GEN_503 = tlMasterXbar_monitor_1__GEN_152 ; 
    wire tlMasterXbar_monitor_1__GEN_504 = tlMasterXbar_monitor_1__GEN_153 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_505 = tlMasterXbar_monitor_1__GEN_20 ; 
    wire tlMasterXbar_monitor_1__GEN_506 = tlMasterXbar_monitor_1__GEN_154 ; 
    wire tlMasterXbar_monitor_1__GEN_507 = tlMasterXbar_monitor_1__GEN_155 ; 
    wire tlMasterXbar_monitor_1__GEN_508 = tlMasterXbar_monitor_1__GEN_156 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_509 = tlMasterXbar_monitor_1__GEN_55 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_510 = tlMasterXbar_monitor_1__GEN_56 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_511 = tlMasterXbar_monitor_1__GEN_33 ; 
    wire tlMasterXbar_monitor_1__GEN_512 = tlMasterXbar_monitor_1__GEN_157 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_513 = tlMasterXbar_monitor_1__GEN_8 ; 
    wire tlMasterXbar_monitor_1__GEN_514 = tlMasterXbar_monitor_1__GEN_158 ; 
    wire tlMasterXbar_monitor_1__GEN_515 = tlMasterXbar_monitor_1__GEN_159 ; 
    wire tlMasterXbar_monitor_1__GEN_516 = tlMasterXbar_monitor_1__GEN_160 ; 
    wire tlMasterXbar_monitor_1__GEN_517 = tlMasterXbar_monitor_1__GEN_161 ; 
    wire tlMasterXbar_monitor_1__GEN_518 = tlMasterXbar_monitor_1__GEN_162 ; 
    wire tlMasterXbar_monitor_1__GEN_519 = tlMasterXbar_monitor_1__GEN_163 ; 
    wire tlMasterXbar_monitor_1__GEN_520 = tlMasterXbar_monitor_1__GEN_164 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_521 = tlMasterXbar_monitor_1__GEN_21 ; 
    wire tlMasterXbar_monitor_1__GEN_522 = tlMasterXbar_monitor_1__GEN_165 ; 
    wire tlMasterXbar_monitor_1__GEN_523 = tlMasterXbar_monitor_1__GEN_166 ; 
    wire tlMasterXbar_monitor_1__GEN_524 = tlMasterXbar_monitor_1__GEN_167 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_525 = tlMasterXbar_monitor_1__GEN_57 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_526 = tlMasterXbar_monitor_1__GEN_58 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_527 = tlMasterXbar_monitor_1__GEN_34 ; 
    wire tlMasterXbar_monitor_1__GEN_528 = tlMasterXbar_monitor_1__GEN_168 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_529 = tlMasterXbar_monitor_1__GEN_9 ; 
    wire tlMasterXbar_monitor_1__GEN_530 = tlMasterXbar_monitor_1__GEN_169 ; 
    wire tlMasterXbar_monitor_1__GEN_531 = tlMasterXbar_monitor_1__GEN_170 ; 
    wire tlMasterXbar_monitor_1__GEN_532 = tlMasterXbar_monitor_1__GEN_171 ; 
    wire tlMasterXbar_monitor_1__GEN_533 = tlMasterXbar_monitor_1__GEN_172 ; 
    wire tlMasterXbar_monitor_1__GEN_534 = tlMasterXbar_monitor_1__GEN_173 ; 
    wire tlMasterXbar_monitor_1__GEN_535 = tlMasterXbar_monitor_1__GEN_174 ; 
    wire tlMasterXbar_monitor_1__GEN_536 = tlMasterXbar_monitor_1__GEN_175 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_537 = tlMasterXbar_monitor_1__GEN_22 ; 
    wire tlMasterXbar_monitor_1__GEN_538 = tlMasterXbar_monitor_1__GEN_176 ; 
    wire tlMasterXbar_monitor_1__GEN_539 =( tlMasterXbar_monitor_1_io_in_d_ready ==1'h0| tlMasterXbar_monitor_1__GEN_523 )==1'h0; 
    wire tlMasterXbar_monitor_1__GEN_540 = tlMasterXbar_monitor_1_c_set_wo_ready != tlMasterXbar_monitor_1_d_clr_wo_ready_1 ==1'h0; reg[31:0] tlMasterXbar_monitor_1_watchdog_1 ;  
    wire tlMasterXbar_monitor_1__GEN_541 =((| tlMasterXbar_monitor_1_inflight_1 )==1'h0| tlMasterXbar_monitor_1__plusarg_reader_1_out ==32'h0| tlMasterXbar_monitor_1_watchdog_1 < tlMasterXbar_monitor_1__plusarg_reader_1_out )==1'h0; 
  always @( posedge  tlMasterXbar_monitor_1_clock )
         begin 
             if ( tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_188 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel has invalid opcode (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries an address illegal for the specified bank visibility\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_193 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_194 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_195 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_196 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_197 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_198 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_192 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_199 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquireBlock is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_201 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_202 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_203 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_204 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_205 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_206 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_207 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_200 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_208 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel AcquirePerm is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_210 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which master claims it can't emit (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_211 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Get type which slave claims it can't support (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_212 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_213 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_214 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_215 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_209 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_216 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Get is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_217 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_218 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutFull type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_217 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_219 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_217 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_220 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_217 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_221 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_217 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_222 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutFull contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_223 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_224 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries PutPartial type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_223 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_225 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_223 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_226 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_223 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_227 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_223 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_228 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel PutPartial contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_229 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_230 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Arithmetic type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_229 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_231 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_229 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_232 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_229 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_233 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_229 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_234 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_235 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_236 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Logical type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_235 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_237 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_235 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_238 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_235 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_239 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical carries invalid opcode param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_235 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_240 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Logical contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_242 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel carries Hint type which is unexpected using diplomatic parameters (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_243 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_244 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint address not aligned to size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_245 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint carries invalid opcode param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_246 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint contains invalid mask (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_241 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_247 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel Hint is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_248 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel has invalid opcode (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_249 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_250 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_249 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_251 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_249 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_252 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_249 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_253 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_249 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_254 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel ReleaseAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_256 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_257 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid sink ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_258 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_259 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_260 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_255 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_261 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel Grant is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_263 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_264 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_265 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData smaller than a beat (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_266 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries invalid cap param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_267 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData carries toN param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_262 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_268 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel GrantData is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_269 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_270 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_269 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_271 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_269 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_272 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_273 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_274 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_273 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_275 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_273 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_276 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel AccessAckData is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_277 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_278 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_277 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_279 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck carries invalid param (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_277 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_280 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is corrupt (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed: 'D' channel HintAck is denied (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_291 )
                 begin 
                     if (1)$error("Assertion failed: 'B' channel valid and not TL-C (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_308 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel valid and not TL-C (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_312 )
                 begin 
                     if (1)$error("Assertion failed: 'E' channel valid and not TL-C (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_317 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_318 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_317 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_319 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel param changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_317 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_320 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel size changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_317 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_321 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel source changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_317 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_322 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel address changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_329 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel opcode changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_330 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel param changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_331 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel size changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_332 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel source changed within multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_333 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel sink changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_328 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_334 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel denied changed with multibeat operation (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_347 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_351 )
                 begin 
                     if (1)$error("Assertion failed: 'A' channel re-used a source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_357 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_358 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_359 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_360 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_359 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_361 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_362 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_363 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper opcode response (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_362 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_364 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_1 & tlMasterXbar_monitor_1_a_first_1 & tlMasterXbar_monitor_1_io_in_a_valid & tlMasterXbar_monitor_1_io_in_a_bits_source == tlMasterXbar_monitor_1_io_in_d_bits_source & tlMasterXbar_monitor_1_d_release_ack ==1'h0& tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_365 )
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_366 )
                 begin 
                     if (1)$error("Assertion failed: 'A' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_367 )
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_445 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_465 )
                 begin 
                     if (1)$error("Assertion failed: 'C' channel re-used a source ID (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_471 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_472 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel acknowledged for nothing inflight (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_471 & tlMasterXbar_monitor_1_same_cycle_resp_1 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_489 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1__GEN_471 &~ tlMasterXbar_monitor_1_same_cycle_resp_1 & tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_490 )
                 begin 
                     if (1)$error("Assertion failed: 'D' channel contains improper response size (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_io_in_d_valid & tlMasterXbar_monitor_1_d_first_2 & tlMasterXbar_monitor_1_c_first & tlMasterXbar_monitor_1__GEN_492 & tlMasterXbar_monitor_1__GEN_512 == tlMasterXbar_monitor_1_io_in_d_bits_source & tlMasterXbar_monitor_1_d_release_ack_1 & tlMasterXbar_monitor_1_c_probe_ack ==1'h0& tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_539 )
                 begin 
                     if (1)$error("Assertion failed: ready check\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ((| tlMasterXbar_monitor_1_c_set_wo_ready )& tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_540 )
                 begin 
                     if (1)$error("Assertion failed: 'C' and 'D' concurrent, despite minlatency 3 (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:49 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_monitor_1_reset ==1'h0& tlMasterXbar_monitor_1__GEN_541 )
                 begin 
                     if (1)$error("Assertion failed: TileLink timeout expired (connected at src/main/scala/rocket/Frontend.scala:387:21)\n    at Monitor.scala:42 assert(cond, message)\n");
                     if (1)$fatal;
                 end 
         end
    wire[32:0] tlMasterXbar_monitor_1__GEN_542 ={1'h0, tlMasterXbar_monitor_1_watchdog_1 }+33'h1; 
    wire tlMasterXbar_monitor_1__GEN_543 = tlMasterXbar_monitor_1__GEN_177 ; 
    wire tlMasterXbar_monitor_1__GEN_544 = tlMasterXbar_monitor_1__GEN_178 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_545 = tlMasterXbar_monitor_1__GEN_59 ; 
    wire[2:0] tlMasterXbar_monitor_1__GEN_546 = tlMasterXbar_monitor_1__GEN_60 ; 
    wire[3:0] tlMasterXbar_monitor_1__GEN_547 = tlMasterXbar_monitor_1__GEN_35 ; 
    wire tlMasterXbar_monitor_1__GEN_548 = tlMasterXbar_monitor_1__GEN_179 ; 
    wire[31:0] tlMasterXbar_monitor_1__GEN_549 = tlMasterXbar_monitor_1__GEN_10 ; 
    wire tlMasterXbar_monitor_1__GEN_550 = tlMasterXbar_monitor_1__GEN_180 ; 
    wire tlMasterXbar_monitor_1__GEN_551 = tlMasterXbar_monitor_1__GEN_181 ; 
    wire tlMasterXbar_monitor_1__GEN_552 = tlMasterXbar_monitor_1__GEN_182 ; 
    wire tlMasterXbar_monitor_1__GEN_553 = tlMasterXbar_monitor_1__GEN_183 ; 
    wire tlMasterXbar_monitor_1__GEN_554 = tlMasterXbar_monitor_1__GEN_184 ; 
    wire tlMasterXbar_monitor_1__GEN_555 = tlMasterXbar_monitor_1__GEN_185 ; 
    wire tlMasterXbar_monitor_1__GEN_556 = tlMasterXbar_monitor_1__GEN_186 ; 
    wire[63:0] tlMasterXbar_monitor_1__GEN_557 = tlMasterXbar_monitor_1__GEN_23 ; 
    wire tlMasterXbar_monitor_1__GEN_558 = tlMasterXbar_monitor_1__GEN_187 ; 
    wire tlMasterXbar_monitor_1__GEN_559 = tlMasterXbar_monitor_1__GEN_543 & tlMasterXbar_monitor_1__GEN_544 | tlMasterXbar_monitor_1_io_in_d_ready & tlMasterXbar_monitor_1_io_in_d_valid ; 
  always @( posedge  tlMasterXbar_monitor_1_clock )
         begin 
             if ( tlMasterXbar_monitor_1_reset )
                 begin  
                     tlMasterXbar_monitor_1_a_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_1_d_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_1_inflight  <=1'h0; 
                     tlMasterXbar_monitor_1_inflight_opcodes  <=4'h0; 
                     tlMasterXbar_monitor_1_inflight_sizes  <=8'h0; 
                     tlMasterXbar_monitor_1_a_first_counter_1  <=9'h0; 
                     tlMasterXbar_monitor_1_d_first_counter_1  <=9'h0; 
                     tlMasterXbar_monitor_1_watchdog  <=32'h0; 
                     tlMasterXbar_monitor_1_inflight_1  <=1'h0; 
                     tlMasterXbar_monitor_1_inflight_opcodes_1  <=4'h0; 
                     tlMasterXbar_monitor_1_inflight_sizes_1  <=8'h0; 
                     tlMasterXbar_monitor_1_c_first_counter  <=9'h0; 
                     tlMasterXbar_monitor_1_d_first_counter_2  <=9'h0; 
                     tlMasterXbar_monitor_1_watchdog_1  <=32'h0;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_monitor_1__GEN_313 )
                         begin 
                             if ( tlMasterXbar_monitor_1_a_first ) 
                                 tlMasterXbar_monitor_1_a_first_counter  <= tlMasterXbar_monitor_1_a_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_1_a_first_counter  <= tlMasterXbar_monitor_1_a_first_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor_1__GEN_324 )
                         begin 
                             if ( tlMasterXbar_monitor_1_d_first ) 
                                 tlMasterXbar_monitor_1_d_first_counter  <= tlMasterXbar_monitor_1_d_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter  <= tlMasterXbar_monitor_1_d_first_counter1 ;
                         end 
                      else 
                         begin 
                         end  
                     tlMasterXbar_monitor_1_inflight  <=( tlMasterXbar_monitor_1_inflight | tlMasterXbar_monitor_1_a_set )&~ tlMasterXbar_monitor_1_d_clr ; 
                     tlMasterXbar_monitor_1_inflight_opcodes  <=( tlMasterXbar_monitor_1_inflight_opcodes | tlMasterXbar_monitor_1_a_opcodes_set )&~ tlMasterXbar_monitor_1_d_opcodes_clr ; 
                     tlMasterXbar_monitor_1_inflight_sizes  <=( tlMasterXbar_monitor_1_inflight_sizes | tlMasterXbar_monitor_1_a_sizes_set )&~ tlMasterXbar_monitor_1_d_sizes_clr ;
                     if ( tlMasterXbar_monitor_1__GEN_336 )
                         begin 
                             if ( tlMasterXbar_monitor_1_a_first_1 ) 
                                 tlMasterXbar_monitor_1_a_first_counter_1  <= tlMasterXbar_monitor_1_a_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_1_a_first_counter_1  <= tlMasterXbar_monitor_1_a_first_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor_1__GEN_340 )
                         begin 
                             if ( tlMasterXbar_monitor_1_d_first_1 ) 
                                 tlMasterXbar_monitor_1_d_first_counter_1  <= tlMasterXbar_monitor_1_d_first_beats1_1 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter_1  <= tlMasterXbar_monitor_1_d_first_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor_1__GEN_369 ) 
                         tlMasterXbar_monitor_1_watchdog  <=32'h0;
                      else  
                         tlMasterXbar_monitor_1_watchdog  <= tlMasterXbar_monitor_1__GEN_368 [31:0]; 
                     tlMasterXbar_monitor_1_inflight_1  <=( tlMasterXbar_monitor_1_inflight_1 | tlMasterXbar_monitor_1_c_set )&~ tlMasterXbar_monitor_1_d_clr_1 ; 
                     tlMasterXbar_monitor_1_inflight_opcodes_1  <=( tlMasterXbar_monitor_1_inflight_opcodes_1 | tlMasterXbar_monitor_1_c_opcodes_set )&~ tlMasterXbar_monitor_1_d_opcodes_clr_1 ; 
                     tlMasterXbar_monitor_1_inflight_sizes_1  <=( tlMasterXbar_monitor_1_inflight_sizes_1 | tlMasterXbar_monitor_1_c_sizes_set )&~ tlMasterXbar_monitor_1_d_sizes_clr_1 ;
                     if ( tlMasterXbar_monitor_1__GEN_370 )
                         begin 
                             if ( tlMasterXbar_monitor_1_c_first ) 
                                 tlMasterXbar_monitor_1_c_first_counter  <= tlMasterXbar_monitor_1_c_first_beats1 ;
                              else  
                                 tlMasterXbar_monitor_1_c_first_counter  <= tlMasterXbar_monitor_1_c_first_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor_1__GEN_374 )
                         begin 
                             if ( tlMasterXbar_monitor_1_d_first_2 ) 
                                 tlMasterXbar_monitor_1_d_first_counter_2  <= tlMasterXbar_monitor_1_d_first_beats1_2 ;
                              else  
                                 tlMasterXbar_monitor_1_d_first_counter_2  <= tlMasterXbar_monitor_1_d_first_counter1_2 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( tlMasterXbar_monitor_1__GEN_559 ) 
                         tlMasterXbar_monitor_1_watchdog_1  <=32'h0;
                      else  
                         tlMasterXbar_monitor_1_watchdog_1  <= tlMasterXbar_monitor_1__GEN_542 [31:0];
                 end 
         end
  always @( posedge  tlMasterXbar_monitor_1_clock )
         begin 
             if ( tlMasterXbar_monitor_1__GEN_323 )
                 begin  
                     tlMasterXbar_monitor_1_opcode  <= tlMasterXbar_monitor_1_io_in_a_bits_opcode ; 
                     tlMasterXbar_monitor_1_param  <= tlMasterXbar_monitor_1_io_in_a_bits_param ; 
                     tlMasterXbar_monitor_1_size  <= tlMasterXbar_monitor_1_io_in_a_bits_size ; 
                     tlMasterXbar_monitor_1_source  <= tlMasterXbar_monitor_1_io_in_a_bits_source ; 
                     tlMasterXbar_monitor_1_address  <= tlMasterXbar_monitor_1_io_in_a_bits_address ;
                 end 
              else 
                 begin 
                 end 
             if ( tlMasterXbar_monitor_1__GEN_335 )
                 begin  
                     tlMasterXbar_monitor_1_opcode_1  <= tlMasterXbar_monitor_1_io_in_d_bits_opcode ; 
                     tlMasterXbar_monitor_1_param_1  <= tlMasterXbar_monitor_1_io_in_d_bits_param ; 
                     tlMasterXbar_monitor_1_size_1  <= tlMasterXbar_monitor_1_io_in_d_bits_size ; 
                     tlMasterXbar_monitor_1_source_1  <= tlMasterXbar_monitor_1_io_in_d_bits_source ; 
                     tlMasterXbar_monitor_1_sink  <= tlMasterXbar_monitor_1_io_in_d_bits_sink ; 
                     tlMasterXbar_monitor_1_denied  <= tlMasterXbar_monitor_1_io_in_d_bits_denied ;
                 end 
              else 
                 begin 
                 end 
         end
 
    assign tlMasterXbar_monitor_1_clock = tlMasterXbar_clock;
    assign tlMasterXbar_monitor_1_reset = tlMasterXbar_reset;
    assign tlMasterXbar_monitor_1_io_in_a_ready = tlMasterXbar_nodeIn_1_a_ready;
    assign tlMasterXbar_monitor_1_io_in_a_valid = tlMasterXbar_nodeIn_1_a_valid;
    assign tlMasterXbar_monitor_1_io_in_a_bits_opcode = tlMasterXbar_nodeIn_1_a_bits_opcode;
    assign tlMasterXbar_monitor_1_io_in_a_bits_param = tlMasterXbar_nodeIn_1_a_bits_param;
    assign tlMasterXbar_monitor_1_io_in_a_bits_size = tlMasterXbar_nodeIn_1_a_bits_size;
    assign tlMasterXbar_monitor_1_io_in_a_bits_source = tlMasterXbar_nodeIn_1_a_bits_source;
    assign tlMasterXbar_monitor_1_io_in_a_bits_address = tlMasterXbar_nodeIn_1_a_bits_address;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_bufferable = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_modifiable = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_readalloc = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_writealloc = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_privileged = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_privileged;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_secure = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_secure;
    assign tlMasterXbar_monitor_1_io_in_a_bits_user_amba_prot_fetch = tlMasterXbar_nodeIn_1_a_bits_user_amba_prot_fetch;
    assign tlMasterXbar_monitor_1_io_in_a_bits_mask = tlMasterXbar_nodeIn_1_a_bits_mask;
    assign tlMasterXbar_monitor_1_io_in_a_bits_data = tlMasterXbar_nodeIn_1_a_bits_data;
    assign tlMasterXbar_monitor_1_io_in_a_bits_corrupt = tlMasterXbar_nodeIn_1_a_bits_corrupt;
    assign tlMasterXbar_monitor_1_io_in_d_ready = tlMasterXbar_nodeIn_1_d_ready;
    assign tlMasterXbar_monitor_1_io_in_d_valid = tlMasterXbar_nodeIn_1_d_valid;
    assign tlMasterXbar_monitor_1_io_in_d_bits_opcode = tlMasterXbar_nodeIn_1_d_bits_opcode;
    assign tlMasterXbar_monitor_1_io_in_d_bits_param = tlMasterXbar_nodeIn_1_d_bits_param;
    assign tlMasterXbar_monitor_1_io_in_d_bits_size = tlMasterXbar_nodeIn_1_d_bits_size;
    assign tlMasterXbar_monitor_1_io_in_d_bits_source = tlMasterXbar_nodeIn_1_d_bits_source;
    assign tlMasterXbar_monitor_1_io_in_d_bits_sink = tlMasterXbar_nodeIn_1_d_bits_sink;
    assign tlMasterXbar_monitor_1_io_in_d_bits_denied = tlMasterXbar_nodeIn_1_d_bits_denied;
    assign tlMasterXbar_monitor_1_io_in_d_bits_data = tlMasterXbar_nodeIn_1_d_bits_data;
    assign tlMasterXbar_monitor_1_io_in_d_bits_corrupt = tlMasterXbar_nodeIn_1_d_bits_corrupt;
     
    wire tlMasterXbar_out_0_a_ready = tlMasterXbar_nodeOut_a_ready ; 
    wire tlMasterXbar_out_0_a_valid ; 
    wire[2:0] tlMasterXbar_out_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_out_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_a_bits_size ; 
    wire[1:0] tlMasterXbar_out_0_a_bits_source ; 
    wire[31:0] tlMasterXbar_out_0_a_bits_address ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_out_0_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar_out_0_a_bits_mask ; 
    wire[63:0] tlMasterXbar_out_0_a_bits_data ; 
    wire tlMasterXbar_out_0_a_bits_corrupt ; 
    wire tlMasterXbar_out_0_b_ready ; 
    wire tlMasterXbar_out_0_b_valid = tlMasterXbar_nodeOut_b_valid ; 
    wire[2:0] tlMasterXbar_out_0_b_bits_opcode = tlMasterXbar_nodeOut_b_bits_opcode ; 
    wire[1:0] tlMasterXbar_out_0_b_bits_param = tlMasterXbar_nodeOut_b_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_b_bits_size = tlMasterXbar_nodeOut_b_bits_size ; 
    wire[1:0] tlMasterXbar_out_0_b_bits_source = tlMasterXbar_nodeOut_b_bits_source ; 
    wire[31:0] tlMasterXbar_out_0_b_bits_address = tlMasterXbar_nodeOut_b_bits_address ; 
    wire[7:0] tlMasterXbar_out_0_b_bits_mask = tlMasterXbar_nodeOut_b_bits_mask ; 
    wire[63:0] tlMasterXbar_out_0_b_bits_data = tlMasterXbar_nodeOut_b_bits_data ; 
    wire tlMasterXbar_out_0_b_bits_corrupt = tlMasterXbar_nodeOut_b_bits_corrupt ; 
    wire tlMasterXbar_out_0_c_ready = tlMasterXbar_nodeOut_c_ready ; 
    wire tlMasterXbar_out_0_c_valid ; 
    wire[2:0] tlMasterXbar_out_0_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_out_0_c_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_c_bits_size ; 
    wire[1:0] tlMasterXbar_out_0_c_bits_source ; 
    wire[31:0] tlMasterXbar_out_0_c_bits_address ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_out_0_c_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_out_0_c_bits_data ; 
    wire tlMasterXbar_out_0_c_bits_corrupt ; 
    wire tlMasterXbar_out_0_d_ready ; 
    wire tlMasterXbar_out_0_d_valid = tlMasterXbar_nodeOut_d_valid ; 
    wire[2:0] tlMasterXbar_out_0_d_bits_opcode = tlMasterXbar_nodeOut_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_out_0_d_bits_param = tlMasterXbar_nodeOut_d_bits_param ; 
    wire[3:0] tlMasterXbar_out_0_d_bits_size = tlMasterXbar_nodeOut_d_bits_size ; 
    wire[1:0] tlMasterXbar_out_0_d_bits_source = tlMasterXbar_nodeOut_d_bits_source ; 
    wire[1:0] tlMasterXbar_out_0_d_bits_sink = tlMasterXbar_nodeOut_d_bits_sink ; 
    wire tlMasterXbar_out_0_d_bits_denied = tlMasterXbar_nodeOut_d_bits_denied ; 
    wire[63:0] tlMasterXbar_out_0_d_bits_data = tlMasterXbar_nodeOut_d_bits_data ; 
    wire tlMasterXbar_out_0_d_bits_corrupt = tlMasterXbar_nodeOut_d_bits_corrupt ; 
    wire tlMasterXbar_out_0_e_ready = tlMasterXbar_nodeOut_e_ready ; 
    wire tlMasterXbar_out_0_e_valid ; 
    wire[1:0] tlMasterXbar_out_0_e_bits_sink ; 
    wire tlMasterXbar_portsAOI_filtered_0_ready ; 
  assign  tlMasterXbar_nodeIn_a_ready = tlMasterXbar_in_0_a_ready ; 
    wire tlMasterXbar_portsAOI_filtered_0_valid = tlMasterXbar_in_0_a_valid ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_0_bits_opcode = tlMasterXbar_in_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_0_bits_param = tlMasterXbar_in_0_a_bits_param ; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_0_bits_size = tlMasterXbar_in_0_a_bits_size ; 
    wire[1:0] tlMasterXbar_portsAOI_filtered_0_bits_source = tlMasterXbar_in_0_a_bits_source ; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_0_bits_address = tlMasterXbar_in_0_a_bits_address ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_bufferable = tlMasterXbar_in_0_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_modifiable = tlMasterXbar_in_0_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_readalloc = tlMasterXbar_in_0_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_writealloc = tlMasterXbar_in_0_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_privileged = tlMasterXbar_in_0_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_secure = tlMasterXbar_in_0_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_fetch = tlMasterXbar_in_0_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar_portsAOI_filtered_0_bits_mask = tlMasterXbar_in_0_a_bits_mask ; 
    wire[63:0] tlMasterXbar_portsAOI_filtered_0_bits_data = tlMasterXbar_in_0_a_bits_data ; 
    wire tlMasterXbar_portsAOI_filtered_0_bits_corrupt = tlMasterXbar_in_0_a_bits_corrupt ; 
    wire tlMasterXbar_portsBIO_filtered_0_ready = tlMasterXbar_in_0_b_ready ; 
    wire tlMasterXbar_portsBIO_filtered_0_valid ; 
  assign  tlMasterXbar_nodeIn_b_valid = tlMasterXbar_in_0_b_valid ; 
    wire[2:0] tlMasterXbar_portsBIO_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_nodeIn_b_bits_opcode = tlMasterXbar_in_0_b_bits_opcode ; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_0_bits_param ; 
  assign  tlMasterXbar_nodeIn_b_bits_param = tlMasterXbar_in_0_b_bits_param ; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_0_bits_size ; 
  assign  tlMasterXbar_nodeIn_b_bits_size = tlMasterXbar_in_0_b_bits_size ; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_0_bits_source ; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_0_bits_address ; 
  assign  tlMasterXbar_nodeIn_b_bits_address = tlMasterXbar_in_0_b_bits_address ; 
    wire[7:0] tlMasterXbar_portsBIO_filtered_0_bits_mask ; 
  assign  tlMasterXbar_nodeIn_b_bits_mask = tlMasterXbar_in_0_b_bits_mask ; 
    wire[63:0] tlMasterXbar_portsBIO_filtered_0_bits_data ; 
  assign  tlMasterXbar_nodeIn_b_bits_data = tlMasterXbar_in_0_b_bits_data ; 
    wire tlMasterXbar_portsBIO_filtered_0_bits_corrupt ; 
  assign  tlMasterXbar_nodeIn_b_bits_corrupt = tlMasterXbar_in_0_b_bits_corrupt ; 
    wire tlMasterXbar_portsCOI_filtered_0_ready ; 
  assign  tlMasterXbar_nodeIn_c_ready = tlMasterXbar_in_0_c_ready ; 
    wire tlMasterXbar_portsCOI_filtered_0_valid = tlMasterXbar_in_0_c_valid ; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_0_bits_opcode = tlMasterXbar_in_0_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_0_bits_param = tlMasterXbar_in_0_c_bits_param ; 
    wire[3:0] tlMasterXbar_portsCOI_filtered_0_bits_size = tlMasterXbar_in_0_c_bits_size ; 
    wire[1:0] tlMasterXbar_portsCOI_filtered_0_bits_source = tlMasterXbar_in_0_c_bits_source ; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_0_bits_address = tlMasterXbar_in_0_c_bits_address ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_bufferable = tlMasterXbar_in_0_c_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_modifiable = tlMasterXbar_in_0_c_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_readalloc = tlMasterXbar_in_0_c_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_writealloc = tlMasterXbar_in_0_c_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_privileged = tlMasterXbar_in_0_c_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_secure = tlMasterXbar_in_0_c_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_fetch = tlMasterXbar_in_0_c_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_portsCOI_filtered_0_bits_data = tlMasterXbar_in_0_c_bits_data ; 
    wire tlMasterXbar_portsCOI_filtered_0_bits_corrupt = tlMasterXbar_in_0_c_bits_corrupt ; 
    wire tlMasterXbar_portsDIO_filtered_0_ready = tlMasterXbar_in_0_d_ready ; 
    wire tlMasterXbar_portsDIO_filtered_0_valid ; 
  assign  tlMasterXbar_nodeIn_d_valid = tlMasterXbar_in_0_d_valid ; 
    wire[2:0] tlMasterXbar_portsDIO_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_nodeIn_d_bits_opcode = tlMasterXbar_in_0_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_0_bits_param ; 
  assign  tlMasterXbar_nodeIn_d_bits_param = tlMasterXbar_in_0_d_bits_param ; 
    wire[3:0] tlMasterXbar_portsDIO_filtered_0_bits_size ; 
  assign  tlMasterXbar_nodeIn_d_bits_size = tlMasterXbar_in_0_d_bits_size ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_0_bits_source ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_0_bits_sink ; 
  assign  tlMasterXbar_nodeIn_d_bits_sink = tlMasterXbar_in_0_d_bits_sink ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_denied ; 
  assign  tlMasterXbar_nodeIn_d_bits_denied = tlMasterXbar_in_0_d_bits_denied ; 
    wire[63:0] tlMasterXbar_portsDIO_filtered_0_bits_data ; 
  assign  tlMasterXbar_nodeIn_d_bits_data = tlMasterXbar_in_0_d_bits_data ; 
    wire tlMasterXbar_portsDIO_filtered_0_bits_corrupt ; 
  assign  tlMasterXbar_nodeIn_d_bits_corrupt = tlMasterXbar_in_0_d_bits_corrupt ; 
    wire tlMasterXbar_portsEOI_filtered_0_ready ; 
  assign  tlMasterXbar_nodeIn_e_ready = tlMasterXbar_in_0_e_ready ; 
    wire tlMasterXbar_portsEOI_filtered_0_valid = tlMasterXbar_in_0_e_valid ; 
    wire[1:0] tlMasterXbar_requestEIO_uncommonBits = tlMasterXbar_in_0_e_bits_sink ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_ready ; 
    wire[1:0] tlMasterXbar_portsEOI_filtered_0_bits_sink = tlMasterXbar_in_0_e_bits_sink ; 
  assign  tlMasterXbar_nodeIn_1_a_ready = tlMasterXbar_in_1_a_ready ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_valid = tlMasterXbar_in_1_a_valid ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_1_0_bits_opcode = tlMasterXbar_in_1_a_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsAOI_filtered_1_0_bits_param = tlMasterXbar_in_1_a_bits_param ; 
    wire[3:0] tlMasterXbar_portsAOI_filtered_1_0_bits_size = tlMasterXbar_in_1_a_bits_size ; 
    wire[1:0] tlMasterXbar_portsAOI_filtered_1_0_bits_source = tlMasterXbar_in_1_a_bits_source ; 
    wire[31:0] tlMasterXbar_portsAOI_filtered_1_0_bits_address = tlMasterXbar_in_1_a_bits_address ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_bufferable = tlMasterXbar_in_1_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_modifiable = tlMasterXbar_in_1_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_readalloc = tlMasterXbar_in_1_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_writealloc = tlMasterXbar_in_1_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_privileged = tlMasterXbar_in_1_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_secure = tlMasterXbar_in_1_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_fetch = tlMasterXbar_in_1_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar_portsAOI_filtered_1_0_bits_mask = tlMasterXbar_in_1_a_bits_mask ; 
    wire[63:0] tlMasterXbar_portsAOI_filtered_1_0_bits_data = tlMasterXbar_in_1_a_bits_data ; 
    wire tlMasterXbar_portsAOI_filtered_1_0_bits_corrupt = tlMasterXbar_in_1_a_bits_corrupt ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_valid = tlMasterXbar_in_1_c_valid ; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_1_0_bits_opcode = tlMasterXbar_in_1_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsCOI_filtered_1_0_bits_param = tlMasterXbar_in_1_c_bits_param ; 
    wire[3:0] tlMasterXbar_portsCOI_filtered_1_0_bits_size = tlMasterXbar_in_1_c_bits_size ; 
    wire[1:0] tlMasterXbar_portsCOI_filtered_1_0_bits_source = tlMasterXbar_in_1_c_bits_source ; 
    wire[31:0] tlMasterXbar_portsCOI_filtered_1_0_bits_address = tlMasterXbar_in_1_c_bits_address ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_bufferable = tlMasterXbar_in_1_c_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_modifiable = tlMasterXbar_in_1_c_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_readalloc = tlMasterXbar_in_1_c_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_writealloc = tlMasterXbar_in_1_c_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_privileged = tlMasterXbar_in_1_c_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_secure = tlMasterXbar_in_1_c_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_user_amba_prot_fetch = tlMasterXbar_in_1_c_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_portsCOI_filtered_1_0_bits_data = tlMasterXbar_in_1_c_bits_data ; 
    wire tlMasterXbar_portsCOI_filtered_1_0_bits_corrupt = tlMasterXbar_in_1_c_bits_corrupt ; 
    wire tlMasterXbar_portsDIO_filtered_1_ready = tlMasterXbar_in_1_d_ready ; 
    wire tlMasterXbar_portsDIO_filtered_1_valid ; 
  assign  tlMasterXbar_nodeIn_1_d_valid = tlMasterXbar_in_1_d_valid ; 
    wire[2:0] tlMasterXbar_portsDIO_filtered_1_bits_opcode ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_opcode = tlMasterXbar_in_1_d_bits_opcode ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_1_bits_param ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_param = tlMasterXbar_in_1_d_bits_param ; 
    wire[3:0] tlMasterXbar_portsDIO_filtered_1_bits_size ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_size = tlMasterXbar_in_1_d_bits_size ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_1_bits_source ; 
    wire[1:0] tlMasterXbar_portsDIO_filtered_1_bits_sink ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_sink = tlMasterXbar_in_1_d_bits_sink ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_denied ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_denied = tlMasterXbar_in_1_d_bits_denied ; 
    wire[63:0] tlMasterXbar_portsDIO_filtered_1_bits_data ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_data = tlMasterXbar_in_1_d_bits_data ; 
    wire tlMasterXbar_portsDIO_filtered_1_bits_corrupt ; 
  assign  tlMasterXbar_nodeIn_1_d_bits_corrupt = tlMasterXbar_in_1_d_bits_corrupt ; 
    wire tlMasterXbar_portsEOI_filtered_1_0_valid = tlMasterXbar_in_1_e_valid ; 
    wire[1:0] tlMasterXbar_requestEIO_uncommonBits_1 = tlMasterXbar_in_1_e_bits_sink ; 
    wire[1:0] tlMasterXbar_portsEOI_filtered_1_0_bits_sink = tlMasterXbar_in_1_e_bits_sink ; 
  assign  tlMasterXbar_in_0_a_bits_source ={1'h0, tlMasterXbar_nodeIn_a_bits_source }; 
    wire[1:0] tlMasterXbar_in_0_b_bits_source ; 
  assign  tlMasterXbar_nodeIn_b_bits_source = tlMasterXbar_in_0_b_bits_source [0]; 
  assign  tlMasterXbar_in_0_c_bits_source ={1'h0, tlMasterXbar_nodeIn_c_bits_source }; 
    wire[1:0] tlMasterXbar_in_0_d_bits_source ; 
  assign  tlMasterXbar_nodeIn_d_bits_source = tlMasterXbar_in_0_d_bits_source [0]; 
  assign  tlMasterXbar_in_1_a_bits_source ={1'h0, tlMasterXbar_nodeIn_1_a_bits_source }|2'h2; 
    wire tlMasterXbar__GEN_89 = tlMasterXbar__GEN_45 ; 
    wire[2:0] tlMasterXbar__GEN_90 = tlMasterXbar__GEN_3 ; 
    wire[1:0] tlMasterXbar__GEN_91 = tlMasterXbar__GEN_12 ; 
    wire[3:0] tlMasterXbar__GEN_92 = tlMasterXbar__GEN_18 ; 
    wire tlMasterXbar__GEN_93 = tlMasterXbar__GEN_47 ; 
    wire[31:0] tlMasterXbar__GEN_94 = tlMasterXbar__GEN_24 ; 
    wire[7:0] tlMasterXbar__GEN_95 = tlMasterXbar__GEN_30 ; 
    wire[63:0] tlMasterXbar__GEN_96 = tlMasterXbar__GEN_33 ; 
    wire tlMasterXbar__GEN_97 = tlMasterXbar__GEN_48 ; 
    wire tlMasterXbar__GEN_98 = tlMasterXbar__GEN_73 ; 
    wire[2:0] tlMasterXbar__GEN_99 = tlMasterXbar__GEN_8 ; 
    wire[2:0] tlMasterXbar__GEN_100 = tlMasterXbar__GEN_9 ; 
    wire[3:0] tlMasterXbar__GEN_101 = tlMasterXbar__GEN_21 ; 
    wire tlMasterXbar__GEN_102 = tlMasterXbar__GEN_74 ; 
    wire[31:0] tlMasterXbar__GEN_103 = tlMasterXbar__GEN_27 ; 
    wire tlMasterXbar__GEN_104 = tlMasterXbar__GEN_75 ; 
    wire tlMasterXbar__GEN_105 = tlMasterXbar__GEN_76 ; 
    wire tlMasterXbar__GEN_106 = tlMasterXbar__GEN_77 ; 
    wire tlMasterXbar__GEN_107 = tlMasterXbar__GEN_78 ; 
    wire tlMasterXbar__GEN_108 = tlMasterXbar__GEN_79 ; 
    wire tlMasterXbar__GEN_109 = tlMasterXbar__GEN_80 ; 
    wire tlMasterXbar__GEN_110 = tlMasterXbar__GEN_81 ; 
    wire[63:0] tlMasterXbar__GEN_111 = tlMasterXbar__GEN_36 ; 
    wire tlMasterXbar__GEN_112 = tlMasterXbar__GEN_82 ; 
    wire[1:0] tlMasterXbar_in_1_d_bits_source ; 
    wire tlMasterXbar__GEN_113 = tlMasterXbar__GEN_88 ; 
    wire[1:0] tlMasterXbar__GEN_114 = tlMasterXbar__GEN_15 ; 
    wire tlMasterXbar_nodeOut_a_valid = tlMasterXbar_out_0_a_valid ; 
    wire[2:0] tlMasterXbar__out_0_a_bits_WIRE_opcode ; 
    wire[2:0] tlMasterXbar_nodeOut_a_bits_opcode = tlMasterXbar_out_0_a_bits_opcode ; 
    wire[2:0] tlMasterXbar__out_0_a_bits_WIRE_param ; 
    wire[2:0] tlMasterXbar_nodeOut_a_bits_param = tlMasterXbar_out_0_a_bits_param ; 
    wire[3:0] tlMasterXbar__out_0_a_bits_WIRE_size ; 
    wire[3:0] tlMasterXbar_nodeOut_a_bits_size = tlMasterXbar_out_0_a_bits_size ; 
    wire[1:0] tlMasterXbar__out_0_a_bits_WIRE_source ; 
    wire[1:0] tlMasterXbar_nodeOut_a_bits_source = tlMasterXbar_out_0_a_bits_source ; 
    wire[31:0] tlMasterXbar__out_0_a_bits_WIRE_address ; 
    wire[31:0] tlMasterXbar_nodeOut_a_bits_address = tlMasterXbar_out_0_a_bits_address ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_bufferable = tlMasterXbar_out_0_a_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_modifiable = tlMasterXbar_out_0_a_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_readalloc = tlMasterXbar_out_0_a_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_writealloc = tlMasterXbar_out_0_a_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_privileged ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_privileged = tlMasterXbar_out_0_a_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_secure ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_secure = tlMasterXbar_out_0_a_bits_user_amba_prot_secure ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_fetch ; 
    wire tlMasterXbar_nodeOut_a_bits_user_amba_prot_fetch = tlMasterXbar_out_0_a_bits_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar__out_0_a_bits_WIRE_mask ; 
    wire[7:0] tlMasterXbar_nodeOut_a_bits_mask = tlMasterXbar_out_0_a_bits_mask ; 
    wire[63:0] tlMasterXbar__out_0_a_bits_WIRE_data ; 
    wire[63:0] tlMasterXbar_nodeOut_a_bits_data = tlMasterXbar_out_0_a_bits_data ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_corrupt ; 
    wire tlMasterXbar_nodeOut_a_bits_corrupt = tlMasterXbar_out_0_a_bits_corrupt ; 
    wire tlMasterXbar__portsBIO_out_0_b_ready_WIRE ; 
    wire tlMasterXbar_nodeOut_b_ready = tlMasterXbar_out_0_b_ready ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_opcode = tlMasterXbar_out_0_b_bits_opcode ; 
    wire[2:0] tlMasterXbar_portsBIO_filtered_1_bits_opcode = tlMasterXbar_out_0_b_bits_opcode ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_param = tlMasterXbar_out_0_b_bits_param ; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_1_bits_param = tlMasterXbar_out_0_b_bits_param ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_size = tlMasterXbar_out_0_b_bits_size ; 
    wire[3:0] tlMasterXbar_portsBIO_filtered_1_bits_size = tlMasterXbar_out_0_b_bits_size ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_source = tlMasterXbar_out_0_b_bits_source ; 
    wire[1:0] tlMasterXbar_portsBIO_filtered_1_bits_source = tlMasterXbar_out_0_b_bits_source ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_address = tlMasterXbar_out_0_b_bits_address ; 
    wire[31:0] tlMasterXbar_portsBIO_filtered_1_bits_address = tlMasterXbar_out_0_b_bits_address ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_mask = tlMasterXbar_out_0_b_bits_mask ; 
    wire[7:0] tlMasterXbar_portsBIO_filtered_1_bits_mask = tlMasterXbar_out_0_b_bits_mask ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_data = tlMasterXbar_out_0_b_bits_data ; 
    wire[63:0] tlMasterXbar_portsBIO_filtered_1_bits_data = tlMasterXbar_out_0_b_bits_data ; 
  assign  tlMasterXbar_portsBIO_filtered_0_bits_corrupt = tlMasterXbar_out_0_b_bits_corrupt ; 
    wire tlMasterXbar_portsBIO_filtered_1_bits_corrupt = tlMasterXbar_out_0_b_bits_corrupt ; 
  assign  tlMasterXbar_portsCOI_filtered_0_ready = tlMasterXbar_out_0_c_ready ; 
    wire tlMasterXbar_nodeOut_c_valid = tlMasterXbar_out_0_c_valid ; 
    wire[2:0] tlMasterXbar_nodeOut_c_bits_opcode = tlMasterXbar_out_0_c_bits_opcode ; 
    wire[2:0] tlMasterXbar_nodeOut_c_bits_param = tlMasterXbar_out_0_c_bits_param ; 
    wire[3:0] tlMasterXbar_nodeOut_c_bits_size = tlMasterXbar_out_0_c_bits_size ; 
    wire[1:0] tlMasterXbar_nodeOut_c_bits_source = tlMasterXbar_out_0_c_bits_source ; 
    wire[31:0] tlMasterXbar_nodeOut_c_bits_address = tlMasterXbar_out_0_c_bits_address ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_bufferable = tlMasterXbar_out_0_c_bits_user_amba_prot_bufferable ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_modifiable = tlMasterXbar_out_0_c_bits_user_amba_prot_modifiable ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_readalloc = tlMasterXbar_out_0_c_bits_user_amba_prot_readalloc ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_writealloc = tlMasterXbar_out_0_c_bits_user_amba_prot_writealloc ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_privileged = tlMasterXbar_out_0_c_bits_user_amba_prot_privileged ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_secure = tlMasterXbar_out_0_c_bits_user_amba_prot_secure ; 
    wire tlMasterXbar_nodeOut_c_bits_user_amba_prot_fetch = tlMasterXbar_out_0_c_bits_user_amba_prot_fetch ; 
    wire[63:0] tlMasterXbar_nodeOut_c_bits_data = tlMasterXbar_out_0_c_bits_data ; 
    wire tlMasterXbar_nodeOut_c_bits_corrupt = tlMasterXbar_out_0_c_bits_corrupt ; 
    wire tlMasterXbar__portsDIO_out_0_d_ready_WIRE ; 
    wire tlMasterXbar_nodeOut_d_ready = tlMasterXbar_out_0_d_ready ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_opcode = tlMasterXbar_out_0_d_bits_opcode ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_opcode = tlMasterXbar_out_0_d_bits_opcode ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_param = tlMasterXbar_out_0_d_bits_param ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_param = tlMasterXbar_out_0_d_bits_param ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_size = tlMasterXbar_out_0_d_bits_size ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_size = tlMasterXbar_out_0_d_bits_size ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_source = tlMasterXbar_out_0_d_bits_source ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_source = tlMasterXbar_out_0_d_bits_source ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_sink = tlMasterXbar_out_0_d_bits_sink ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_sink = tlMasterXbar_out_0_d_bits_sink ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_denied = tlMasterXbar_out_0_d_bits_denied ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_denied = tlMasterXbar_out_0_d_bits_denied ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_data = tlMasterXbar_out_0_d_bits_data ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_data = tlMasterXbar_out_0_d_bits_data ; 
  assign  tlMasterXbar_portsDIO_filtered_0_bits_corrupt = tlMasterXbar_out_0_d_bits_corrupt ; 
  assign  tlMasterXbar_portsDIO_filtered_1_bits_corrupt = tlMasterXbar_out_0_d_bits_corrupt ; 
  assign  tlMasterXbar_portsEOI_filtered_0_ready = tlMasterXbar_out_0_e_ready ; 
    wire tlMasterXbar_nodeOut_e_valid = tlMasterXbar_out_0_e_valid ; 
    wire[1:0] tlMasterXbar_nodeOut_e_bits_sink = tlMasterXbar_out_0_e_bits_sink ; 
    wire tlMasterXbar_requestBOI_uncommonBits = tlMasterXbar_out_0_b_bits_source [0]; 
    wire tlMasterXbar_requestBOI_0_0 = tlMasterXbar_out_0_b_bits_source [1]==1'h0&1'h0<= tlMasterXbar_requestBOI_uncommonBits & tlMasterXbar_requestBOI_uncommonBits <=1'h1; 
    wire tlMasterXbar_requestBOI_0_1 = tlMasterXbar_out_0_b_bits_source ==2'h2; 
    wire tlMasterXbar_requestDOI_uncommonBits = tlMasterXbar_out_0_d_bits_source [0]; 
    wire tlMasterXbar_requestDOI_0_0 = tlMasterXbar_out_0_d_bits_source [1]==1'h0&1'h0<= tlMasterXbar_requestDOI_uncommonBits & tlMasterXbar_requestDOI_uncommonBits <=1'h1; 
    wire tlMasterXbar_requestDOI_0_1 = tlMasterXbar_out_0_d_bits_source ==2'h2; 
    wire tlMasterXbar_requestEIO_0_0 =2'h0<= tlMasterXbar_requestEIO_uncommonBits &1'h1& tlMasterXbar_requestEIO_uncommonBits <=2'h3; 
    wire tlMasterXbar_requestEIO_1_0 =2'h0<= tlMasterXbar_requestEIO_uncommonBits_1 &1'h1& tlMasterXbar_requestEIO_uncommonBits_1 <=2'h3; 
    wire[26:0] tlMasterXbar__GEN_115 =27'hFFF<< tlMasterXbar_in_0_a_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_116 =~( tlMasterXbar__GEN_115 [11:0]); 
    wire[8:0] tlMasterXbar_beatsAI_decode = tlMasterXbar__GEN_116 [11:3]; 
    wire tlMasterXbar_beatsAI_opdata = tlMasterXbar_in_0_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_beatsAI_0 = tlMasterXbar_beatsAI_opdata  ?  tlMasterXbar_beatsAI_decode :9'h0; 
    wire[26:0] tlMasterXbar__GEN_117 =27'hFFF<< tlMasterXbar_in_1_a_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_118 =~( tlMasterXbar__GEN_117 [11:0]); 
    wire[8:0] tlMasterXbar_beatsAI_decode_1 = tlMasterXbar__GEN_118 [11:3]; 
    wire tlMasterXbar_beatsAI_opdata_1 = tlMasterXbar_in_1_a_bits_opcode [2]==1'h0; 
    wire[8:0] tlMasterXbar_beatsAI_1 = tlMasterXbar_beatsAI_opdata_1  ?  tlMasterXbar_beatsAI_decode_1 :9'h0; 
    wire[26:0] tlMasterXbar__GEN_119 =27'hFFF<< tlMasterXbar_out_0_b_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_120 =~( tlMasterXbar__GEN_119 [11:0]); 
    wire[8:0] tlMasterXbar_beatsBO_decode = tlMasterXbar__GEN_120 [11:3]; 
    wire tlMasterXbar_beatsBO_opdata = tlMasterXbar_out_0_b_bits_opcode [2]==1'h0; 
    wire[26:0] tlMasterXbar__GEN_121 =27'hFFF<< tlMasterXbar_in_0_c_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_122 =~( tlMasterXbar__GEN_121 [11:0]); 
    wire[8:0] tlMasterXbar_beatsCI_decode = tlMasterXbar__GEN_122 [11:3]; 
    wire tlMasterXbar_beatsCI_opdata = tlMasterXbar_in_0_c_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_beatsCI_0 = tlMasterXbar_beatsCI_opdata  ?  tlMasterXbar_beatsCI_decode :9'h0; 
    wire[26:0] tlMasterXbar__GEN_123 =27'hFFF<< tlMasterXbar_in_1_c_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_124 =~( tlMasterXbar__GEN_123 [11:0]); 
    wire[8:0] tlMasterXbar_beatsCI_decode_1 = tlMasterXbar__GEN_124 [11:3]; 
    wire tlMasterXbar_beatsCI_opdata_1 = tlMasterXbar_in_1_c_bits_opcode [0]; 
    wire[26:0] tlMasterXbar__GEN_125 =27'hFFF<< tlMasterXbar_out_0_d_bits_size ; 
    wire[11:0] tlMasterXbar__GEN_126 =~( tlMasterXbar__GEN_125 [11:0]); 
    wire[8:0] tlMasterXbar_beatsDO_decode = tlMasterXbar__GEN_126 [11:3]; 
    wire tlMasterXbar_beatsDO_opdata = tlMasterXbar_out_0_d_bits_opcode [0]; 
    wire[8:0] tlMasterXbar_beatsDO_0 = tlMasterXbar_beatsDO_opdata  ?  tlMasterXbar_beatsDO_decode :9'h0; 
  assign  tlMasterXbar_in_0_a_ready = tlMasterXbar_portsAOI_filtered_0_ready ; 
  assign  tlMasterXbar_in_1_a_ready = tlMasterXbar_portsAOI_filtered_1_0_ready ; 
  assign  tlMasterXbar_in_0_b_valid = tlMasterXbar_portsBIO_filtered_0_valid ; 
  assign  tlMasterXbar_in_0_b_bits_opcode = tlMasterXbar_portsBIO_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_in_0_b_bits_param = tlMasterXbar_portsBIO_filtered_0_bits_param ; 
  assign  tlMasterXbar_in_0_b_bits_size = tlMasterXbar_portsBIO_filtered_0_bits_size ; 
  assign  tlMasterXbar_in_0_b_bits_source = tlMasterXbar_portsBIO_filtered_0_bits_source ; 
  assign  tlMasterXbar_in_0_b_bits_address = tlMasterXbar_portsBIO_filtered_0_bits_address ; 
  assign  tlMasterXbar_in_0_b_bits_mask = tlMasterXbar_portsBIO_filtered_0_bits_mask ; 
  assign  tlMasterXbar_in_0_b_bits_data = tlMasterXbar_portsBIO_filtered_0_bits_data ; 
  assign  tlMasterXbar_in_0_b_bits_corrupt = tlMasterXbar_portsBIO_filtered_0_bits_corrupt ; 
  assign  tlMasterXbar_portsBIO_filtered_0_valid = tlMasterXbar_out_0_b_valid & tlMasterXbar_requestBOI_0_0 ; 
    wire tlMasterXbar_portsBIO_filtered_1_valid = tlMasterXbar_out_0_b_valid & tlMasterXbar_requestBOI_0_1 ; 
  assign  tlMasterXbar__portsBIO_out_0_b_ready_WIRE =( tlMasterXbar_requestBOI_0_0  ?  tlMasterXbar_portsBIO_filtered_0_ready :1'h0)|( tlMasterXbar_requestBOI_0_1  ?  tlMasterXbar_portsBIO_filtered_1_ready :1'h0); 
  assign  tlMasterXbar_out_0_b_ready = tlMasterXbar__portsBIO_out_0_b_ready_WIRE ; 
  assign  tlMasterXbar_in_0_c_ready = tlMasterXbar_portsCOI_filtered_0_ready ; 
  assign  tlMasterXbar_out_0_c_valid = tlMasterXbar_portsCOI_filtered_0_valid ; 
  assign  tlMasterXbar_out_0_c_bits_opcode = tlMasterXbar_portsCOI_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_out_0_c_bits_param = tlMasterXbar_portsCOI_filtered_0_bits_param ; 
  assign  tlMasterXbar_out_0_c_bits_size = tlMasterXbar_portsCOI_filtered_0_bits_size ; 
  assign  tlMasterXbar_out_0_c_bits_source = tlMasterXbar_portsCOI_filtered_0_bits_source ; 
  assign  tlMasterXbar_out_0_c_bits_address = tlMasterXbar_portsCOI_filtered_0_bits_address ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_bufferable = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_bufferable ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_modifiable = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_modifiable ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_readalloc = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_readalloc ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_writealloc = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_writealloc ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_privileged = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_privileged ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_secure = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_secure ; 
  assign  tlMasterXbar_out_0_c_bits_user_amba_prot_fetch = tlMasterXbar_portsCOI_filtered_0_bits_user_amba_prot_fetch ; 
  assign  tlMasterXbar_out_0_c_bits_data = tlMasterXbar_portsCOI_filtered_0_bits_data ; 
  assign  tlMasterXbar_out_0_c_bits_corrupt = tlMasterXbar_portsCOI_filtered_0_bits_corrupt ; 
    wire tlMasterXbar_in_1_c_ready = tlMasterXbar_portsCOI_filtered_1_0_ready ; 
  assign  tlMasterXbar_in_0_d_valid = tlMasterXbar_portsDIO_filtered_0_valid ; 
  assign  tlMasterXbar_in_0_d_bits_opcode = tlMasterXbar_portsDIO_filtered_0_bits_opcode ; 
  assign  tlMasterXbar_in_0_d_bits_param = tlMasterXbar_portsDIO_filtered_0_bits_param ; 
  assign  tlMasterXbar_in_0_d_bits_size = tlMasterXbar_portsDIO_filtered_0_bits_size ; 
  assign  tlMasterXbar_in_0_d_bits_source = tlMasterXbar_portsDIO_filtered_0_bits_source ; 
  assign  tlMasterXbar_in_0_d_bits_sink = tlMasterXbar_portsDIO_filtered_0_bits_sink ; 
  assign  tlMasterXbar_in_0_d_bits_denied = tlMasterXbar_portsDIO_filtered_0_bits_denied ; 
  assign  tlMasterXbar_in_0_d_bits_data = tlMasterXbar_portsDIO_filtered_0_bits_data ; 
  assign  tlMasterXbar_in_0_d_bits_corrupt = tlMasterXbar_portsDIO_filtered_0_bits_corrupt ; 
  assign  tlMasterXbar_in_1_d_valid = tlMasterXbar_portsDIO_filtered_1_valid ; 
  assign  tlMasterXbar_in_1_d_bits_opcode = tlMasterXbar_portsDIO_filtered_1_bits_opcode ; 
  assign  tlMasterXbar_in_1_d_bits_param = tlMasterXbar_portsDIO_filtered_1_bits_param ; 
  assign  tlMasterXbar_in_1_d_bits_size = tlMasterXbar_portsDIO_filtered_1_bits_size ; 
  assign  tlMasterXbar_in_1_d_bits_source = tlMasterXbar_portsDIO_filtered_1_bits_source ; 
  assign  tlMasterXbar_in_1_d_bits_sink = tlMasterXbar_portsDIO_filtered_1_bits_sink ; 
  assign  tlMasterXbar_in_1_d_bits_denied = tlMasterXbar_portsDIO_filtered_1_bits_denied ; 
  assign  tlMasterXbar_in_1_d_bits_data = tlMasterXbar_portsDIO_filtered_1_bits_data ; 
  assign  tlMasterXbar_in_1_d_bits_corrupt = tlMasterXbar_portsDIO_filtered_1_bits_corrupt ; 
  assign  tlMasterXbar_portsDIO_filtered_0_valid = tlMasterXbar_out_0_d_valid & tlMasterXbar_requestDOI_0_0 ; 
  assign  tlMasterXbar_portsDIO_filtered_1_valid = tlMasterXbar_out_0_d_valid & tlMasterXbar_requestDOI_0_1 ; 
  assign  tlMasterXbar__portsDIO_out_0_d_ready_WIRE =( tlMasterXbar_requestDOI_0_0  ?  tlMasterXbar_portsDIO_filtered_0_ready :1'h0)|( tlMasterXbar_requestDOI_0_1  ?  tlMasterXbar_portsDIO_filtered_1_ready :1'h0); 
  assign  tlMasterXbar_out_0_d_ready = tlMasterXbar__portsDIO_out_0_d_ready_WIRE ; 
  assign  tlMasterXbar_in_0_e_ready = tlMasterXbar_portsEOI_filtered_0_ready ; 
  assign  tlMasterXbar_out_0_e_valid = tlMasterXbar_portsEOI_filtered_0_valid ; 
  assign  tlMasterXbar_out_0_e_bits_sink = tlMasterXbar_portsEOI_filtered_0_bits_sink ; 
    wire tlMasterXbar_in_1_e_ready = tlMasterXbar_portsEOI_filtered_1_0_ready ; reg[8:0] tlMasterXbar_beatsLeft ; 
    wire tlMasterXbar_idle = tlMasterXbar_beatsLeft ==9'h0; 
    wire tlMasterXbar_latch = tlMasterXbar_idle & tlMasterXbar_out_0_a_ready ; 
    wire[1:0] tlMasterXbar_readys_valid ={ tlMasterXbar_portsAOI_filtered_1_0_valid , tlMasterXbar_portsAOI_filtered_0_valid }; 
    wire tlMasterXbar__GEN_127 = tlMasterXbar_readys_valid == tlMasterXbar_readys_valid ==1'h0; reg[1:0] tlMasterXbar_readys_mask ; 
    wire[3:0] tlMasterXbar_readys_filter ={ tlMasterXbar_readys_valid &~ tlMasterXbar_readys_mask , tlMasterXbar_readys_valid }; 
    wire[3:0] tlMasterXbar__GEN_128 = tlMasterXbar_readys_filter |{1'h0, tlMasterXbar_readys_filter [3:1]}; 
    wire[3:0] tlMasterXbar_readys_unready ={1'h0, tlMasterXbar__GEN_128 [3:1]}|{ tlMasterXbar_readys_mask ,2'h0}; 
    wire[1:0] tlMasterXbar_readys_readys =~( tlMasterXbar_readys_unready [3:2]& tlMasterXbar_readys_unready [1:0]); 
    wire tlMasterXbar__GEN_129 = tlMasterXbar_latch &(| tlMasterXbar_readys_valid ); 
    wire[1:0] tlMasterXbar__GEN_130 = tlMasterXbar_readys_readys & tlMasterXbar_readys_valid ; 
    wire[2:0] tlMasterXbar__GEN_131 ={ tlMasterXbar__GEN_130 ,1'h0}; 
    wire[1:0] tlMasterXbar__GEN_132 = tlMasterXbar__GEN_130 | tlMasterXbar__GEN_131 [1:0]; 
    wire tlMasterXbar_readys_0 = tlMasterXbar_readys_readys [0]; 
    wire tlMasterXbar_readys_1 = tlMasterXbar_readys_readys [1]; 
    wire tlMasterXbar_winner_0 = tlMasterXbar_readys_0 & tlMasterXbar_portsAOI_filtered_0_valid ; 
    wire tlMasterXbar_winner_1 = tlMasterXbar_readys_1 & tlMasterXbar_portsAOI_filtered_1_0_valid ; 
    wire tlMasterXbar_prefixOR_1 = tlMasterXbar_winner_0 |1'h0; 
    wire tlMasterXbar__GEN_133 =(( tlMasterXbar_prefixOR_1 ==1'h0| tlMasterXbar_winner_1 ==1'h0)&1'h1)==1'h0; 
    wire tlMasterXbar__GEN_134 =(( tlMasterXbar_portsAOI_filtered_0_valid | tlMasterXbar_portsAOI_filtered_1_0_valid )==1'h0| tlMasterXbar_winner_0 | tlMasterXbar_winner_1 )==1'h0; 
  always @( posedge  tlMasterXbar_clock )
         begin 
             if ( tlMasterXbar_reset ==1'h0& tlMasterXbar__GEN_127 )
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:22 assert (valid === valids)\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_reset ==1'h0& tlMasterXbar__GEN_133 )
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:77 assert((prefixOR zip winner) map { case (p,w) => !p || !w } reduce {_ && _})\n");
                     if (1)$fatal;
                 end 
             if ( tlMasterXbar_reset ==1'h0& tlMasterXbar__GEN_134 )
                 begin 
                     if (1)$error("Assertion failed\n    at Arbiter.scala:79 assert (!valids.reduce(_||_) || winner.reduce(_||_))\n");
                     if (1)$fatal;
                 end 
         end
    wire[8:0] tlMasterXbar_maskedBeats_0 = tlMasterXbar_winner_0  ?  tlMasterXbar_beatsAI_0 :9'h0; 
    wire[8:0] tlMasterXbar_maskedBeats_1 = tlMasterXbar_winner_1  ?  tlMasterXbar_beatsAI_1 :9'h0; 
    wire[8:0] tlMasterXbar_initBeats = tlMasterXbar_maskedBeats_0 | tlMasterXbar_maskedBeats_1 ; 
    wire[9:0] tlMasterXbar__GEN_135 ={1'h0, tlMasterXbar_beatsLeft }-{9'h0, tlMasterXbar_out_0_a_ready & tlMasterXbar_out_0_a_valid }; 
    reg tlMasterXbar_state_0 ; 
    reg tlMasterXbar_state_1 ; 
    wire tlMasterXbar_muxState_0 = tlMasterXbar_idle  ?  tlMasterXbar_winner_0 : tlMasterXbar_state_0 ; 
    wire tlMasterXbar_muxState_1 = tlMasterXbar_idle  ?  tlMasterXbar_winner_1 : tlMasterXbar_state_1 ; 
    wire tlMasterXbar_allowed_0 = tlMasterXbar_idle  ?  tlMasterXbar_readys_0 : tlMasterXbar_state_0 ; 
    wire tlMasterXbar_allowed_1 = tlMasterXbar_idle  ?  tlMasterXbar_readys_1 : tlMasterXbar_state_1 ; 
  assign  tlMasterXbar_portsAOI_filtered_0_ready = tlMasterXbar_out_0_a_ready & tlMasterXbar_allowed_0 ; 
  assign  tlMasterXbar_portsAOI_filtered_1_0_ready = tlMasterXbar_out_0_a_ready & tlMasterXbar_allowed_1 ; 
    wire tlMasterXbar__out_0_a_valid_WIRE =( tlMasterXbar_state_0  ?  tlMasterXbar_portsAOI_filtered_0_valid :1'h0)|( tlMasterXbar_state_1  ?  tlMasterXbar_portsAOI_filtered_1_0_valid :1'h0); 
  assign  tlMasterXbar_out_0_a_valid = tlMasterXbar_idle  ?  tlMasterXbar_portsAOI_filtered_0_valid | tlMasterXbar_portsAOI_filtered_1_0_valid : tlMasterXbar__out_0_a_valid_WIRE ; 
    wire[2:0] tlMasterXbar__out_0_a_bits_WIRE_18 ; 
  assign  tlMasterXbar_out_0_a_bits_opcode = tlMasterXbar__out_0_a_bits_WIRE_opcode ; 
    wire[2:0] tlMasterXbar__out_0_a_bits_WIRE_17 ; 
  assign  tlMasterXbar_out_0_a_bits_param = tlMasterXbar__out_0_a_bits_WIRE_param ; 
    wire[3:0] tlMasterXbar__out_0_a_bits_WIRE_16 ; 
  assign  tlMasterXbar_out_0_a_bits_size = tlMasterXbar__out_0_a_bits_WIRE_size ; 
    wire[1:0] tlMasterXbar__out_0_a_bits_WIRE_15 ; 
  assign  tlMasterXbar_out_0_a_bits_source = tlMasterXbar__out_0_a_bits_WIRE_source ; 
    wire[31:0] tlMasterXbar__out_0_a_bits_WIRE_14 ; 
  assign  tlMasterXbar_out_0_a_bits_address = tlMasterXbar__out_0_a_bits_WIRE_address ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_bufferable ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_bufferable = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_bufferable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_modifiable ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_modifiable = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_modifiable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_readalloc ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_readalloc = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_readalloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_writealloc ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_writealloc = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_writealloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_privileged ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_privileged = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_privileged ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_secure ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_secure = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_secure ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_fetch ; 
  assign  tlMasterXbar_out_0_a_bits_user_amba_prot_fetch = tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_fetch ; 
    wire[7:0] tlMasterXbar__out_0_a_bits_WIRE_3 ; 
  assign  tlMasterXbar_out_0_a_bits_mask = tlMasterXbar__out_0_a_bits_WIRE_mask ; 
    wire[63:0] tlMasterXbar__out_0_a_bits_WIRE_2 ; 
  assign  tlMasterXbar_out_0_a_bits_data = tlMasterXbar__out_0_a_bits_WIRE_data ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_1 ; 
  assign  tlMasterXbar_out_0_a_bits_corrupt = tlMasterXbar__out_0_a_bits_WIRE_corrupt ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_1 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_corrupt :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_corrupt :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_corrupt = tlMasterXbar__out_0_a_bits_WIRE_1 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_2 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_data :64'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_data :64'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_data = tlMasterXbar__out_0_a_bits_WIRE_2 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_3 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_mask :8'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_mask :8'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_mask = tlMasterXbar__out_0_a_bits_WIRE_3 ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_bufferable ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_bufferable = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_bufferable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_modifiable ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_modifiable = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_modifiable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_readalloc ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_readalloc = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_readalloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_writealloc ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_writealloc = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_writealloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_privileged ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_privileged = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_privileged ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_secure ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_secure = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_secure ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_6_fetch ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_user_amba_prot_fetch = tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_fetch ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_13 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_bufferable = tlMasterXbar__out_0_a_bits_WIRE_6_bufferable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_12 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_modifiable = tlMasterXbar__out_0_a_bits_WIRE_6_modifiable ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_11 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_readalloc = tlMasterXbar__out_0_a_bits_WIRE_6_readalloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_10 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_writealloc = tlMasterXbar__out_0_a_bits_WIRE_6_writealloc ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_9 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_privileged = tlMasterXbar__out_0_a_bits_WIRE_6_privileged ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_8 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_secure = tlMasterXbar__out_0_a_bits_WIRE_6_secure ; 
    wire tlMasterXbar__out_0_a_bits_WIRE_7 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_5_amba_prot_fetch = tlMasterXbar__out_0_a_bits_WIRE_6_fetch ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_7 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_fetch :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_fetch :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_fetch = tlMasterXbar__out_0_a_bits_WIRE_7 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_8 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_secure :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_secure :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_secure = tlMasterXbar__out_0_a_bits_WIRE_8 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_9 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_privileged :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_privileged :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_privileged = tlMasterXbar__out_0_a_bits_WIRE_9 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_10 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_writealloc :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_writealloc :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_writealloc = tlMasterXbar__out_0_a_bits_WIRE_10 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_11 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_readalloc :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_readalloc :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_readalloc = tlMasterXbar__out_0_a_bits_WIRE_11 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_12 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_modifiable :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_modifiable :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_modifiable = tlMasterXbar__out_0_a_bits_WIRE_12 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_13 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_user_amba_prot_bufferable :1'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_user_amba_prot_bufferable :1'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_6_bufferable = tlMasterXbar__out_0_a_bits_WIRE_13 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_14 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_address :32'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_address :32'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_address = tlMasterXbar__out_0_a_bits_WIRE_14 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_15 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_source :2'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_source :2'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_source = tlMasterXbar__out_0_a_bits_WIRE_15 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_16 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_size :4'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_size :4'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_size = tlMasterXbar__out_0_a_bits_WIRE_16 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_17 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_param :3'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_param :3'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_param = tlMasterXbar__out_0_a_bits_WIRE_17 ; 
  assign  tlMasterXbar__out_0_a_bits_WIRE_18 =( tlMasterXbar_muxState_0  ?  tlMasterXbar_portsAOI_filtered_0_bits_opcode :3'h0)|( tlMasterXbar_muxState_1  ?  tlMasterXbar_portsAOI_filtered_1_0_bits_opcode :3'h0); 
  assign  tlMasterXbar__out_0_a_bits_WIRE_opcode = tlMasterXbar__out_0_a_bits_WIRE_18 ; 
  always @( posedge  tlMasterXbar_clock )
         begin 
             if ( tlMasterXbar_reset )
                 begin  
                     tlMasterXbar_beatsLeft  <=9'h0; 
                     tlMasterXbar_readys_mask  <=2'h3; 
                     tlMasterXbar_state_0  <= tlMasterXbar__state_WIRE_0 ; 
                     tlMasterXbar_state_1  <= tlMasterXbar__state_WIRE_1 ;
                 end 
              else 
                 begin 
                     if ( tlMasterXbar_latch ) 
                         tlMasterXbar_beatsLeft  <= tlMasterXbar_initBeats ;
                      else  
                         tlMasterXbar_beatsLeft  <= tlMasterXbar__GEN_135 [8:0];
                     if ( tlMasterXbar__GEN_129 ) 
                         tlMasterXbar_readys_mask  <= tlMasterXbar__GEN_132 ;
                      else 
                         begin 
                         end  
                     tlMasterXbar_state_0  <= tlMasterXbar_muxState_0 ; 
                     tlMasterXbar_state_1  <= tlMasterXbar_muxState_1 ;
                 end 
         end
  assign  tlMasterXbar_auto_in_1_a_ready = tlMasterXbar_nodeIn_1_a_ready ; 
  assign  tlMasterXbar_auto_in_1_d_valid = tlMasterXbar_nodeIn_1_d_valid ; 
  assign  tlMasterXbar_auto_in_1_d_bits_opcode = tlMasterXbar_nodeIn_1_d_bits_opcode ; 
  assign  tlMasterXbar_auto_in_1_d_bits_param = tlMasterXbar_nodeIn_1_d_bits_param ; 
  assign  tlMasterXbar_auto_in_1_d_bits_size = tlMasterXbar_nodeIn_1_d_bits_size ; 
  assign  tlMasterXbar_auto_in_1_d_bits_source = tlMasterXbar_nodeIn_1_d_bits_source ; 
  assign  tlMasterXbar_auto_in_1_d_bits_sink = tlMasterXbar_nodeIn_1_d_bits_sink ; 
  assign  tlMasterXbar_auto_in_1_d_bits_denied = tlMasterXbar_nodeIn_1_d_bits_denied ; 
  assign  tlMasterXbar_auto_in_1_d_bits_data = tlMasterXbar_nodeIn_1_d_bits_data ; 
  assign  tlMasterXbar_auto_in_1_d_bits_corrupt = tlMasterXbar_nodeIn_1_d_bits_corrupt ; 
  assign  tlMasterXbar_auto_in_0_a_ready = tlMasterXbar_nodeIn_a_ready ; 
  assign  tlMasterXbar_auto_in_0_b_valid = tlMasterXbar_nodeIn_b_valid ; 
  assign  tlMasterXbar_auto_in_0_b_bits_opcode = tlMasterXbar_nodeIn_b_bits_opcode ; 
  assign  tlMasterXbar_auto_in_0_b_bits_param = tlMasterXbar_nodeIn_b_bits_param ; 
  assign  tlMasterXbar_auto_in_0_b_bits_size = tlMasterXbar_nodeIn_b_bits_size ; 
  assign  tlMasterXbar_auto_in_0_b_bits_source = tlMasterXbar_nodeIn_b_bits_source ; 
  assign  tlMasterXbar_auto_in_0_b_bits_address = tlMasterXbar_nodeIn_b_bits_address ; 
  assign  tlMasterXbar_auto_in_0_b_bits_mask = tlMasterXbar_nodeIn_b_bits_mask ; 
  assign  tlMasterXbar_auto_in_0_b_bits_data = tlMasterXbar_nodeIn_b_bits_data ; 
  assign  tlMasterXbar_auto_in_0_b_bits_corrupt = tlMasterXbar_nodeIn_b_bits_corrupt ; 
  assign  tlMasterXbar_auto_in_0_c_ready = tlMasterXbar_nodeIn_c_ready ; 
  assign  tlMasterXbar_auto_in_0_d_valid = tlMasterXbar_nodeIn_d_valid ; 
  assign  tlMasterXbar_auto_in_0_d_bits_opcode = tlMasterXbar_nodeIn_d_bits_opcode ; 
  assign  tlMasterXbar_auto_in_0_d_bits_param = tlMasterXbar_nodeIn_d_bits_param ; 
  assign  tlMasterXbar_auto_in_0_d_bits_size = tlMasterXbar_nodeIn_d_bits_size ; 
  assign  tlMasterXbar_auto_in_0_d_bits_source = tlMasterXbar_nodeIn_d_bits_source ; 
  assign  tlMasterXbar_auto_in_0_d_bits_sink = tlMasterXbar_nodeIn_d_bits_sink ; 
  assign  tlMasterXbar_auto_in_0_d_bits_denied = tlMasterXbar_nodeIn_d_bits_denied ; 
  assign  tlMasterXbar_auto_in_0_d_bits_data = tlMasterXbar_nodeIn_d_bits_data ; 
  assign  tlMasterXbar_auto_in_0_d_bits_corrupt = tlMasterXbar_nodeIn_d_bits_corrupt ; 
  assign  tlMasterXbar_auto_in_0_e_ready = tlMasterXbar_nodeIn_e_ready ; 
  assign  tlMasterXbar_auto_out_a_valid = tlMasterXbar_nodeOut_a_valid ; 
  assign  tlMasterXbar_auto_out_a_bits_opcode = tlMasterXbar_nodeOut_a_bits_opcode ; 
  assign  tlMasterXbar_auto_out_a_bits_param = tlMasterXbar_nodeOut_a_bits_param ; 
  assign  tlMasterXbar_auto_out_a_bits_size = tlMasterXbar_nodeOut_a_bits_size ; 
  assign  tlMasterXbar_auto_out_a_bits_source = tlMasterXbar_nodeOut_a_bits_source ; 
  assign  tlMasterXbar_auto_out_a_bits_address = tlMasterXbar_nodeOut_a_bits_address ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable = tlMasterXbar_nodeOut_a_bits_user_amba_prot_bufferable ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable = tlMasterXbar_nodeOut_a_bits_user_amba_prot_modifiable ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc = tlMasterXbar_nodeOut_a_bits_user_amba_prot_readalloc ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc = tlMasterXbar_nodeOut_a_bits_user_amba_prot_writealloc ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged = tlMasterXbar_nodeOut_a_bits_user_amba_prot_privileged ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_secure = tlMasterXbar_nodeOut_a_bits_user_amba_prot_secure ; 
  assign  tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch = tlMasterXbar_nodeOut_a_bits_user_amba_prot_fetch ; 
  assign  tlMasterXbar_auto_out_a_bits_mask = tlMasterXbar_nodeOut_a_bits_mask ; 
  assign  tlMasterXbar_auto_out_a_bits_data = tlMasterXbar_nodeOut_a_bits_data ; 
  assign  tlMasterXbar_auto_out_a_bits_corrupt = tlMasterXbar_nodeOut_a_bits_corrupt ; 
  assign  tlMasterXbar_auto_out_b_ready = tlMasterXbar_nodeOut_b_ready ; 
  assign  tlMasterXbar_auto_out_c_valid = tlMasterXbar_nodeOut_c_valid ; 
  assign  tlMasterXbar_auto_out_c_bits_opcode = tlMasterXbar_nodeOut_c_bits_opcode ; 
  assign  tlMasterXbar_auto_out_c_bits_param = tlMasterXbar_nodeOut_c_bits_param ; 
  assign  tlMasterXbar_auto_out_c_bits_size = tlMasterXbar_nodeOut_c_bits_size ; 
  assign  tlMasterXbar_auto_out_c_bits_source = tlMasterXbar_nodeOut_c_bits_source ; 
  assign  tlMasterXbar_auto_out_c_bits_address = tlMasterXbar_nodeOut_c_bits_address ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_bufferable = tlMasterXbar_nodeOut_c_bits_user_amba_prot_bufferable ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_modifiable = tlMasterXbar_nodeOut_c_bits_user_amba_prot_modifiable ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_readalloc = tlMasterXbar_nodeOut_c_bits_user_amba_prot_readalloc ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_writealloc = tlMasterXbar_nodeOut_c_bits_user_amba_prot_writealloc ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_privileged = tlMasterXbar_nodeOut_c_bits_user_amba_prot_privileged ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_secure = tlMasterXbar_nodeOut_c_bits_user_amba_prot_secure ; 
  assign  tlMasterXbar_auto_out_c_bits_user_amba_prot_fetch = tlMasterXbar_nodeOut_c_bits_user_amba_prot_fetch ; 
  assign  tlMasterXbar_auto_out_c_bits_data = tlMasterXbar_nodeOut_c_bits_data ; 
  assign  tlMasterXbar_auto_out_c_bits_corrupt = tlMasterXbar_nodeOut_c_bits_corrupt ; 
  assign  tlMasterXbar_auto_out_d_ready = tlMasterXbar_nodeOut_d_ready ; 
  assign  tlMasterXbar_auto_out_e_valid = tlMasterXbar_nodeOut_e_valid ; 
  assign  tlMasterXbar_auto_out_e_bits_sink = tlMasterXbar_nodeOut_e_bits_sink ;
    assign tlMasterXbar_clock = clock;
    assign tlMasterXbar_reset = reset;
    assign widget_1_auto_out_a_ready = tlMasterXbar_auto_in_1_a_ready;
    assign tlMasterXbar_auto_in_1_a_valid = widget_1_auto_out_a_valid;
    assign tlMasterXbar_auto_in_1_a_bits_opcode = widget_1_auto_out_a_bits_opcode;
    assign tlMasterXbar_auto_in_1_a_bits_param = widget_1_auto_out_a_bits_param;
    assign tlMasterXbar_auto_in_1_a_bits_size = widget_1_auto_out_a_bits_size;
    assign tlMasterXbar_auto_in_1_a_bits_source = widget_1_auto_out_a_bits_source;
    assign tlMasterXbar_auto_in_1_a_bits_address = widget_1_auto_out_a_bits_address;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_bufferable = widget_1_auto_out_a_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_modifiable = widget_1_auto_out_a_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_readalloc = widget_1_auto_out_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_writealloc = widget_1_auto_out_a_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_privileged = widget_1_auto_out_a_bits_user_amba_prot_privileged;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_secure = widget_1_auto_out_a_bits_user_amba_prot_secure;
    assign tlMasterXbar_auto_in_1_a_bits_user_amba_prot_fetch = widget_1_auto_out_a_bits_user_amba_prot_fetch;
    assign tlMasterXbar_auto_in_1_a_bits_mask = widget_1_auto_out_a_bits_mask;
    assign tlMasterXbar_auto_in_1_a_bits_data = widget_1_auto_out_a_bits_data;
    assign tlMasterXbar_auto_in_1_a_bits_corrupt = widget_1_auto_out_a_bits_corrupt;
    assign tlMasterXbar_auto_in_1_d_ready = widget_1_auto_out_d_ready;
    assign widget_1_auto_out_d_valid = tlMasterXbar_auto_in_1_d_valid;
    assign widget_1_auto_out_d_bits_opcode = tlMasterXbar_auto_in_1_d_bits_opcode;
    assign widget_1_auto_out_d_bits_param = tlMasterXbar_auto_in_1_d_bits_param;
    assign widget_1_auto_out_d_bits_size = tlMasterXbar_auto_in_1_d_bits_size;
    assign widget_1_auto_out_d_bits_source = tlMasterXbar_auto_in_1_d_bits_source;
    assign widget_1_auto_out_d_bits_sink = tlMasterXbar_auto_in_1_d_bits_sink;
    assign widget_1_auto_out_d_bits_denied = tlMasterXbar_auto_in_1_d_bits_denied;
    assign widget_1_auto_out_d_bits_data = tlMasterXbar_auto_in_1_d_bits_data;
    assign widget_1_auto_out_d_bits_corrupt = tlMasterXbar_auto_in_1_d_bits_corrupt;
    assign widget_auto_out_a_ready = tlMasterXbar_auto_in_0_a_ready;
    assign tlMasterXbar_auto_in_0_a_valid = widget_auto_out_a_valid;
    assign tlMasterXbar_auto_in_0_a_bits_opcode = widget_auto_out_a_bits_opcode;
    assign tlMasterXbar_auto_in_0_a_bits_param = widget_auto_out_a_bits_param;
    assign tlMasterXbar_auto_in_0_a_bits_size = widget_auto_out_a_bits_size;
    assign tlMasterXbar_auto_in_0_a_bits_source = widget_auto_out_a_bits_source;
    assign tlMasterXbar_auto_in_0_a_bits_address = widget_auto_out_a_bits_address;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_bufferable = widget_auto_out_a_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_modifiable = widget_auto_out_a_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_readalloc = widget_auto_out_a_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_writealloc = widget_auto_out_a_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_privileged = widget_auto_out_a_bits_user_amba_prot_privileged;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_secure = widget_auto_out_a_bits_user_amba_prot_secure;
    assign tlMasterXbar_auto_in_0_a_bits_user_amba_prot_fetch = widget_auto_out_a_bits_user_amba_prot_fetch;
    assign tlMasterXbar_auto_in_0_a_bits_mask = widget_auto_out_a_bits_mask;
    assign tlMasterXbar_auto_in_0_a_bits_data = widget_auto_out_a_bits_data;
    assign tlMasterXbar_auto_in_0_a_bits_corrupt = widget_auto_out_a_bits_corrupt;
    assign tlMasterXbar_auto_in_0_b_ready = widget_auto_out_b_ready;
    assign widget_auto_out_b_valid = tlMasterXbar_auto_in_0_b_valid;
    assign widget_auto_out_b_bits_opcode = tlMasterXbar_auto_in_0_b_bits_opcode;
    assign widget_auto_out_b_bits_param = tlMasterXbar_auto_in_0_b_bits_param;
    assign widget_auto_out_b_bits_size = tlMasterXbar_auto_in_0_b_bits_size;
    assign widget_auto_out_b_bits_source = tlMasterXbar_auto_in_0_b_bits_source;
    assign widget_auto_out_b_bits_address = tlMasterXbar_auto_in_0_b_bits_address;
    assign widget_auto_out_b_bits_mask = tlMasterXbar_auto_in_0_b_bits_mask;
    assign widget_auto_out_b_bits_data = tlMasterXbar_auto_in_0_b_bits_data;
    assign widget_auto_out_b_bits_corrupt = tlMasterXbar_auto_in_0_b_bits_corrupt;
    assign widget_auto_out_c_ready = tlMasterXbar_auto_in_0_c_ready;
    assign tlMasterXbar_auto_in_0_c_valid = widget_auto_out_c_valid;
    assign tlMasterXbar_auto_in_0_c_bits_opcode = widget_auto_out_c_bits_opcode;
    assign tlMasterXbar_auto_in_0_c_bits_param = widget_auto_out_c_bits_param;
    assign tlMasterXbar_auto_in_0_c_bits_size = widget_auto_out_c_bits_size;
    assign tlMasterXbar_auto_in_0_c_bits_source = widget_auto_out_c_bits_source;
    assign tlMasterXbar_auto_in_0_c_bits_address = widget_auto_out_c_bits_address;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_bufferable = widget_auto_out_c_bits_user_amba_prot_bufferable;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_modifiable = widget_auto_out_c_bits_user_amba_prot_modifiable;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_readalloc = widget_auto_out_c_bits_user_amba_prot_readalloc;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_writealloc = widget_auto_out_c_bits_user_amba_prot_writealloc;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_privileged = widget_auto_out_c_bits_user_amba_prot_privileged;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_secure = widget_auto_out_c_bits_user_amba_prot_secure;
    assign tlMasterXbar_auto_in_0_c_bits_user_amba_prot_fetch = widget_auto_out_c_bits_user_amba_prot_fetch;
    assign tlMasterXbar_auto_in_0_c_bits_data = widget_auto_out_c_bits_data;
    assign tlMasterXbar_auto_in_0_c_bits_corrupt = widget_auto_out_c_bits_corrupt;
    assign tlMasterXbar_auto_in_0_d_ready = widget_auto_out_d_ready;
    assign widget_auto_out_d_valid = tlMasterXbar_auto_in_0_d_valid;
    assign widget_auto_out_d_bits_opcode = tlMasterXbar_auto_in_0_d_bits_opcode;
    assign widget_auto_out_d_bits_param = tlMasterXbar_auto_in_0_d_bits_param;
    assign widget_auto_out_d_bits_size = tlMasterXbar_auto_in_0_d_bits_size;
    assign widget_auto_out_d_bits_source = tlMasterXbar_auto_in_0_d_bits_source;
    assign widget_auto_out_d_bits_sink = tlMasterXbar_auto_in_0_d_bits_sink;
    assign widget_auto_out_d_bits_denied = tlMasterXbar_auto_in_0_d_bits_denied;
    assign widget_auto_out_d_bits_data = tlMasterXbar_auto_in_0_d_bits_data;
    assign widget_auto_out_d_bits_corrupt = tlMasterXbar_auto_in_0_d_bits_corrupt;
    assign widget_auto_out_e_ready = tlMasterXbar_auto_in_0_e_ready;
    assign tlMasterXbar_auto_in_0_e_valid = widget_auto_out_e_valid;
    assign tlMasterXbar_auto_in_0_e_bits_sink = widget_auto_out_e_bits_sink;
    assign tlMasterXbar_auto_out_a_ready = tlOtherMastersNodeIn_a_ready;
    assign tlOtherMastersNodeIn_a_valid = tlMasterXbar_auto_out_a_valid;
    assign tlOtherMastersNodeIn_a_bits_opcode = tlMasterXbar_auto_out_a_bits_opcode;
    assign tlOtherMastersNodeIn_a_bits_param = tlMasterXbar_auto_out_a_bits_param;
    assign tlOtherMastersNodeIn_a_bits_size = tlMasterXbar_auto_out_a_bits_size;
    assign tlOtherMastersNodeIn_a_bits_source = tlMasterXbar_auto_out_a_bits_source;
    assign tlOtherMastersNodeIn_a_bits_address = tlMasterXbar_auto_out_a_bits_address;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_bufferable = tlMasterXbar_auto_out_a_bits_user_amba_prot_bufferable;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_modifiable = tlMasterXbar_auto_out_a_bits_user_amba_prot_modifiable;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_readalloc = tlMasterXbar_auto_out_a_bits_user_amba_prot_readalloc;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_writealloc = tlMasterXbar_auto_out_a_bits_user_amba_prot_writealloc;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_privileged = tlMasterXbar_auto_out_a_bits_user_amba_prot_privileged;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_secure = tlMasterXbar_auto_out_a_bits_user_amba_prot_secure;
    assign tlOtherMastersNodeIn_a_bits_user_amba_prot_fetch = tlMasterXbar_auto_out_a_bits_user_amba_prot_fetch;
    assign tlOtherMastersNodeIn_a_bits_mask = tlMasterXbar_auto_out_a_bits_mask;
    assign tlOtherMastersNodeIn_a_bits_data = tlMasterXbar_auto_out_a_bits_data;
    assign tlOtherMastersNodeIn_a_bits_corrupt = tlMasterXbar_auto_out_a_bits_corrupt;
    assign tlOtherMastersNodeIn_b_ready = tlMasterXbar_auto_out_b_ready;
    assign tlMasterXbar_auto_out_b_valid = tlOtherMastersNodeIn_b_valid;
    assign tlMasterXbar_auto_out_b_bits_opcode = tlOtherMastersNodeIn_b_bits_opcode;
    assign tlMasterXbar_auto_out_b_bits_param = tlOtherMastersNodeIn_b_bits_param;
    assign tlMasterXbar_auto_out_b_bits_size = tlOtherMastersNodeIn_b_bits_size;
    assign tlMasterXbar_auto_out_b_bits_source = tlOtherMastersNodeIn_b_bits_source;
    assign tlMasterXbar_auto_out_b_bits_address = tlOtherMastersNodeIn_b_bits_address;
    assign tlMasterXbar_auto_out_b_bits_mask = tlOtherMastersNodeIn_b_bits_mask;
    assign tlMasterXbar_auto_out_b_bits_data = tlOtherMastersNodeIn_b_bits_data;
    assign tlMasterXbar_auto_out_b_bits_corrupt = tlOtherMastersNodeIn_b_bits_corrupt;
    assign tlMasterXbar_auto_out_c_ready = tlOtherMastersNodeIn_c_ready;
    assign tlOtherMastersNodeIn_c_valid = tlMasterXbar_auto_out_c_valid;
    assign tlOtherMastersNodeIn_c_bits_opcode = tlMasterXbar_auto_out_c_bits_opcode;
    assign tlOtherMastersNodeIn_c_bits_param = tlMasterXbar_auto_out_c_bits_param;
    assign tlOtherMastersNodeIn_c_bits_size = tlMasterXbar_auto_out_c_bits_size;
    assign tlOtherMastersNodeIn_c_bits_source = tlMasterXbar_auto_out_c_bits_source;
    assign tlOtherMastersNodeIn_c_bits_address = tlMasterXbar_auto_out_c_bits_address;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_bufferable = tlMasterXbar_auto_out_c_bits_user_amba_prot_bufferable;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_modifiable = tlMasterXbar_auto_out_c_bits_user_amba_prot_modifiable;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_readalloc = tlMasterXbar_auto_out_c_bits_user_amba_prot_readalloc;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_writealloc = tlMasterXbar_auto_out_c_bits_user_amba_prot_writealloc;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_privileged = tlMasterXbar_auto_out_c_bits_user_amba_prot_privileged;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_secure = tlMasterXbar_auto_out_c_bits_user_amba_prot_secure;
    assign tlOtherMastersNodeIn_c_bits_user_amba_prot_fetch = tlMasterXbar_auto_out_c_bits_user_amba_prot_fetch;
    assign tlOtherMastersNodeIn_c_bits_data = tlMasterXbar_auto_out_c_bits_data;
    assign tlOtherMastersNodeIn_c_bits_corrupt = tlMasterXbar_auto_out_c_bits_corrupt;
    assign tlOtherMastersNodeIn_d_ready = tlMasterXbar_auto_out_d_ready;
    assign tlMasterXbar_auto_out_d_valid = tlOtherMastersNodeIn_d_valid;
    assign tlMasterXbar_auto_out_d_bits_opcode = tlOtherMastersNodeIn_d_bits_opcode;
    assign tlMasterXbar_auto_out_d_bits_param = tlOtherMastersNodeIn_d_bits_param;
    assign tlMasterXbar_auto_out_d_bits_size = tlOtherMastersNodeIn_d_bits_size;
    assign tlMasterXbar_auto_out_d_bits_source = tlOtherMastersNodeIn_d_bits_source;
    assign tlMasterXbar_auto_out_d_bits_sink = tlOtherMastersNodeIn_d_bits_sink;
    assign tlMasterXbar_auto_out_d_bits_denied = tlOtherMastersNodeIn_d_bits_denied;
    assign tlMasterXbar_auto_out_d_bits_data = tlOtherMastersNodeIn_d_bits_data;
    assign tlMasterXbar_auto_out_d_bits_corrupt = tlOtherMastersNodeIn_d_bits_corrupt;
    assign tlMasterXbar_auto_out_e_ready = tlOtherMastersNodeIn_e_ready;
    assign tlOtherMastersNodeIn_e_valid = tlMasterXbar_auto_out_e_valid;
    assign tlOtherMastersNodeIn_e_bits_sink = tlMasterXbar_auto_out_e_bits_sink;
    
  wire tlSlaveXbar_clock;
    wire tlSlaveXbar_reset;

    
    assign tlSlaveXbar_clock = clock;
    assign tlSlaveXbar_reset = reset;
    
  wire        int_localOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        x1_int_localOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        x1_int_localOut_1;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        x1_int_localOut_1_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire intXbar_clock;
    wire intXbar_reset;
    wire intXbar_auto_int_in_2_0;
    wire intXbar_auto_int_in_1_0;
    wire intXbar_auto_int_in_1_1;
    wire intXbar_auto_int_in_0_0;
    wire intXbar_auto_int_out_0;
    wire intXbar_auto_int_out_1;
    wire intXbar_auto_int_out_2;
    wire intXbar_auto_int_out_3;

    wire intXbar_intnodeIn_0 = intXbar_auto_int_in_0_0 ; 
    wire intXbar_intnodeIn_1_0 = intXbar_auto_int_in_1_0 ; 
    wire intXbar_intnodeIn_1_1 = intXbar_auto_int_in_1_1 ; 
    wire intXbar_intnodeIn_2_0 = intXbar_auto_int_in_2_0 ; 
    wire intXbar_intnodeOut_0 = intXbar_intnodeIn_0 ; 
    wire intXbar_intnodeOut_1 = intXbar_intnodeIn_1_0 ; 
    wire intXbar_intnodeOut_2 = intXbar_intnodeIn_1_1 ; 
    wire intXbar_intnodeOut_3 = intXbar_intnodeIn_2_0 ; 
  assign  intXbar_auto_int_out_0 = intXbar_intnodeOut_0 ; 
  assign  intXbar_auto_int_out_1 = intXbar_intnodeOut_1 ; 
  assign  intXbar_auto_int_out_2 = intXbar_intnodeOut_2 ; 
  assign  intXbar_auto_int_out_3 = intXbar_intnodeOut_3 ;
    assign intXbar_clock = clock;
    assign intXbar_reset = reset;
    assign intXbar_auto_int_in_2_0 = x1_int_localOut_1_0;
    assign intXbar_auto_int_in_1_0 = x1_int_localOut_0;
    assign intXbar_auto_int_in_1_1 = x1_int_localOut_1;
    assign intXbar_auto_int_in_0_0 = int_localOut_0;
    assign intSinkNodeIn_0 = intXbar_auto_int_out_0;
    assign intSinkNodeIn_1 = intXbar_auto_int_out_1;
    assign intSinkNodeIn_2 = intXbar_auto_int_out_2;
    assign intSinkNodeIn_3 = intXbar_auto_int_out_3;
    
  wire        hartidOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_nodeIn = broadcast_auto_in;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        hartIdSinkNodeIn = broadcast_auto_out;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign broadcast_nodeOut = broadcast_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_auto_out = broadcast_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] reset_vectorOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_1_nodeIn = broadcast_1_auto_in;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_1_x1_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_1_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] resetVectorSinkNodeIn = broadcast_1_auto_out_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign broadcast_1_nodeOut = broadcast_1_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_1_x1_nodeOut = broadcast_1_nodeIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_1_auto_out_0 = broadcast_1_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_1_auto_out_1 = broadcast_1_x1_nodeOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        nmiOut_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_2_nodeIn_rnmi = broadcast_2_auto_in_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] nmiOut_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_2_nodeIn_rnmi_interrupt_vector =
    broadcast_2_auto_in_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] nmiOut_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_2_nodeIn_rnmi_exception_vector =
    broadcast_2_auto_in_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_2_nodeOut_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_2_nodeOut_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        nmiSinkNodeIn_rnmi = broadcast_2_auto_out_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] broadcast_2_nodeOut_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] nmiSinkNodeIn_rnmi_interrupt_vector =
    broadcast_2_auto_out_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] nmiSinkNodeIn_rnmi_exception_vector =
    broadcast_2_auto_out_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign broadcast_2_nodeOut_rnmi = broadcast_2_nodeIn_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_2_nodeOut_rnmi_interrupt_vector =
    broadcast_2_nodeIn_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_2_nodeOut_rnmi_exception_vector =
    broadcast_2_nodeIn_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_2_auto_out_rnmi = broadcast_2_nodeOut_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_2_auto_out_rnmi_interrupt_vector =
    broadcast_2_nodeOut_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_2_auto_out_rnmi_exception_vector =
    broadcast_2_nodeOut_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        traceSourceNodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeIn_insns_0_valid = broadcast_3_auto_in_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [33:0] traceSourceNodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_nodeIn_insns_0_iaddr = broadcast_3_auto_in_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] traceSourceNodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeIn_insns_0_insn = broadcast_3_auto_in_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  traceSourceNodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  broadcast_3_nodeIn_insns_0_priv = broadcast_3_auto_in_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        traceSourceNodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeIn_insns_0_exception =
    broadcast_3_auto_in_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        traceSourceNodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeIn_insns_0_interrupt =
    broadcast_3_auto_in_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] traceSourceNodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeIn_insns_0_cause = broadcast_3_auto_in_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [33:0] traceSourceNodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_nodeIn_insns_0_tval = broadcast_3_auto_in_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] traceSourceNodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeIn_time = broadcast_3_auto_in_time;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        broadcast_3_nodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_nodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_nodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  broadcast_3_nodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_nodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_nodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_nodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_nodeOut_insns_0_valid = broadcast_3_nodeIn_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_iaddr = broadcast_3_nodeIn_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_insn = broadcast_3_nodeIn_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_priv = broadcast_3_nodeIn_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_exception = broadcast_3_nodeIn_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_interrupt = broadcast_3_nodeIn_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_cause = broadcast_3_nodeIn_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_insns_0_tval = broadcast_3_nodeIn_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_nodeOut_time = broadcast_3_nodeIn_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        broadcast_3_auto_out_insns_0_valid = broadcast_3_nodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_auto_out_insns_0_iaddr = broadcast_3_nodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] broadcast_3_auto_out_insns_0_insn = broadcast_3_nodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  broadcast_3_auto_out_insns_0_priv = broadcast_3_nodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_auto_out_insns_0_exception =
    broadcast_3_nodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_3_auto_out_insns_0_interrupt =
    broadcast_3_nodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_auto_out_insns_0_cause = broadcast_3_nodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [33:0] broadcast_3_auto_out_insns_0_tval = broadcast_3_nodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] broadcast_3_auto_out_time = broadcast_3_nodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        nexus_1_nodeOut_enable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        nexus_1_nodeOut_stall;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        traceAuxSinkNodeIn_enable = nexus_1_auto_out_enable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        traceAuxSinkNodeIn_stall = nexus_1_auto_out_stall;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign nexus_1_auto_out_enable = nexus_1_nodeOut_enable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign nexus_1_auto_out_stall = nexus_1_nodeOut_stall;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign nexus_1_nodeOut_enable = nexus_1_defaultWireOpt_enable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:294:19
  assign nexus_1_nodeOut_stall = nexus_1_defaultWireOpt_stall;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/BaseTile.scala:294:19
  wire        bpwatchSourceNodeOut_0_valid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_4_nodeIn_0_valid_0 = broadcast_4_auto_in_0_valid_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        bpwatchSourceNodeOut_0_rvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_4_nodeIn_0_rvalid_0 = broadcast_4_auto_in_0_rvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        bpwatchSourceNodeOut_0_wvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_4_nodeIn_0_wvalid_0 = broadcast_4_auto_in_0_wvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        bpwatchSourceNodeOut_0_ivalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        broadcast_4_nodeIn_0_ivalid_0 = broadcast_4_auto_in_0_ivalid_0;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  bpwatchSourceNodeOut_0_action;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  broadcast_4_nodeIn_0_action = broadcast_4_auto_in_0_action;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_valid = widget_auto_in_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_a_bits_opcode = widget_auto_in_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_a_bits_param = widget_auto_in_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_a_bits_size = widget_auto_in_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_source = widget_auto_in_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_nodeIn_a_bits_address = widget_auto_in_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_bufferable =
    widget_auto_in_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_modifiable =
    widget_auto_in_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_readalloc =
    widget_auto_in_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_writealloc =
    widget_auto_in_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_privileged =
    widget_auto_in_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_secure =
    widget_auto_in_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_user_amba_prot_fetch =
    widget_auto_in_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  widget_nodeIn_a_bits_mask = widget_auto_in_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_nodeIn_a_bits_data = widget_auto_in_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_a_bits_corrupt = widget_auto_in_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_b_ready = widget_auto_in_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_nodeIn_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_nodeIn_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  widget_nodeIn_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_nodeIn_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_valid = widget_auto_in_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_c_bits_opcode = widget_auto_in_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_c_bits_param = widget_auto_in_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_c_bits_size = widget_auto_in_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_source = widget_auto_in_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_nodeIn_c_bits_address = widget_auto_in_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_bufferable =
    widget_auto_in_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_modifiable =
    widget_auto_in_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_readalloc =
    widget_auto_in_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_writealloc =
    widget_auto_in_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_privileged =
    widget_auto_in_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_secure =
    widget_auto_in_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_user_amba_prot_fetch =
    widget_auto_in_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_nodeIn_c_bits_data = widget_auto_in_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_c_bits_corrupt = widget_auto_in_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_ready = widget_auto_in_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeIn_e_valid = widget_auto_in_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_nodeIn_e_bits_sink = widget_auto_in_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_nodeOut_a_ready = widget_auto_out_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  widget_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_b_valid = widget_auto_out_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_b_bits_opcode = widget_auto_out_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_nodeOut_b_bits_param = widget_auto_out_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_nodeOut_b_bits_size = widget_auto_out_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_b_bits_source = widget_auto_out_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_nodeOut_b_bits_address = widget_auto_out_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  widget_nodeOut_b_bits_mask = widget_auto_out_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_nodeOut_b_bits_data = widget_auto_out_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_b_bits_corrupt = widget_auto_out_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_ready = widget_auto_out_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_nodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_nodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_nodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_valid = widget_auto_out_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_nodeOut_d_bits_opcode = widget_auto_out_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_nodeOut_d_bits_param = widget_auto_out_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_nodeOut_d_bits_size = widget_auto_out_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_source = widget_auto_out_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_nodeOut_d_bits_sink = widget_auto_out_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_denied = widget_auto_out_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_nodeOut_d_bits_data = widget_auto_out_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_d_bits_corrupt = widget_auto_out_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_e_ready = widget_auto_out_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_nodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_nodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_nodeIn_a_ready = widget_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_auto_out_a_valid = widget_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_opcode = widget_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_param = widget_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_size = widget_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_source = widget_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_address = widget_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_bufferable =
    widget_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_modifiable =
    widget_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_readalloc =
    widget_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_writealloc =
    widget_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_privileged =
    widget_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_secure =
    widget_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_user_amba_prot_fetch =
    widget_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_mask = widget_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_data = widget_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_a_bits_corrupt = widget_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_b_ready = widget_nodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_nodeIn_b_valid = widget_nodeOut_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_opcode = widget_nodeOut_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_param = widget_nodeOut_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_size = widget_nodeOut_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_source = widget_nodeOut_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_address = widget_nodeOut_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_mask = widget_nodeOut_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_data = widget_nodeOut_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_b_bits_corrupt = widget_nodeOut_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_c_ready = widget_nodeOut_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_auto_out_c_valid = widget_nodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_opcode = widget_nodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_param = widget_nodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_size = widget_nodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_source = widget_nodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_address = widget_nodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_bufferable =
    widget_nodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_modifiable =
    widget_nodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_readalloc =
    widget_nodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_writealloc =
    widget_nodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_privileged =
    widget_nodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_secure =
    widget_nodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_user_amba_prot_fetch =
    widget_nodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_data = widget_nodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_c_bits_corrupt = widget_nodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_d_ready = widget_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_nodeIn_d_valid = widget_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_opcode = widget_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_param = widget_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_size = widget_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_source = widget_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_sink = widget_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_denied = widget_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_data = widget_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_d_bits_corrupt = widget_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeIn_e_ready = widget_nodeOut_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_auto_out_e_valid = widget_nodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_auto_out_e_bits_sink = widget_nodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_auto_in_a_ready = widget_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_nodeOut_a_valid = widget_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_opcode = widget_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_param = widget_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_size = widget_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_source = widget_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_address = widget_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_bufferable =
    widget_nodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_modifiable =
    widget_nodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_readalloc =
    widget_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_writealloc =
    widget_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_privileged =
    widget_nodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_secure =
    widget_nodeIn_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_user_amba_prot_fetch =
    widget_nodeIn_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_mask = widget_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_data = widget_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_a_bits_corrupt = widget_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_b_ready = widget_nodeIn_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_auto_in_b_valid = widget_nodeIn_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_auto_in_b_bits_opcode = widget_nodeIn_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_auto_in_b_bits_param = widget_nodeIn_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_auto_in_b_bits_size = widget_nodeIn_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_b_bits_source = widget_nodeIn_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_auto_in_b_bits_address = widget_nodeIn_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  widget_auto_in_b_bits_mask = widget_nodeIn_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_auto_in_b_bits_data = widget_nodeIn_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_b_bits_corrupt = widget_nodeIn_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_c_ready = widget_nodeIn_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_nodeOut_c_valid = widget_nodeIn_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_opcode = widget_nodeIn_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_param = widget_nodeIn_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_size = widget_nodeIn_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_source = widget_nodeIn_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_address = widget_nodeIn_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_bufferable =
    widget_nodeIn_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_modifiable =
    widget_nodeIn_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_readalloc =
    widget_nodeIn_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_writealloc =
    widget_nodeIn_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_privileged =
    widget_nodeIn_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_secure =
    widget_nodeIn_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_user_amba_prot_fetch =
    widget_nodeIn_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_data = widget_nodeIn_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_c_bits_corrupt = widget_nodeIn_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_d_ready = widget_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        widget_auto_in_d_valid = widget_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_auto_in_d_bits_opcode = widget_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_auto_in_d_bits_param = widget_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_auto_in_d_bits_size = widget_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_d_bits_source = widget_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_auto_in_d_bits_sink = widget_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_d_bits_denied = widget_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_auto_in_d_bits_data = widget_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_d_bits_corrupt = widget_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_auto_in_e_ready = widget_nodeIn_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_nodeOut_e_valid = widget_nodeIn_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_nodeOut_e_bits_sink = widget_nodeIn_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire dcache_clock;
    wire dcache_reset;
    wire dcache_auto_out_a_ready;
    wire dcache_auto_out_a_valid;
    wire[2:0] dcache_auto_out_a_bits_opcode;
    wire[2:0] dcache_auto_out_a_bits_param;
    wire[3:0] dcache_auto_out_a_bits_size;
    wire dcache_auto_out_a_bits_source;
    wire[31:0] dcache_auto_out_a_bits_address;
    wire dcache_auto_out_a_bits_user_amba_prot_bufferable;
    wire dcache_auto_out_a_bits_user_amba_prot_modifiable;
    wire dcache_auto_out_a_bits_user_amba_prot_readalloc;
    wire dcache_auto_out_a_bits_user_amba_prot_writealloc;
    wire dcache_auto_out_a_bits_user_amba_prot_privileged;
    wire dcache_auto_out_a_bits_user_amba_prot_secure;
    wire dcache_auto_out_a_bits_user_amba_prot_fetch;
    wire[7:0] dcache_auto_out_a_bits_mask;
    wire[63:0] dcache_auto_out_a_bits_data;
    wire dcache_auto_out_a_bits_corrupt;
    wire dcache_auto_out_b_ready;
    wire dcache_auto_out_b_valid;
    wire[2:0] dcache_auto_out_b_bits_opcode;
    wire[1:0] dcache_auto_out_b_bits_param;
    wire[3:0] dcache_auto_out_b_bits_size;
    wire dcache_auto_out_b_bits_source;
    wire[31:0] dcache_auto_out_b_bits_address;
    wire[7:0] dcache_auto_out_b_bits_mask;
    wire[63:0] dcache_auto_out_b_bits_data;
    wire dcache_auto_out_b_bits_corrupt;
    wire dcache_auto_out_c_ready;
    wire dcache_auto_out_c_valid;
    wire[2:0] dcache_auto_out_c_bits_opcode;
    wire[2:0] dcache_auto_out_c_bits_param;
    wire[3:0] dcache_auto_out_c_bits_size;
    wire dcache_auto_out_c_bits_source;
    wire[31:0] dcache_auto_out_c_bits_address;
    wire dcache_auto_out_c_bits_user_amba_prot_bufferable;
    wire dcache_auto_out_c_bits_user_amba_prot_modifiable;
    wire dcache_auto_out_c_bits_user_amba_prot_readalloc;
    wire dcache_auto_out_c_bits_user_amba_prot_writealloc;
    wire dcache_auto_out_c_bits_user_amba_prot_privileged;
    wire dcache_auto_out_c_bits_user_amba_prot_secure;
    wire dcache_auto_out_c_bits_user_amba_prot_fetch;
    wire[63:0] dcache_auto_out_c_bits_data;
    wire dcache_auto_out_c_bits_corrupt;
    wire dcache_auto_out_d_ready;
    wire dcache_auto_out_d_valid;
    wire[2:0] dcache_auto_out_d_bits_opcode;
    wire[1:0] dcache_auto_out_d_bits_param;
    wire[3:0] dcache_auto_out_d_bits_size;
    wire dcache_auto_out_d_bits_source;
    wire[1:0] dcache_auto_out_d_bits_sink;
    wire dcache_auto_out_d_bits_denied;
    wire[63:0] dcache_auto_out_d_bits_data;
    wire dcache_auto_out_d_bits_corrupt;
    wire dcache_auto_out_e_ready;
    wire dcache_auto_out_e_valid;
    wire[1:0] dcache_auto_out_e_bits_sink;
    wire dcache_io_cpu_req_ready;
    wire dcache_io_cpu_req_valid;
    wire[33:0] dcache_io_cpu_req_bits_addr;
    wire[5:0] dcache_io_cpu_req_bits_tag;
    wire[4:0] dcache_io_cpu_req_bits_cmd;
    wire[1:0] dcache_io_cpu_req_bits_size;
    wire dcache_io_cpu_req_bits_signed;
    wire[1:0] dcache_io_cpu_req_bits_dprv;
    wire dcache_io_cpu_req_bits_dv;
    wire dcache_io_cpu_req_bits_phys;
    wire dcache_io_cpu_req_bits_no_alloc;
    wire dcache_io_cpu_req_bits_no_xcpt;
    wire[63:0] dcache_io_cpu_req_bits_data;
    wire[7:0] dcache_io_cpu_req_bits_mask;
    wire dcache_io_cpu_s1_kill;
    wire[63:0] dcache_io_cpu_s1_data_data;
    wire[7:0] dcache_io_cpu_s1_data_mask;
    wire dcache_io_cpu_s2_nack;
    wire dcache_io_cpu_s2_nack_cause_raw;
    wire dcache_io_cpu_s2_kill;
    wire dcache_io_cpu_s2_uncached;
    wire[31:0] dcache_io_cpu_s2_paddr;
    wire dcache_io_cpu_resp_valid;
    wire[33:0] dcache_io_cpu_resp_bits_addr;
    wire[5:0] dcache_io_cpu_resp_bits_tag;
    wire[4:0] dcache_io_cpu_resp_bits_cmd;
    wire[1:0] dcache_io_cpu_resp_bits_size;
    wire dcache_io_cpu_resp_bits_signed;
    wire[1:0] dcache_io_cpu_resp_bits_dprv;
    wire dcache_io_cpu_resp_bits_dv;
    wire[63:0] dcache_io_cpu_resp_bits_data;
    wire[7:0] dcache_io_cpu_resp_bits_mask;
    wire dcache_io_cpu_resp_bits_replay;
    wire dcache_io_cpu_resp_bits_has_data;
    wire[63:0] dcache_io_cpu_resp_bits_data_word_bypass;
    wire[63:0] dcache_io_cpu_resp_bits_data_raw;
    wire[63:0] dcache_io_cpu_resp_bits_store_data;
    wire dcache_io_cpu_replay_next;
    wire dcache_io_cpu_s2_xcpt_ma_ld;
    wire dcache_io_cpu_s2_xcpt_ma_st;
    wire dcache_io_cpu_s2_xcpt_pf_ld;
    wire dcache_io_cpu_s2_xcpt_pf_st;
    wire dcache_io_cpu_s2_xcpt_gf_ld;
    wire dcache_io_cpu_s2_xcpt_gf_st;
    wire dcache_io_cpu_s2_xcpt_ae_ld;
    wire dcache_io_cpu_s2_xcpt_ae_st;
    wire[33:0] dcache_io_cpu_s2_gpa;
    wire dcache_io_cpu_s2_gpa_is_pte;
    wire dcache_io_cpu_ordered;
    wire dcache_io_cpu_perf_acquire;
    wire dcache_io_cpu_perf_release;
    wire dcache_io_cpu_perf_grant;
    wire dcache_io_cpu_perf_tlbMiss;
    wire dcache_io_cpu_perf_blocked;
    wire dcache_io_cpu_perf_canAcceptStoreThenLoad;
    wire dcache_io_cpu_perf_canAcceptStoreThenRMW;
    wire dcache_io_cpu_perf_canAcceptLoadThenLoad;
    wire dcache_io_cpu_perf_storeBufferEmptyAfterLoad;
    wire dcache_io_cpu_perf_storeBufferEmptyAfterStore;
    wire dcache_io_cpu_keep_clock_enabled;
    wire dcache_io_cpu_clock_enabled;
    wire dcache_io_ptw_req_ready;
    wire dcache_io_ptw_req_valid;
    wire dcache_io_ptw_req_bits_valid;
    wire[20:0] dcache_io_ptw_req_bits_bits_addr;
    wire dcache_io_ptw_req_bits_bits_need_gpa;
    wire dcache_io_ptw_req_bits_bits_vstage1;
    wire dcache_io_ptw_req_bits_bits_stage2;
    wire dcache_io_ptw_resp_valid;
    wire dcache_io_ptw_resp_bits_ae_ptw;
    wire dcache_io_ptw_resp_bits_ae_final;
    wire dcache_io_ptw_resp_bits_pf;
    wire dcache_io_ptw_resp_bits_gf;
    wire dcache_io_ptw_resp_bits_hr;
    wire dcache_io_ptw_resp_bits_hw;
    wire dcache_io_ptw_resp_bits_hx;
    wire[9:0] dcache_io_ptw_resp_bits_pte_reserved_for_future;
    wire[43:0] dcache_io_ptw_resp_bits_pte_ppn;
    wire[1:0] dcache_io_ptw_resp_bits_pte_reserved_for_software;
    wire dcache_io_ptw_resp_bits_pte_d;
    wire dcache_io_ptw_resp_bits_pte_a;
    wire dcache_io_ptw_resp_bits_pte_g;
    wire dcache_io_ptw_resp_bits_pte_u;
    wire dcache_io_ptw_resp_bits_pte_x;
    wire dcache_io_ptw_resp_bits_pte_w;
    wire dcache_io_ptw_resp_bits_pte_r;
    wire dcache_io_ptw_resp_bits_pte_v;
    wire[1:0] dcache_io_ptw_resp_bits_level;
    wire dcache_io_ptw_resp_bits_fragmented_superpage;
    wire dcache_io_ptw_resp_bits_homogeneous;
    wire dcache_io_ptw_resp_bits_gpa_valid;
    wire[32:0] dcache_io_ptw_resp_bits_gpa_bits;
    wire dcache_io_ptw_resp_bits_gpa_is_pte;
    wire[3:0] dcache_io_ptw_ptbr_mode;
    wire[15:0] dcache_io_ptw_ptbr_asid;
    wire[43:0] dcache_io_ptw_ptbr_ppn;
    wire[3:0] dcache_io_ptw_hgatp_mode;
    wire[15:0] dcache_io_ptw_hgatp_asid;
    wire[43:0] dcache_io_ptw_hgatp_ppn;
    wire[3:0] dcache_io_ptw_vsatp_mode;
    wire[15:0] dcache_io_ptw_vsatp_asid;
    wire[43:0] dcache_io_ptw_vsatp_ppn;
    wire dcache_io_ptw_status_debug;
    wire dcache_io_ptw_status_cease;
    wire dcache_io_ptw_status_wfi;
    wire[31:0] dcache_io_ptw_status_isa;
    wire[1:0] dcache_io_ptw_status_dprv;
    wire dcache_io_ptw_status_dv;
    wire[1:0] dcache_io_ptw_status_prv;
    wire dcache_io_ptw_status_v;
    wire dcache_io_ptw_status_sd;
    wire[22:0] dcache_io_ptw_status_zero2;
    wire dcache_io_ptw_status_mpv;
    wire dcache_io_ptw_status_gva;
    wire dcache_io_ptw_status_mbe;
    wire dcache_io_ptw_status_sbe;
    wire[1:0] dcache_io_ptw_status_sxl;
    wire[1:0] dcache_io_ptw_status_uxl;
    wire dcache_io_ptw_status_sd_rv32;
    wire[7:0] dcache_io_ptw_status_zero1;
    wire dcache_io_ptw_status_tsr;
    wire dcache_io_ptw_status_tw;
    wire dcache_io_ptw_status_tvm;
    wire dcache_io_ptw_status_mxr;
    wire dcache_io_ptw_status_sum;
    wire dcache_io_ptw_status_mprv;
    wire[1:0] dcache_io_ptw_status_xs;
    wire[1:0] dcache_io_ptw_status_fs;
    wire[1:0] dcache_io_ptw_status_mpp;
    wire[1:0] dcache_io_ptw_status_vs;
    wire dcache_io_ptw_status_spp;
    wire dcache_io_ptw_status_mpie;
    wire dcache_io_ptw_status_ube;
    wire dcache_io_ptw_status_spie;
    wire dcache_io_ptw_status_upie;
    wire dcache_io_ptw_status_mie;
    wire dcache_io_ptw_status_hie;
    wire dcache_io_ptw_status_sie;
    wire dcache_io_ptw_status_uie;
    wire[29:0] dcache_io_ptw_hstatus_zero6;
    wire[1:0] dcache_io_ptw_hstatus_vsxl;
    wire[8:0] dcache_io_ptw_hstatus_zero5;
    wire dcache_io_ptw_hstatus_vtsr;
    wire dcache_io_ptw_hstatus_vtw;
    wire dcache_io_ptw_hstatus_vtvm;
    wire[1:0] dcache_io_ptw_hstatus_zero3;
    wire[5:0] dcache_io_ptw_hstatus_vgein;
    wire[1:0] dcache_io_ptw_hstatus_zero2;
    wire dcache_io_ptw_hstatus_hu;
    wire dcache_io_ptw_hstatus_spvp;
    wire dcache_io_ptw_hstatus_spv;
    wire dcache_io_ptw_hstatus_gva;
    wire dcache_io_ptw_hstatus_vsbe;
    wire[4:0] dcache_io_ptw_hstatus_zero1;
    wire dcache_io_ptw_gstatus_debug;
    wire dcache_io_ptw_gstatus_cease;
    wire dcache_io_ptw_gstatus_wfi;
    wire[31:0] dcache_io_ptw_gstatus_isa;
    wire[1:0] dcache_io_ptw_gstatus_dprv;
    wire dcache_io_ptw_gstatus_dv;
    wire[1:0] dcache_io_ptw_gstatus_prv;
    wire dcache_io_ptw_gstatus_v;
    wire dcache_io_ptw_gstatus_sd;
    wire[22:0] dcache_io_ptw_gstatus_zero2;
    wire dcache_io_ptw_gstatus_mpv;
    wire dcache_io_ptw_gstatus_gva;
    wire dcache_io_ptw_gstatus_mbe;
    wire dcache_io_ptw_gstatus_sbe;
    wire[1:0] dcache_io_ptw_gstatus_sxl;
    wire[1:0] dcache_io_ptw_gstatus_uxl;
    wire dcache_io_ptw_gstatus_sd_rv32;
    wire[7:0] dcache_io_ptw_gstatus_zero1;
    wire dcache_io_ptw_gstatus_tsr;
    wire dcache_io_ptw_gstatus_tw;
    wire dcache_io_ptw_gstatus_tvm;
    wire dcache_io_ptw_gstatus_mxr;
    wire dcache_io_ptw_gstatus_sum;
    wire dcache_io_ptw_gstatus_mprv;
    wire[1:0] dcache_io_ptw_gstatus_xs;
    wire[1:0] dcache_io_ptw_gstatus_fs;
    wire[1:0] dcache_io_ptw_gstatus_mpp;
    wire[1:0] dcache_io_ptw_gstatus_vs;
    wire dcache_io_ptw_gstatus_spp;
    wire dcache_io_ptw_gstatus_mpie;
    wire dcache_io_ptw_gstatus_ube;
    wire dcache_io_ptw_gstatus_spie;
    wire dcache_io_ptw_gstatus_upie;
    wire dcache_io_ptw_gstatus_mie;
    wire dcache_io_ptw_gstatus_hie;
    wire dcache_io_ptw_gstatus_sie;
    wire dcache_io_ptw_gstatus_uie;
    wire dcache_io_ptw_pmp_0_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_0_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_0_cfg_a;
    wire dcache_io_ptw_pmp_0_cfg_x;
    wire dcache_io_ptw_pmp_0_cfg_w;
    wire dcache_io_ptw_pmp_0_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_0_addr;
    wire[31:0] dcache_io_ptw_pmp_0_mask;
    wire dcache_io_ptw_pmp_1_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_1_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_1_cfg_a;
    wire dcache_io_ptw_pmp_1_cfg_x;
    wire dcache_io_ptw_pmp_1_cfg_w;
    wire dcache_io_ptw_pmp_1_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_1_addr;
    wire[31:0] dcache_io_ptw_pmp_1_mask;
    wire dcache_io_ptw_pmp_2_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_2_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_2_cfg_a;
    wire dcache_io_ptw_pmp_2_cfg_x;
    wire dcache_io_ptw_pmp_2_cfg_w;
    wire dcache_io_ptw_pmp_2_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_2_addr;
    wire[31:0] dcache_io_ptw_pmp_2_mask;
    wire dcache_io_ptw_pmp_3_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_3_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_3_cfg_a;
    wire dcache_io_ptw_pmp_3_cfg_x;
    wire dcache_io_ptw_pmp_3_cfg_w;
    wire dcache_io_ptw_pmp_3_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_3_addr;
    wire[31:0] dcache_io_ptw_pmp_3_mask;
    wire dcache_io_ptw_pmp_4_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_4_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_4_cfg_a;
    wire dcache_io_ptw_pmp_4_cfg_x;
    wire dcache_io_ptw_pmp_4_cfg_w;
    wire dcache_io_ptw_pmp_4_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_4_addr;
    wire[31:0] dcache_io_ptw_pmp_4_mask;
    wire dcache_io_ptw_pmp_5_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_5_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_5_cfg_a;
    wire dcache_io_ptw_pmp_5_cfg_x;
    wire dcache_io_ptw_pmp_5_cfg_w;
    wire dcache_io_ptw_pmp_5_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_5_addr;
    wire[31:0] dcache_io_ptw_pmp_5_mask;
    wire dcache_io_ptw_pmp_6_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_6_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_6_cfg_a;
    wire dcache_io_ptw_pmp_6_cfg_x;
    wire dcache_io_ptw_pmp_6_cfg_w;
    wire dcache_io_ptw_pmp_6_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_6_addr;
    wire[31:0] dcache_io_ptw_pmp_6_mask;
    wire dcache_io_ptw_pmp_7_cfg_l;
    wire[1:0] dcache_io_ptw_pmp_7_cfg_res;
    wire[1:0] dcache_io_ptw_pmp_7_cfg_a;
    wire dcache_io_ptw_pmp_7_cfg_x;
    wire dcache_io_ptw_pmp_7_cfg_w;
    wire dcache_io_ptw_pmp_7_cfg_r;
    wire[29:0] dcache_io_ptw_pmp_7_addr;
    wire[31:0] dcache_io_ptw_pmp_7_mask;
    wire dcache_io_ptw_customCSRs_csrs_0_ren;
    wire dcache_io_ptw_customCSRs_csrs_0_wen;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_0_wdata;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_0_value;
    wire dcache_io_ptw_customCSRs_csrs_0_stall;
    wire dcache_io_ptw_customCSRs_csrs_0_set;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_0_sdata;
    wire dcache_io_ptw_customCSRs_csrs_1_ren;
    wire dcache_io_ptw_customCSRs_csrs_1_wen;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_1_wdata;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_1_value;
    wire dcache_io_ptw_customCSRs_csrs_1_stall;
    wire dcache_io_ptw_customCSRs_csrs_1_set;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_1_sdata;
    wire dcache_io_ptw_customCSRs_csrs_2_ren;
    wire dcache_io_ptw_customCSRs_csrs_2_wen;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_2_wdata;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_2_value;
    wire dcache_io_ptw_customCSRs_csrs_2_stall;
    wire dcache_io_ptw_customCSRs_csrs_2_set;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_2_sdata;
    wire dcache_io_ptw_customCSRs_csrs_3_ren;
    wire dcache_io_ptw_customCSRs_csrs_3_wen;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_3_wdata;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_3_value;
    wire dcache_io_ptw_customCSRs_csrs_3_stall;
    wire dcache_io_ptw_customCSRs_csrs_3_set;
    wire[63:0] dcache_io_ptw_customCSRs_csrs_3_sdata;
    wire dcache_io_errors_bus_valid;
    wire[31:0] dcache_io_errors_bus_bits;
    wire dcache_tlb_port_req_ready;
    wire dcache_tlb_port_req_valid;
    wire[33:0] dcache_tlb_port_req_bits_vaddr;
    wire dcache_tlb_port_req_bits_passthrough;
    wire[1:0] dcache_tlb_port_req_bits_size;
    wire[4:0] dcache_tlb_port_req_bits_cmd;
    wire[1:0] dcache_tlb_port_req_bits_prv;
    wire dcache_tlb_port_req_bits_v;
    wire dcache_tlb_port_s1_resp_miss;
    wire[31:0] dcache_tlb_port_s1_resp_paddr;
    wire[33:0] dcache_tlb_port_s1_resp_gpa;
    wire dcache_tlb_port_s1_resp_gpa_is_pte;
    wire dcache_tlb_port_s1_resp_pf_ld;
    wire dcache_tlb_port_s1_resp_pf_st;
    wire dcache_tlb_port_s1_resp_pf_inst;
    wire dcache_tlb_port_s1_resp_gf_ld;
    wire dcache_tlb_port_s1_resp_gf_st;
    wire dcache_tlb_port_s1_resp_gf_inst;
    wire dcache_tlb_port_s1_resp_ae_ld;
    wire dcache_tlb_port_s1_resp_ae_st;
    wire dcache_tlb_port_s1_resp_ae_inst;
    wire dcache_tlb_port_s1_resp_ma_ld;
    wire dcache_tlb_port_s1_resp_ma_st;
    wire dcache_tlb_port_s1_resp_ma_inst;
    wire dcache_tlb_port_s1_resp_cacheable;
    wire dcache_tlb_port_s1_resp_must_alloc;
    wire dcache_tlb_port_s1_resp_prefetchable;
    wire dcache_tlb_port_s2_kill;

    wire[1:0] dcache_newCoh_state ; 
    wire[19:0] dcache_s2_meta_corrected_0_tag ; 
    wire dcache_tl_out_a_bits_corrupt ; 
    wire[63:0] dcache_tl_out_a_bits_data ; 
    wire[7:0] dcache_tl_out_a_bits_mask ; 
    wire dcache_tl_out_a_bits_user_amba_prot_privileged ; 
    wire dcache_tl_out_a_bits_user_amba_prot_writealloc ; 
    wire dcache_tl_out_a_bits_user_amba_prot_readalloc ; 
    wire dcache_tl_out_a_bits_user_amba_prot_modifiable ; 
    wire dcache_tl_out_a_bits_user_amba_prot_bufferable ; 
    wire[31:0] dcache_tl_out_a_bits_address ; 
    wire dcache_tl_out_a_bits_source ; 
    wire[3:0] dcache_tl_out_a_bits_size ; 
    wire[2:0] dcache_tl_out_a_bits_param ; 
    wire[2:0] dcache_tl_out_a_bits_opcode ; 
    wire dcache_tl_out_a_valid ; 
    wire[63:0] dcache_dataArb_io_in_1_bits_wdata ; 
    wire[63:0] dcache_s1_all_data_ways_0 ; 
    wire dcache__GEN ; 
    wire[21:0] dcache_tag_array_s1_meta_data_0 ; 
    wire[21:0] dcache_metaArb_io_out_bits_data ; 
    wire[5:0] dcache_metaArb_io_out_bits_idx ; 
    wire[21:0] dcache_metaArb_io_in_4_bits_data ; 
    wire dcache_metaArb_io_in_4_bits_way_en ; 
    wire[1:0] dcache__pma_checker_mpu_priv_1to0 ; 
    wire[31:0] dcache__pma_checker_mpu_physaddr_31to0 ; 
    wire[1:0] dcache__tlb_mpu_priv_1to0 ; 
    wire[31:0] dcache__tlb_mpu_physaddr_31to0 ; 
    wire dcache__lfsr_prng_io_out_0 ; 
    wire dcache__lfsr_prng_io_out_1 ; 
    wire dcache__lfsr_prng_io_out_2 ; 
    wire dcache__lfsr_prng_io_out_3 ; 
    wire dcache__lfsr_prng_io_out_4 ; 
    wire dcache__lfsr_prng_io_out_5 ; 
    wire dcache__lfsr_prng_io_out_6 ; 
    wire dcache__lfsr_prng_io_out_7 ; 
    wire dcache__lfsr_prng_io_out_8 ; 
    wire dcache__lfsr_prng_io_out_9 ; 
    wire dcache__lfsr_prng_io_out_10 ; 
    wire dcache__lfsr_prng_io_out_11 ; 
    wire dcache__lfsr_prng_io_out_12 ; 
    wire dcache__lfsr_prng_io_out_13 ; 
    wire dcache__lfsr_prng_io_out_14 ; 
    wire dcache__lfsr_prng_io_out_15 ; 
    wire[19:0] dcache__pma_checker_entries_barrier_5_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_5_io_y_hr ; 
    wire[19:0] dcache__pma_checker_entries_barrier_4_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_4_io_y_c ; 
    wire[19:0] dcache__pma_checker_entries_barrier_3_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_3_io_y_c ; 
    wire[19:0] dcache__pma_checker_entries_barrier_2_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_2_io_y_c ; 
    wire[19:0] dcache__pma_checker_entries_barrier_1_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_1_io_y_c ; 
    wire[19:0] dcache__pma_checker_entries_barrier_io_y_ppn ; 
    wire dcache__pma_checker_entries_barrier_io_y_u ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_ptw ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_final ; 
    wire dcache__pma_checker_entries_barrier_io_y_ae_stage2 ; 
    wire dcache__pma_checker_entries_barrier_io_y_pf ; 
    wire dcache__pma_checker_entries_barrier_io_y_gf ; 
    wire dcache__pma_checker_entries_barrier_io_y_sw ; 
    wire dcache__pma_checker_entries_barrier_io_y_sx ; 
    wire dcache__pma_checker_entries_barrier_io_y_sr ; 
    wire dcache__pma_checker_entries_barrier_io_y_hw ; 
    wire dcache__pma_checker_entries_barrier_io_y_hx ; 
    wire dcache__pma_checker_entries_barrier_io_y_hr ; 
    wire dcache__pma_checker_entries_barrier_io_y_pw ; 
    wire dcache__pma_checker_entries_barrier_io_y_px ; 
    wire dcache__pma_checker_entries_barrier_io_y_pr ; 
    wire dcache__pma_checker_entries_barrier_io_y_ppp ; 
    wire dcache__pma_checker_entries_barrier_io_y_pal ; 
    wire dcache__pma_checker_entries_barrier_io_y_paa ; 
    wire dcache__pma_checker_entries_barrier_io_y_eff ; 
    wire dcache__pma_checker_entries_barrier_io_y_c ; 
    wire dcache__pma_checker_pmp_io_r ; 
    wire dcache__pma_checker_pmp_io_w ; 
    wire dcache__pma_checker_pmp_io_x ; 
    wire[19:0] dcache__pma_checker_mpu_ppn_barrier_io_y_ppn ; 
    wire[19:0] dcache__tlb_entries_barrier_5_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_5_io_y_u ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_5_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_5_io_y_pf ; 
    wire dcache__tlb_entries_barrier_5_io_y_gf ; 
    wire dcache__tlb_entries_barrier_5_io_y_sw ; 
    wire dcache__tlb_entries_barrier_5_io_y_sx ; 
    wire dcache__tlb_entries_barrier_5_io_y_sr ; 
    wire dcache__tlb_entries_barrier_5_io_y_hw ; 
    wire dcache__tlb_entries_barrier_5_io_y_hx ; 
    wire dcache__tlb_entries_barrier_5_io_y_hr ; 
    wire[19:0] dcache__tlb_entries_barrier_4_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_4_io_y_u ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_4_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_4_io_y_pf ; 
    wire dcache__tlb_entries_barrier_4_io_y_gf ; 
    wire dcache__tlb_entries_barrier_4_io_y_sw ; 
    wire dcache__tlb_entries_barrier_4_io_y_sx ; 
    wire dcache__tlb_entries_barrier_4_io_y_sr ; 
    wire dcache__tlb_entries_barrier_4_io_y_hw ; 
    wire dcache__tlb_entries_barrier_4_io_y_hx ; 
    wire dcache__tlb_entries_barrier_4_io_y_hr ; 
    wire dcache__tlb_entries_barrier_4_io_y_pw ; 
    wire dcache__tlb_entries_barrier_4_io_y_px ; 
    wire dcache__tlb_entries_barrier_4_io_y_pr ; 
    wire dcache__tlb_entries_barrier_4_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_4_io_y_pal ; 
    wire dcache__tlb_entries_barrier_4_io_y_paa ; 
    wire dcache__tlb_entries_barrier_4_io_y_eff ; 
    wire dcache__tlb_entries_barrier_4_io_y_c ; 
    wire[19:0] dcache__tlb_entries_barrier_3_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_3_io_y_u ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_3_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_3_io_y_pf ; 
    wire dcache__tlb_entries_barrier_3_io_y_gf ; 
    wire dcache__tlb_entries_barrier_3_io_y_sw ; 
    wire dcache__tlb_entries_barrier_3_io_y_sx ; 
    wire dcache__tlb_entries_barrier_3_io_y_sr ; 
    wire dcache__tlb_entries_barrier_3_io_y_hw ; 
    wire dcache__tlb_entries_barrier_3_io_y_hx ; 
    wire dcache__tlb_entries_barrier_3_io_y_hr ; 
    wire dcache__tlb_entries_barrier_3_io_y_pw ; 
    wire dcache__tlb_entries_barrier_3_io_y_px ; 
    wire dcache__tlb_entries_barrier_3_io_y_pr ; 
    wire dcache__tlb_entries_barrier_3_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_3_io_y_pal ; 
    wire dcache__tlb_entries_barrier_3_io_y_paa ; 
    wire dcache__tlb_entries_barrier_3_io_y_eff ; 
    wire dcache__tlb_entries_barrier_3_io_y_c ; 
    wire[19:0] dcache__tlb_entries_barrier_2_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_2_io_y_u ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_2_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_2_io_y_pf ; 
    wire dcache__tlb_entries_barrier_2_io_y_gf ; 
    wire dcache__tlb_entries_barrier_2_io_y_sw ; 
    wire dcache__tlb_entries_barrier_2_io_y_sx ; 
    wire dcache__tlb_entries_barrier_2_io_y_sr ; 
    wire dcache__tlb_entries_barrier_2_io_y_hw ; 
    wire dcache__tlb_entries_barrier_2_io_y_hx ; 
    wire dcache__tlb_entries_barrier_2_io_y_hr ; 
    wire dcache__tlb_entries_barrier_2_io_y_pw ; 
    wire dcache__tlb_entries_barrier_2_io_y_px ; 
    wire dcache__tlb_entries_barrier_2_io_y_pr ; 
    wire dcache__tlb_entries_barrier_2_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_2_io_y_pal ; 
    wire dcache__tlb_entries_barrier_2_io_y_paa ; 
    wire dcache__tlb_entries_barrier_2_io_y_eff ; 
    wire dcache__tlb_entries_barrier_2_io_y_c ; 
    wire[19:0] dcache__tlb_entries_barrier_1_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_1_io_y_u ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_1_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_1_io_y_pf ; 
    wire dcache__tlb_entries_barrier_1_io_y_gf ; 
    wire dcache__tlb_entries_barrier_1_io_y_sw ; 
    wire dcache__tlb_entries_barrier_1_io_y_sx ; 
    wire dcache__tlb_entries_barrier_1_io_y_sr ; 
    wire dcache__tlb_entries_barrier_1_io_y_hw ; 
    wire dcache__tlb_entries_barrier_1_io_y_hx ; 
    wire dcache__tlb_entries_barrier_1_io_y_hr ; 
    wire dcache__tlb_entries_barrier_1_io_y_pw ; 
    wire dcache__tlb_entries_barrier_1_io_y_px ; 
    wire dcache__tlb_entries_barrier_1_io_y_pr ; 
    wire dcache__tlb_entries_barrier_1_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_1_io_y_pal ; 
    wire dcache__tlb_entries_barrier_1_io_y_paa ; 
    wire dcache__tlb_entries_barrier_1_io_y_eff ; 
    wire dcache__tlb_entries_barrier_1_io_y_c ; 
    wire[19:0] dcache__tlb_entries_barrier_io_y_ppn ; 
    wire dcache__tlb_entries_barrier_io_y_u ; 
    wire dcache__tlb_entries_barrier_io_y_ae_ptw ; 
    wire dcache__tlb_entries_barrier_io_y_ae_final ; 
    wire dcache__tlb_entries_barrier_io_y_ae_stage2 ; 
    wire dcache__tlb_entries_barrier_io_y_pf ; 
    wire dcache__tlb_entries_barrier_io_y_gf ; 
    wire dcache__tlb_entries_barrier_io_y_sw ; 
    wire dcache__tlb_entries_barrier_io_y_sx ; 
    wire dcache__tlb_entries_barrier_io_y_sr ; 
    wire dcache__tlb_entries_barrier_io_y_hw ; 
    wire dcache__tlb_entries_barrier_io_y_hx ; 
    wire dcache__tlb_entries_barrier_io_y_hr ; 
    wire dcache__tlb_entries_barrier_io_y_pw ; 
    wire dcache__tlb_entries_barrier_io_y_px ; 
    wire dcache__tlb_entries_barrier_io_y_pr ; 
    wire dcache__tlb_entries_barrier_io_y_ppp ; 
    wire dcache__tlb_entries_barrier_io_y_pal ; 
    wire dcache__tlb_entries_barrier_io_y_paa ; 
    wire dcache__tlb_entries_barrier_io_y_eff ; 
    wire dcache__tlb_entries_barrier_io_y_c ; 
    wire dcache__tlb_pmp_io_r ; 
    wire dcache__tlb_pmp_io_w ; 
    wire dcache__tlb_pmp_io_x ; 
    wire[19:0] dcache__tlb_mpu_ppn_barrier_io_y_ppn ; 
    wire dcache_nodeOut_a_ready = dcache_auto_out_a_ready ; 
    wire dcache_nodeOut_b_valid = dcache_auto_out_b_valid ; 
    wire[2:0] dcache_nodeOut_b_bits_opcode = dcache_auto_out_b_bits_opcode ; 
    wire[1:0] dcache_nodeOut_b_bits_param = dcache_auto_out_b_bits_param ; 
    wire[3:0] dcache_nodeOut_b_bits_size = dcache_auto_out_b_bits_size ; 
    wire dcache_nodeOut_b_bits_source = dcache_auto_out_b_bits_source ; 
    wire[31:0] dcache_nodeOut_b_bits_address = dcache_auto_out_b_bits_address ; 
    wire[7:0] dcache_nodeOut_b_bits_mask = dcache_auto_out_b_bits_mask ; 
    wire[63:0] dcache_nodeOut_b_bits_data = dcache_auto_out_b_bits_data ; 
    wire dcache_nodeOut_b_bits_corrupt = dcache_auto_out_b_bits_corrupt ; 
    wire dcache_nodeOut_c_ready = dcache_auto_out_c_ready ; 
    wire dcache_nodeOut_d_valid = dcache_auto_out_d_valid ; 
    wire[2:0] dcache_nodeOut_d_bits_opcode = dcache_auto_out_d_bits_opcode ; 
    wire[1:0] dcache_nodeOut_d_bits_param = dcache_auto_out_d_bits_param ; 
    wire[3:0] dcache_nodeOut_d_bits_size = dcache_auto_out_d_bits_size ; 
    wire dcache_nodeOut_d_bits_source = dcache_auto_out_d_bits_source ; 
    wire[1:0] dcache_nodeOut_d_bits_sink = dcache_auto_out_d_bits_sink ; 
    wire dcache_nodeOut_d_bits_denied = dcache_auto_out_d_bits_denied ; 
    wire[63:0] dcache_nodeOut_d_bits_data = dcache_auto_out_d_bits_data ; 
    wire dcache_nodeOut_d_bits_corrupt = dcache_auto_out_d_bits_corrupt ; 
    wire dcache_nodeOut_e_ready = dcache_auto_out_e_ready ; 
    wire dcache_tlb_clock = dcache_clock ; 
    wire dcache_tlb_reset = dcache_reset ; 
    wire dcache_tlb_io_ptw_req_ready = dcache_io_ptw_req_ready ; 
    wire dcache_tlb_io_ptw_resp_valid = dcache_io_ptw_resp_valid ; 
    wire dcache_tlb_io_ptw_resp_bits_ae_ptw = dcache_io_ptw_resp_bits_ae_ptw ; 
    wire dcache_tlb_io_ptw_resp_bits_ae_final = dcache_io_ptw_resp_bits_ae_final ; 
    wire dcache_tlb_io_ptw_resp_bits_pf = dcache_io_ptw_resp_bits_pf ; 
    wire dcache_tlb_io_ptw_resp_bits_gf = dcache_io_ptw_resp_bits_gf ; 
    wire dcache_tlb_io_ptw_resp_bits_hr = dcache_io_ptw_resp_bits_hr ; 
    wire dcache_tlb_io_ptw_resp_bits_hw = dcache_io_ptw_resp_bits_hw ; 
    wire dcache_tlb_io_ptw_resp_bits_hx = dcache_io_ptw_resp_bits_hx ; 
    wire[9:0] dcache_tlb_io_ptw_resp_bits_pte_reserved_for_future = dcache_io_ptw_resp_bits_pte_reserved_for_future ; 
    wire[43:0] dcache_tlb_io_ptw_resp_bits_pte_ppn = dcache_io_ptw_resp_bits_pte_ppn ; 
    wire[1:0] dcache_tlb_io_ptw_resp_bits_pte_reserved_for_software = dcache_io_ptw_resp_bits_pte_reserved_for_software ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_d = dcache_io_ptw_resp_bits_pte_d ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_a = dcache_io_ptw_resp_bits_pte_a ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_g = dcache_io_ptw_resp_bits_pte_g ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_u = dcache_io_ptw_resp_bits_pte_u ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_x = dcache_io_ptw_resp_bits_pte_x ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_w = dcache_io_ptw_resp_bits_pte_w ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_r = dcache_io_ptw_resp_bits_pte_r ; 
    wire dcache_tlb_io_ptw_resp_bits_pte_v = dcache_io_ptw_resp_bits_pte_v ; 
    wire[1:0] dcache_tlb_io_ptw_resp_bits_level = dcache_io_ptw_resp_bits_level ; 
    wire dcache_tlb_io_ptw_resp_bits_fragmented_superpage = dcache_io_ptw_resp_bits_fragmented_superpage ; 
    wire dcache_tlb_io_ptw_resp_bits_homogeneous = dcache_io_ptw_resp_bits_homogeneous ; 
    wire dcache_tlb_io_ptw_resp_bits_gpa_valid = dcache_io_ptw_resp_bits_gpa_valid ; 
    wire[32:0] dcache_tlb_io_ptw_resp_bits_gpa_bits = dcache_io_ptw_resp_bits_gpa_bits ; 
    wire dcache_tlb_io_ptw_resp_bits_gpa_is_pte = dcache_io_ptw_resp_bits_gpa_is_pte ; 
    wire[3:0] dcache_tlb_io_ptw_ptbr_mode = dcache_io_ptw_ptbr_mode ; 
    wire[15:0] dcache_tlb_io_ptw_ptbr_asid = dcache_io_ptw_ptbr_asid ; 
    wire[43:0] dcache_tlb_io_ptw_ptbr_ppn = dcache_io_ptw_ptbr_ppn ; 
    wire[3:0] dcache_tlb_io_ptw_hgatp_mode = dcache_io_ptw_hgatp_mode ; 
    wire[15:0] dcache_tlb_io_ptw_hgatp_asid = dcache_io_ptw_hgatp_asid ; 
    wire[43:0] dcache_tlb_io_ptw_hgatp_ppn = dcache_io_ptw_hgatp_ppn ; 
    wire[3:0] dcache_tlb_io_ptw_vsatp_mode = dcache_io_ptw_vsatp_mode ; 
    wire[15:0] dcache_tlb_io_ptw_vsatp_asid = dcache_io_ptw_vsatp_asid ; 
    wire[43:0] dcache_tlb_io_ptw_vsatp_ppn = dcache_io_ptw_vsatp_ppn ; 
    wire dcache_tlb_io_ptw_status_debug = dcache_io_ptw_status_debug ; 
    wire dcache_tlb_io_ptw_status_cease = dcache_io_ptw_status_cease ; 
    wire dcache_tlb_io_ptw_status_wfi = dcache_io_ptw_status_wfi ; 
    wire[31:0] dcache_tlb_io_ptw_status_isa = dcache_io_ptw_status_isa ; 
    wire[1:0] dcache_tlb_io_ptw_status_dprv = dcache_io_ptw_status_dprv ; 
    wire dcache_tlb_io_ptw_status_dv = dcache_io_ptw_status_dv ; 
    wire[1:0] dcache_tlb_io_ptw_status_prv = dcache_io_ptw_status_prv ; 
    wire dcache_tlb_io_ptw_status_v = dcache_io_ptw_status_v ; 
    wire dcache_tlb_io_ptw_status_sd = dcache_io_ptw_status_sd ; 
    wire[22:0] dcache_tlb_io_ptw_status_zero2 = dcache_io_ptw_status_zero2 ; 
    wire dcache_tlb_io_ptw_status_mpv = dcache_io_ptw_status_mpv ; 
    wire dcache_tlb_io_ptw_status_gva = dcache_io_ptw_status_gva ; 
    wire dcache_tlb_io_ptw_status_mbe = dcache_io_ptw_status_mbe ; 
    wire dcache_tlb_io_ptw_status_sbe = dcache_io_ptw_status_sbe ; 
    wire[1:0] dcache_tlb_io_ptw_status_sxl = dcache_io_ptw_status_sxl ; 
    wire[1:0] dcache_tlb_io_ptw_status_uxl = dcache_io_ptw_status_uxl ; 
    wire dcache_tlb_io_ptw_status_sd_rv32 = dcache_io_ptw_status_sd_rv32 ; 
    wire[7:0] dcache_tlb_io_ptw_status_zero1 = dcache_io_ptw_status_zero1 ; 
    wire dcache_tlb_io_ptw_status_tsr = dcache_io_ptw_status_tsr ; 
    wire dcache_tlb_io_ptw_status_tw = dcache_io_ptw_status_tw ; 
    wire dcache_tlb_io_ptw_status_tvm = dcache_io_ptw_status_tvm ; 
    wire dcache_tlb_io_ptw_status_mxr = dcache_io_ptw_status_mxr ; 
    wire dcache_tlb_io_ptw_status_sum = dcache_io_ptw_status_sum ; 
    wire dcache_tlb_io_ptw_status_mprv = dcache_io_ptw_status_mprv ; 
    wire[1:0] dcache_tlb_io_ptw_status_xs = dcache_io_ptw_status_xs ; 
    wire[1:0] dcache_tlb_io_ptw_status_fs = dcache_io_ptw_status_fs ; 
    wire[1:0] dcache_tlb_io_ptw_status_mpp = dcache_io_ptw_status_mpp ; 
    wire[1:0] dcache_tlb_io_ptw_status_vs = dcache_io_ptw_status_vs ; 
    wire dcache_tlb_io_ptw_status_spp = dcache_io_ptw_status_spp ; 
    wire dcache_tlb_io_ptw_status_mpie = dcache_io_ptw_status_mpie ; 
    wire dcache_tlb_io_ptw_status_ube = dcache_io_ptw_status_ube ; 
    wire dcache_tlb_io_ptw_status_spie = dcache_io_ptw_status_spie ; 
    wire dcache_tlb_io_ptw_status_upie = dcache_io_ptw_status_upie ; 
    wire dcache_tlb_io_ptw_status_mie = dcache_io_ptw_status_mie ; 
    wire dcache_tlb_io_ptw_status_hie = dcache_io_ptw_status_hie ; 
    wire dcache_tlb_io_ptw_status_sie = dcache_io_ptw_status_sie ; 
    wire dcache_tlb_io_ptw_status_uie = dcache_io_ptw_status_uie ; 
    wire[29:0] dcache_tlb_io_ptw_hstatus_zero6 = dcache_io_ptw_hstatus_zero6 ; 
    wire[1:0] dcache_tlb_io_ptw_hstatus_vsxl = dcache_io_ptw_hstatus_vsxl ; 
    wire[8:0] dcache_tlb_io_ptw_hstatus_zero5 = dcache_io_ptw_hstatus_zero5 ; 
    wire dcache_tlb_io_ptw_hstatus_vtsr = dcache_io_ptw_hstatus_vtsr ; 
    wire dcache_tlb_io_ptw_hstatus_vtw = dcache_io_ptw_hstatus_vtw ; 
    wire dcache_tlb_io_ptw_hstatus_vtvm = dcache_io_ptw_hstatus_vtvm ; 
    wire[1:0] dcache_tlb_io_ptw_hstatus_zero3 = dcache_io_ptw_hstatus_zero3 ; 
    wire[5:0] dcache_tlb_io_ptw_hstatus_vgein = dcache_io_ptw_hstatus_vgein ; 
    wire[1:0] dcache_tlb_io_ptw_hstatus_zero2 = dcache_io_ptw_hstatus_zero2 ; 
    wire dcache_tlb_io_ptw_hstatus_hu = dcache_io_ptw_hstatus_hu ; 
    wire dcache_tlb_io_ptw_hstatus_spvp = dcache_io_ptw_hstatus_spvp ; 
    wire dcache_tlb_io_ptw_hstatus_spv = dcache_io_ptw_hstatus_spv ; 
    wire dcache_tlb_io_ptw_hstatus_gva = dcache_io_ptw_hstatus_gva ; 
    wire dcache_tlb_io_ptw_hstatus_vsbe = dcache_io_ptw_hstatus_vsbe ; 
    wire[4:0] dcache_tlb_io_ptw_hstatus_zero1 = dcache_io_ptw_hstatus_zero1 ; 
    wire dcache_tlb_io_ptw_gstatus_debug = dcache_io_ptw_gstatus_debug ; 
    wire dcache_tlb_io_ptw_gstatus_cease = dcache_io_ptw_gstatus_cease ; 
    wire dcache_tlb_io_ptw_gstatus_wfi = dcache_io_ptw_gstatus_wfi ; 
    wire[31:0] dcache_tlb_io_ptw_gstatus_isa = dcache_io_ptw_gstatus_isa ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_dprv = dcache_io_ptw_gstatus_dprv ; 
    wire dcache_tlb_io_ptw_gstatus_dv = dcache_io_ptw_gstatus_dv ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_prv = dcache_io_ptw_gstatus_prv ; 
    wire dcache_tlb_io_ptw_gstatus_v = dcache_io_ptw_gstatus_v ; 
    wire dcache_tlb_io_ptw_gstatus_sd = dcache_io_ptw_gstatus_sd ; 
    wire[22:0] dcache_tlb_io_ptw_gstatus_zero2 = dcache_io_ptw_gstatus_zero2 ; 
    wire dcache_tlb_io_ptw_gstatus_mpv = dcache_io_ptw_gstatus_mpv ; 
    wire dcache_tlb_io_ptw_gstatus_gva = dcache_io_ptw_gstatus_gva ; 
    wire dcache_tlb_io_ptw_gstatus_mbe = dcache_io_ptw_gstatus_mbe ; 
    wire dcache_tlb_io_ptw_gstatus_sbe = dcache_io_ptw_gstatus_sbe ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_sxl = dcache_io_ptw_gstatus_sxl ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_uxl = dcache_io_ptw_gstatus_uxl ; 
    wire dcache_tlb_io_ptw_gstatus_sd_rv32 = dcache_io_ptw_gstatus_sd_rv32 ; 
    wire[7:0] dcache_tlb_io_ptw_gstatus_zero1 = dcache_io_ptw_gstatus_zero1 ; 
    wire dcache_tlb_io_ptw_gstatus_tsr = dcache_io_ptw_gstatus_tsr ; 
    wire dcache_tlb_io_ptw_gstatus_tw = dcache_io_ptw_gstatus_tw ; 
    wire dcache_tlb_io_ptw_gstatus_tvm = dcache_io_ptw_gstatus_tvm ; 
    wire dcache_tlb_io_ptw_gstatus_mxr = dcache_io_ptw_gstatus_mxr ; 
    wire dcache_tlb_io_ptw_gstatus_sum = dcache_io_ptw_gstatus_sum ; 
    wire dcache_tlb_io_ptw_gstatus_mprv = dcache_io_ptw_gstatus_mprv ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_xs = dcache_io_ptw_gstatus_xs ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_fs = dcache_io_ptw_gstatus_fs ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_mpp = dcache_io_ptw_gstatus_mpp ; 
    wire[1:0] dcache_tlb_io_ptw_gstatus_vs = dcache_io_ptw_gstatus_vs ; 
    wire dcache_tlb_io_ptw_gstatus_spp = dcache_io_ptw_gstatus_spp ; 
    wire dcache_tlb_io_ptw_gstatus_mpie = dcache_io_ptw_gstatus_mpie ; 
    wire dcache_tlb_io_ptw_gstatus_ube = dcache_io_ptw_gstatus_ube ; 
    wire dcache_tlb_io_ptw_gstatus_spie = dcache_io_ptw_gstatus_spie ; 
    wire dcache_tlb_io_ptw_gstatus_upie = dcache_io_ptw_gstatus_upie ; 
    wire dcache_tlb_io_ptw_gstatus_mie = dcache_io_ptw_gstatus_mie ; 
    wire dcache_tlb_io_ptw_gstatus_hie = dcache_io_ptw_gstatus_hie ; 
    wire dcache_tlb_io_ptw_gstatus_sie = dcache_io_ptw_gstatus_sie ; 
    wire dcache_tlb_io_ptw_gstatus_uie = dcache_io_ptw_gstatus_uie ; 
    wire dcache_tlb_io_ptw_pmp_0_cfg_l = dcache_io_ptw_pmp_0_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_0_cfg_res = dcache_io_ptw_pmp_0_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_0_cfg_a = dcache_io_ptw_pmp_0_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_0_cfg_x = dcache_io_ptw_pmp_0_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_0_cfg_w = dcache_io_ptw_pmp_0_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_0_cfg_r = dcache_io_ptw_pmp_0_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_0_addr = dcache_io_ptw_pmp_0_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_0_mask = dcache_io_ptw_pmp_0_mask ; 
    wire dcache_tlb_io_ptw_pmp_1_cfg_l = dcache_io_ptw_pmp_1_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_1_cfg_res = dcache_io_ptw_pmp_1_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_1_cfg_a = dcache_io_ptw_pmp_1_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_1_cfg_x = dcache_io_ptw_pmp_1_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_1_cfg_w = dcache_io_ptw_pmp_1_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_1_cfg_r = dcache_io_ptw_pmp_1_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_1_addr = dcache_io_ptw_pmp_1_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_1_mask = dcache_io_ptw_pmp_1_mask ; 
    wire dcache_tlb_io_ptw_pmp_2_cfg_l = dcache_io_ptw_pmp_2_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_2_cfg_res = dcache_io_ptw_pmp_2_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_2_cfg_a = dcache_io_ptw_pmp_2_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_2_cfg_x = dcache_io_ptw_pmp_2_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_2_cfg_w = dcache_io_ptw_pmp_2_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_2_cfg_r = dcache_io_ptw_pmp_2_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_2_addr = dcache_io_ptw_pmp_2_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_2_mask = dcache_io_ptw_pmp_2_mask ; 
    wire dcache_tlb_io_ptw_pmp_3_cfg_l = dcache_io_ptw_pmp_3_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_3_cfg_res = dcache_io_ptw_pmp_3_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_3_cfg_a = dcache_io_ptw_pmp_3_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_3_cfg_x = dcache_io_ptw_pmp_3_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_3_cfg_w = dcache_io_ptw_pmp_3_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_3_cfg_r = dcache_io_ptw_pmp_3_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_3_addr = dcache_io_ptw_pmp_3_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_3_mask = dcache_io_ptw_pmp_3_mask ; 
    wire dcache_tlb_io_ptw_pmp_4_cfg_l = dcache_io_ptw_pmp_4_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_4_cfg_res = dcache_io_ptw_pmp_4_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_4_cfg_a = dcache_io_ptw_pmp_4_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_4_cfg_x = dcache_io_ptw_pmp_4_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_4_cfg_w = dcache_io_ptw_pmp_4_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_4_cfg_r = dcache_io_ptw_pmp_4_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_4_addr = dcache_io_ptw_pmp_4_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_4_mask = dcache_io_ptw_pmp_4_mask ; 
    wire dcache_tlb_io_ptw_pmp_5_cfg_l = dcache_io_ptw_pmp_5_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_5_cfg_res = dcache_io_ptw_pmp_5_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_5_cfg_a = dcache_io_ptw_pmp_5_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_5_cfg_x = dcache_io_ptw_pmp_5_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_5_cfg_w = dcache_io_ptw_pmp_5_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_5_cfg_r = dcache_io_ptw_pmp_5_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_5_addr = dcache_io_ptw_pmp_5_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_5_mask = dcache_io_ptw_pmp_5_mask ; 
    wire dcache_tlb_io_ptw_pmp_6_cfg_l = dcache_io_ptw_pmp_6_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_6_cfg_res = dcache_io_ptw_pmp_6_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_6_cfg_a = dcache_io_ptw_pmp_6_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_6_cfg_x = dcache_io_ptw_pmp_6_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_6_cfg_w = dcache_io_ptw_pmp_6_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_6_cfg_r = dcache_io_ptw_pmp_6_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_6_addr = dcache_io_ptw_pmp_6_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_6_mask = dcache_io_ptw_pmp_6_mask ; 
    wire dcache_tlb_io_ptw_pmp_7_cfg_l = dcache_io_ptw_pmp_7_cfg_l ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_7_cfg_res = dcache_io_ptw_pmp_7_cfg_res ; 
    wire[1:0] dcache_tlb_io_ptw_pmp_7_cfg_a = dcache_io_ptw_pmp_7_cfg_a ; 
    wire dcache_tlb_io_ptw_pmp_7_cfg_x = dcache_io_ptw_pmp_7_cfg_x ; 
    wire dcache_tlb_io_ptw_pmp_7_cfg_w = dcache_io_ptw_pmp_7_cfg_w ; 
    wire dcache_tlb_io_ptw_pmp_7_cfg_r = dcache_io_ptw_pmp_7_cfg_r ; 
    wire[29:0] dcache_tlb_io_ptw_pmp_7_addr = dcache_io_ptw_pmp_7_addr ; 
    wire[31:0] dcache_tlb_io_ptw_pmp_7_mask = dcache_io_ptw_pmp_7_mask ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_0_ren = dcache_io_ptw_customCSRs_csrs_0_ren ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_0_wen = dcache_io_ptw_customCSRs_csrs_0_wen ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_0_wdata = dcache_io_ptw_customCSRs_csrs_0_wdata ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_0_value = dcache_io_ptw_customCSRs_csrs_0_value ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_1_ren = dcache_io_ptw_customCSRs_csrs_1_ren ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_1_wen = dcache_io_ptw_customCSRs_csrs_1_wen ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_1_wdata = dcache_io_ptw_customCSRs_csrs_1_wdata ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_1_value = dcache_io_ptw_customCSRs_csrs_1_value ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_2_ren = dcache_io_ptw_customCSRs_csrs_2_ren ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_2_wen = dcache_io_ptw_customCSRs_csrs_2_wen ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_2_wdata = dcache_io_ptw_customCSRs_csrs_2_wdata ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_2_value = dcache_io_ptw_customCSRs_csrs_2_value ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_3_ren = dcache_io_ptw_customCSRs_csrs_3_ren ; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_3_wen = dcache_io_ptw_customCSRs_csrs_3_wen ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_3_wdata = dcache_io_ptw_customCSRs_csrs_3_wdata ; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_3_value = dcache_io_ptw_customCSRs_csrs_3_value ; 
    wire dcache_pma_checker_clock = dcache_clock ; 
    wire dcache_pma_checker_reset = dcache_reset ; 
    wire dcache_metaArb_clock = dcache_clock ; 
    wire dcache_metaArb_reset = dcache_reset ; 
    wire dcache_metaArb_io_in_7_valid = dcache_io_cpu_req_valid ; 
    wire[33:0] dcache_metaArb_io_in_7_bits_addr = dcache_io_cpu_req_bits_addr ; 
    wire dcache_tag_array_MPORT_clk = dcache_clock ; 
    wire dcache_tag_array_s1_meta_clk = dcache_clock ; 
    wire dcache_dataArb_clock = dcache_clock ; 
    wire dcache_dataArb_reset = dcache_reset ; 
    wire[5:0] dcache_s0_req_tag = dcache_io_cpu_req_bits_tag ; 
    wire[4:0] dcache_s0_req_cmd = dcache_io_cpu_req_bits_cmd ; 
    wire[1:0] dcache_s0_req_size = dcache_io_cpu_req_bits_size ; 
    wire dcache_s0_req_signed = dcache_io_cpu_req_bits_signed ; 
    wire[1:0] dcache_s0_req_dprv = dcache_io_cpu_req_bits_dprv ; 
    wire dcache_s0_req_dv = dcache_io_cpu_req_bits_dv ; 
    wire dcache_s0_req_no_alloc = dcache_io_cpu_req_bits_no_alloc ; 
    wire dcache_s0_req_no_xcpt = dcache_io_cpu_req_bits_no_xcpt ; 
    wire[63:0] dcache_s0_req_data = dcache_io_cpu_req_bits_data ; 
    wire[7:0] dcache_s0_req_mask = dcache_io_cpu_req_bits_mask ; 
    wire[2:0] dcache_atomics_a_param =3'h3; 
    wire[2:0] dcache_atomics_a_8_param =3'h3; 
    wire[2:0] dcache_atomics_a_2_param =3'h1; 
    wire[2:0] dcache_atomics_a_6_param =3'h1; 
    wire[2:0] dcache_atomics_a_3_param =3'h2; 
    wire[2:0] dcache_atomics_a_7_param =3'h2; 
    wire[9:0] dcache_pma_checker_io_ptw_resp_bits_pte_reserved_for_future =10'h0; 
    wire[15:0] dcache_pma_checker_io_ptw_ptbr_asid =16'h0; 
    wire[15:0] dcache_pma_checker_io_ptw_hgatp_asid =16'h0; 
    wire[15:0] dcache_pma_checker_io_ptw_vsatp_asid =16'h0; 
    wire[43:0] dcache_pma_checker_io_ptw_resp_bits_pte_ppn =44'h0; 
    wire[43:0] dcache_pma_checker_io_ptw_ptbr_ppn =44'h0; 
    wire[43:0] dcache_pma_checker_io_ptw_hgatp_ppn =44'h0; 
    wire[43:0] dcache_pma_checker_io_ptw_vsatp_ppn =44'h0; 
    wire[8:0] dcache_pma_checker_io_ptw_hstatus_zero5 =9'h0; 
    wire[22:0] dcache_pma_checker_io_ptw_status_zero2 =23'h0; 
    wire[22:0] dcache_pma_checker_io_ptw_gstatus_zero2 =23'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_status_isa =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_gstatus_isa =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_0_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_1_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_2_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_3_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_4_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_5_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_6_mask =32'h0; 
    wire[31:0] dcache_pma_checker_io_ptw_pmp_7_mask =32'h0; 
    wire[31:0] dcache__atomics_WIRE_address =32'h0; 
    wire[31:0] dcache__io_cpu_s2_xcpt_WIRE_paddr =32'h0; 
    wire[7:0] dcache_dataArb_io_in_1_bits_eccMask =8'hFF; 
    wire[7:0] dcache_dataArb_io_in_2_bits_eccMask =8'hFF; 
    wire[7:0] dcache_dataArb_io_in_3_bits_eccMask =8'hFF; 
    wire[2:0] dcache_nackResponseMessage_param =3'h5; 
    wire[2:0] dcache_dirtyReleaseMessage_opcode =3'h5; 
    wire[2:0] dcache_get_opcode =3'h4; 
    wire[2:0] dcache_atomics_a_4_param =3'h4; 
    wire[2:0] dcache_nackResponseMessage_opcode =3'h4; 
    wire[2:0] dcache_cleanReleaseMessage_opcode =3'h4; 
    wire[2:0] dcache_nodeOut_c_bits_c_1_opcode =3'h7; 
    wire[2:0] dcache_tl_out_a_bits_a_opcode =3'h6; 
    wire[2:0] dcache_nodeOut_c_bits_c_opcode =3'h6; 
    wire[33:0] dcache__io_cpu_s2_xcpt_WIRE_gpa =34'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_hstatus_zero6 =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_0_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_1_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_2_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_3_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_4_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_5_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_6_addr =30'h0; 
    wire[29:0] dcache_pma_checker_io_ptw_pmp_7_addr =30'h0; 
    wire[3:0] dcache_pma_checker_io_ptw_ptbr_mode =4'h0; 
    wire[3:0] dcache_pma_checker_io_ptw_hgatp_mode =4'h0; 
    wire[3:0] dcache_pma_checker_io_ptw_vsatp_mode =4'h0; 
    wire[3:0] dcache__atomics_WIRE_size =4'h0; 
    wire[3:0] dcache_probe_bits_res_size =4'h0; 
    wire[4:0] dcache_pma_checker_io_ptw_hstatus_zero1 =5'h0; 
    wire[1:0] dcache_tl_out_a_bits_a_mask_sizeOH_shiftAmount =2'h2; 
    wire[2:0] dcache__atomics_WIRE_opcode =3'h0; 
    wire[2:0] dcache__atomics_WIRE_param =3'h0; 
    wire[2:0] dcache_atomics_a_1_param =3'h0; 
    wire[2:0] dcache_atomics_a_5_param =3'h0; 
    wire[2:0] dcache_probe_bits_res_opcode =3'h0; 
    wire[32:0] dcache_pma_checker_io_sfence_bits_addr =33'h0; 
    wire[32:0] dcache_pma_checker_io_ptw_resp_bits_gpa_bits =33'h0; 
    wire[7:0] dcache_pma_checker_io_ptw_status_zero1 =8'h0; 
    wire[7:0] dcache_pma_checker_io_ptw_gstatus_zero1 =8'h0; 
    wire[7:0] dcache__atomics_WIRE_mask =8'h0; 
    wire[7:0] dcache_probe_bits_res_mask =8'h0; 
    wire[5:0] dcache_tlb_stage1_bypass =6'h0; 
    wire[5:0] dcache_pma_checker_io_ptw_hstatus_vgein =6'h0; 
    wire[5:0] dcache_pma_checker_stage1_bypass =6'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_resp_bits_pte_reserved_for_software =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_resp_bits_level =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_dprv =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_prv =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_sxl =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_uxl =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_xs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_fs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_mpp =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_status_vs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_hstatus_vsxl =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_hstatus_zero3 =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_hstatus_zero2 =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_dprv =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_prv =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_sxl =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_uxl =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_xs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_fs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_mpp =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_gstatus_vs =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_0_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_0_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_1_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_1_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_2_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_2_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_3_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_3_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_4_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_4_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_5_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_5_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_6_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_6_cfg_a =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_7_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_io_ptw_pmp_7_cfg_a =2'h0; 
    wire[1:0] dcache_s1_meta_hit_state_meta_state =2'h0; 
    wire[1:0] dcache_metaArb_io_in_1_bits_data_new_meta_coh_meta_state =2'h0; 
    wire[1:0] dcache_probe_bits_res_param =2'h0; 
    wire[1:0] dcache_metaArb_io_in_0_bits_data_meta_state =2'h0; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_0_sdata =64'h0; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_1_sdata =64'h0; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_2_sdata =64'h0; 
    wire[63:0] dcache_tlb_io_ptw_customCSRs_csrs_3_sdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_0_wdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_0_value =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_0_sdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_1_wdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_1_value =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_1_sdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_2_wdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_2_value =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_2_sdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_3_wdata =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_3_value =64'h0; 
    wire[63:0] dcache_pma_checker_io_ptw_customCSRs_csrs_3_sdata =64'h0; 
    wire[63:0] dcache__atomics_WIRE_data =64'h0; 
    wire[63:0] dcache_probe_bits_res_data =64'h0; 
    wire dcache_nodeOut_c_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_tlb_io_resp_ma_inst =1'h0; 
    wire dcache_tlb_io_resp_prefetchable =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_0_stall =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_0_set =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_1_stall =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_1_set =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_2_stall =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_2_set =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_3_stall =1'h0; 
    wire dcache_tlb_io_ptw_customCSRs_csrs_3_set =1'h0; 
    wire dcache_tlb_priv_v =1'h0; 
    wire dcache_tlb_stage1_en =1'h0; 
    wire dcache_tlb_vstage1_en =1'h0; 
    wire dcache_tlb_stage2_en =1'h0; 
    wire dcache_tlb_do_refill =1'h0; 
    wire dcache_tlb_cmd_readx =1'h0; 
    wire dcache_pma_checker_io_req_valid =1'h0; 
    wire dcache_pma_checker_io_resp_ma_inst =1'h0; 
    wire dcache_pma_checker_io_resp_prefetchable =1'h0; 
    wire dcache_pma_checker_io_sfence_valid =1'h0; 
    wire dcache_pma_checker_io_sfence_bits_rs1 =1'h0; 
    wire dcache_pma_checker_io_sfence_bits_rs2 =1'h0; 
    wire dcache_pma_checker_io_sfence_bits_asid =1'h0; 
    wire dcache_pma_checker_io_sfence_bits_hv =1'h0; 
    wire dcache_pma_checker_io_sfence_bits_hg =1'h0; 
    wire dcache_pma_checker_io_ptw_req_ready =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_valid =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_ae_ptw =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_ae_final =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pf =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_gf =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_hr =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_hw =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_hx =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_d =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_a =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_g =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_u =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_x =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_w =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_r =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_pte_v =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_fragmented_superpage =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_homogeneous =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_gpa_valid =1'h0; 
    wire dcache_pma_checker_io_ptw_resp_bits_gpa_is_pte =1'h0; 
    wire dcache_pma_checker_io_ptw_status_debug =1'h0; 
    wire dcache_pma_checker_io_ptw_status_cease =1'h0; 
    wire dcache_pma_checker_io_ptw_status_wfi =1'h0; 
    wire dcache_pma_checker_io_ptw_status_dv =1'h0; 
    wire dcache_pma_checker_io_ptw_status_v =1'h0; 
    wire dcache_pma_checker_io_ptw_status_sd =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mpv =1'h0; 
    wire dcache_pma_checker_io_ptw_status_gva =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mbe =1'h0; 
    wire dcache_pma_checker_io_ptw_status_sbe =1'h0; 
    wire dcache_pma_checker_io_ptw_status_sd_rv32 =1'h0; 
    wire dcache_pma_checker_io_ptw_status_tsr =1'h0; 
    wire dcache_pma_checker_io_ptw_status_tw =1'h0; 
    wire dcache_pma_checker_io_ptw_status_tvm =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mxr =1'h0; 
    wire dcache_pma_checker_io_ptw_status_sum =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mprv =1'h0; 
    wire dcache_pma_checker_io_ptw_status_spp =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mpie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_ube =1'h0; 
    wire dcache_pma_checker_io_ptw_status_spie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_upie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_mie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_hie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_sie =1'h0; 
    wire dcache_pma_checker_io_ptw_status_uie =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_vtsr =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_vtw =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_vtvm =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_hu =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_spvp =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_spv =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_gva =1'h0; 
    wire dcache_pma_checker_io_ptw_hstatus_vsbe =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_debug =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_cease =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_wfi =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_dv =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_v =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_sd =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mpv =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_gva =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mbe =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_sbe =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_sd_rv32 =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_tsr =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_tw =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_tvm =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mxr =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_sum =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mprv =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_spp =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mpie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_ube =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_spie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_upie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_mie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_hie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_sie =1'h0; 
    wire dcache_pma_checker_io_ptw_gstatus_uie =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_0_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_0_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_0_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_0_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_1_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_1_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_1_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_1_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_2_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_2_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_2_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_2_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_3_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_3_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_3_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_3_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_4_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_4_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_4_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_4_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_5_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_5_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_5_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_5_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_6_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_6_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_6_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_6_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_7_cfg_l =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_7_cfg_x =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_7_cfg_w =1'h0; 
    wire dcache_pma_checker_io_ptw_pmp_7_cfg_r =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_0_ren =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_0_wen =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_0_stall =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_0_set =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_1_ren =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_1_wen =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_1_stall =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_1_set =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_2_ren =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_2_wen =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_2_stall =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_2_set =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_3_ren =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_3_wen =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_3_stall =1'h0; 
    wire dcache_pma_checker_io_ptw_customCSRs_csrs_3_set =1'h0; 
    wire dcache_pma_checker_io_kill =1'h0; 
    wire dcache_pma_checker_priv_v =1'h0; 
    wire dcache_pma_checker_stage1_en =1'h0; 
    wire dcache_pma_checker_vstage1_en =1'h0; 
    wire dcache_pma_checker_stage2_en =1'h0; 
    wire dcache_pma_checker_do_refill =1'h0; 
    wire dcache_pma_checker_cmd_readx =1'h0; 
    wire dcache_metaArb_io_in_5_bits_write =1'h0; 
    wire dcache_metaArb_io_in_6_bits_write =1'h0; 
    wire dcache_metaArb_io_in_7_bits_write =1'h0; 
    wire dcache_dataArb_io_in_2_bits_write =1'h0; 
    wire dcache_dataArb_io_in_3_bits_write =1'h0; 
    wire dcache_tl_out_a_bits_user_amba_prot_fetch =1'h0; 
    wire dcache_s1_waw_hazard =1'h0; 
    wire dcache__uncachedInFlight_WIRE_0 =1'h0; 
    wire dcache_s1_victim_way =1'h0; 
    wire dcache_s2_store_merge =1'h0; 
    wire dcache_s2_data_error =1'h0; 
    wire dcache_s2_data_error_uncorrectable =1'h0; 
    wire dcache_s2_correct =1'h0; 
    wire dcache_dataArb_io_in_0_valid_s2_kill =1'h0; 
    wire dcache_get_user_amba_prot_bufferable =1'h0; 
    wire dcache_get_user_amba_prot_modifiable =1'h0; 
    wire dcache_get_user_amba_prot_readalloc =1'h0; 
    wire dcache_get_user_amba_prot_writealloc =1'h0; 
    wire dcache_get_user_amba_prot_privileged =1'h0; 
    wire dcache_get_user_amba_prot_secure =1'h0; 
    wire dcache_get_user_amba_prot_fetch =1'h0; 
    wire dcache_get_corrupt =1'h0; 
    wire dcache_put_user_amba_prot_bufferable =1'h0; 
    wire dcache_put_user_amba_prot_modifiable =1'h0; 
    wire dcache_put_user_amba_prot_readalloc =1'h0; 
    wire dcache_put_user_amba_prot_writealloc =1'h0; 
    wire dcache_put_user_amba_prot_privileged =1'h0; 
    wire dcache_put_user_amba_prot_secure =1'h0; 
    wire dcache_put_user_amba_prot_fetch =1'h0; 
    wire dcache_put_corrupt =1'h0; 
    wire dcache_putpartial_user_amba_prot_bufferable =1'h0; 
    wire dcache_putpartial_user_amba_prot_modifiable =1'h0; 
    wire dcache_putpartial_user_amba_prot_readalloc =1'h0; 
    wire dcache_putpartial_user_amba_prot_writealloc =1'h0; 
    wire dcache_putpartial_user_amba_prot_privileged =1'h0; 
    wire dcache_putpartial_user_amba_prot_secure =1'h0; 
    wire dcache_putpartial_user_amba_prot_fetch =1'h0; 
    wire dcache_putpartial_corrupt =1'h0; 
    wire dcache__atomics_WIRE_source =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_bufferable =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_modifiable =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_readalloc =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_writealloc =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_privileged =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_secure =1'h0; 
    wire dcache__atomics_WIRE_user_amba_prot_fetch =1'h0; 
    wire dcache__atomics_WIRE_corrupt =1'h0; 
    wire dcache_atomics_a_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_corrupt =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_1_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_1_corrupt =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_2_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_2_corrupt =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_3_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_3_corrupt =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_4_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_4_corrupt =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_5_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_5_corrupt =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_6_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_6_corrupt =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_7_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_7_corrupt =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_bufferable =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_modifiable =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_readalloc =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_writealloc =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_privileged =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_secure =1'h0; 
    wire dcache_atomics_a_8_user_amba_prot_fetch =1'h0; 
    wire dcache_atomics_a_8_corrupt =1'h0; 
    wire dcache_tl_out_a_bits_a_source =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_bufferable =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_modifiable =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_readalloc =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_writealloc =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_privileged =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_secure =1'h0; 
    wire dcache_tl_out_a_bits_a_user_amba_prot_fetch =1'h0; 
    wire dcache_tl_out_a_bits_a_corrupt =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_nackResponseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_nackResponseMessage_corrupt =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_cleanReleaseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_cleanReleaseMessage_corrupt =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_bufferable =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_modifiable =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_readalloc =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_writealloc =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_privileged =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_secure =1'h0; 
    wire dcache_dirtyReleaseMessage_user_amba_prot_fetch =1'h0; 
    wire dcache_dirtyReleaseMessage_corrupt =1'h0; 
    wire dcache_probe_bits_res_source =1'h0; 
    wire dcache_probe_bits_res_corrupt =1'h0; 
    wire dcache_nodeOut_c_bits_legal =1'h0; 
    wire dcache_nodeOut_c_bits_c_source =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_bufferable =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_modifiable =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_readalloc =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_writealloc =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_privileged =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_secure =1'h0; 
    wire dcache_nodeOut_c_bits_c_user_amba_prot_fetch =1'h0; 
    wire dcache_nodeOut_c_bits_c_corrupt =1'h0; 
    wire dcache_nodeOut_c_bits_legal_1 =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_source =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_bufferable =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_modifiable =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_readalloc =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_writealloc =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_privileged =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_secure =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_user_amba_prot_fetch =1'h0; 
    wire dcache_nodeOut_c_bits_c_1_corrupt =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_miss =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_gpa_is_pte =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_pf_ld =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_pf_st =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_pf_inst =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_gf_ld =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_gf_st =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_gf_inst =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ae_ld =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ae_st =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ae_inst =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ma_ld =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ma_st =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_ma_inst =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_cacheable =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_must_alloc =1'h0; 
    wire dcache__io_cpu_s2_xcpt_WIRE_prefetchable =1'h0; 
    wire dcache_io_cpu_resp_bits_data_doZero =1'h0; 
    wire dcache_io_cpu_resp_bits_data_doZero_1 =1'h0; 
    wire dcache_io_cpu_resp_bits_data_word_bypass_doZero =1'h0; 
    wire dcache_nodeOut_c_bits_user_amba_prot_bufferable =1'h1; 
    wire dcache_nodeOut_c_bits_user_amba_prot_modifiable =1'h1; 
    wire dcache_nodeOut_c_bits_user_amba_prot_readalloc =1'h1; 
    wire dcache_nodeOut_c_bits_user_amba_prot_writealloc =1'h1; 
    wire dcache_nodeOut_c_bits_user_amba_prot_privileged =1'h1; 
    wire dcache_nodeOut_c_bits_user_amba_prot_secure =1'h1; 
    wire dcache_pma_checker_io_req_bits_passthrough =1'h1; 
    wire dcache_metaArb_io_in_0_bits_write =1'h1; 
    wire dcache_metaArb_io_in_0_bits_way_en =1'h1; 
    wire dcache_metaArb_io_in_1_bits_write =1'h1; 
    wire dcache_metaArb_io_in_3_bits_write =1'h1; 
    wire dcache_metaArb_io_in_4_bits_write =1'h1; 
    wire dcache_tag_array_MPORT_mask_0 =1'h1; 
    wire dcache_dataArb_io_in_1_bits_wordMask =1'h1; 
    wire dcache_dataArb_io_in_2_bits_wordMask =1'h1; 
    wire dcache_dataArb_io_in_2_bits_way_en =1'h1; 
    wire dcache_dataArb_io_in_3_bits_wordMask =1'h1; 
    wire dcache_dataArb_io_in_3_bits_way_en =1'h1; 
    wire dcache_dataArb_io_out_ready =1'h1; 
    wire dcache_tl_out_a_bits_user_amba_prot_secure =1'h1; 
    wire dcache_tl_out_a_bits_a_mask_acc =1'h1; 
    wire dcache_tl_out_a_bits_a_mask_acc_1 =1'h1; 
    wire dcache_tlb_io_ptw_req_valid ; 
    wire dcache_nodeOut_a_deq_ready = dcache_nodeOut_a_ready ; 
    wire dcache_nodeOut_a_deq_valid ; 
    wire[2:0] dcache_nodeOut_a_deq_bits_opcode ; 
    wire[2:0] dcache_nodeOut_a_deq_bits_param ; 
    wire[3:0] dcache_nodeOut_a_deq_bits_size ; 
    wire dcache_nodeOut_a_deq_bits_source ; 
    wire[31:0] dcache_nodeOut_a_deq_bits_address ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_privileged ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_secure ; 
    wire dcache_nodeOut_a_deq_bits_user_amba_prot_fetch ; 
    wire[7:0] dcache_nodeOut_a_deq_bits_mask ; 
    wire[63:0] dcache_nodeOut_a_deq_bits_data ; 
    wire dcache_nodeOut_a_deq_bits_corrupt ; 
    wire[63:0] dcache_s2_data_corrected ; 
    wire dcache_uncachedRespIdxOH_shiftAmount = dcache_nodeOut_d_bits_source ; 
    wire[1:0] dcache_nodeOut_e_bits_e_sink = dcache_nodeOut_d_bits_sink ; 
    wire[63:0] dcache_s1_uncached_data_word = dcache_nodeOut_d_bits_data ; 
    reg dcache_clock_en_reg ; 
    wire dcache__tlb_port_req_ready_output = dcache_clock_en_reg ; 
    wire dcache_metaArb_io_out_ready = dcache_clock_en_reg ; 
    wire dcache__io_ptw_req_valid_output = dcache_tlb_io_ptw_req_valid ; 
    wire dcache_tlb_newEntry_ae_ptw = dcache_tlb_io_ptw_resp_bits_ae_ptw ; 
    wire dcache_tlb_newEntry_ae_final = dcache_tlb_io_ptw_resp_bits_ae_final ; 
    wire dcache_tlb_newEntry_pf = dcache_tlb_io_ptw_resp_bits_pf ; 
    wire dcache_tlb_newEntry_gf = dcache_tlb_io_ptw_resp_bits_gf ; 
    wire dcache_tlb_newEntry_hr = dcache_tlb_io_ptw_resp_bits_hr ; 
    wire dcache_tlb_newEntry_hw = dcache_tlb_io_ptw_resp_bits_hw ; 
    wire dcache_tlb_newEntry_hx = dcache_tlb_io_ptw_resp_bits_hx ; 
    wire dcache_tlb_newEntry_u = dcache_tlb_io_ptw_resp_bits_pte_u ; 
    wire dcache_tlb_newEntry_fragmented_superpage = dcache_tlb_io_ptw_resp_bits_fragmented_superpage ; 
    wire[33:0] dcache_tlb_io_req_bits_vaddr ; 
    wire[20:0] dcache_tlb_vpn = dcache_tlb_io_req_bits_vaddr [32:12]; reg[1:0] dcache_tlb_sectored_entries_0_0_level ; reg[20:0] dcache_tlb_sectored_entries_0_0_tag_vpn ; 
    reg dcache_tlb_sectored_entries_0_0_tag_v ; reg[41:0] dcache_tlb_sectored_entries_0_0_data_0 ; reg[41:0] dcache_tlb_sectored_entries_0_0_data_1 ; reg[41:0] dcache_tlb_sectored_entries_0_0_data_2 ; reg[41:0] dcache_tlb_sectored_entries_0_0_data_3 ; 
    reg dcache_tlb_sectored_entries_0_0_valid_0 ; 
    reg dcache_tlb_sectored_entries_0_0_valid_1 ; 
    reg dcache_tlb_sectored_entries_0_0_valid_2 ; 
    reg dcache_tlb_sectored_entries_0_0_valid_3 ; reg[1:0] dcache_tlb_superpage_entries_0_level ; reg[20:0] dcache_tlb_superpage_entries_0_tag_vpn ; 
    reg dcache_tlb_superpage_entries_0_tag_v ; reg[41:0] dcache_tlb_superpage_entries_0_data_0 ; 
    wire[41:0] dcache_tlb__entries_WIRE_3 = dcache_tlb_superpage_entries_0_data_0 ; 
    reg dcache_tlb_superpage_entries_0_valid_0 ; reg[1:0] dcache_tlb_superpage_entries_1_level ; reg[20:0] dcache_tlb_superpage_entries_1_tag_vpn ; 
    reg dcache_tlb_superpage_entries_1_tag_v ; reg[41:0] dcache_tlb_superpage_entries_1_data_0 ; 
    wire[41:0] dcache_tlb__entries_WIRE_5 = dcache_tlb_superpage_entries_1_data_0 ; 
    reg dcache_tlb_superpage_entries_1_valid_0 ; reg[1:0] dcache_tlb_superpage_entries_2_level ; reg[20:0] dcache_tlb_superpage_entries_2_tag_vpn ; 
    reg dcache_tlb_superpage_entries_2_tag_v ; reg[41:0] dcache_tlb_superpage_entries_2_data_0 ; 
    wire[41:0] dcache_tlb__entries_WIRE_7 = dcache_tlb_superpage_entries_2_data_0 ; 
    reg dcache_tlb_superpage_entries_2_valid_0 ; reg[1:0] dcache_tlb_superpage_entries_3_level ; reg[20:0] dcache_tlb_superpage_entries_3_tag_vpn ; 
    reg dcache_tlb_superpage_entries_3_tag_v ; reg[41:0] dcache_tlb_superpage_entries_3_data_0 ; 
    wire[41:0] dcache_tlb__entries_WIRE_9 = dcache_tlb_superpage_entries_3_data_0 ; 
    reg dcache_tlb_superpage_entries_3_valid_0 ; reg[1:0] dcache_tlb_special_entry_level ; reg[20:0] dcache_tlb_special_entry_tag_vpn ; 
    reg dcache_tlb_special_entry_tag_v ; reg[41:0] dcache_tlb_special_entry_data_0 ; 
    wire[41:0] dcache_tlb__mpu_ppn_WIRE_1 = dcache_tlb_special_entry_data_0 ; 
    wire[41:0] dcache_tlb__entries_WIRE_11 = dcache_tlb_special_entry_data_0 ; 
    reg dcache_tlb_special_entry_valid_0 ; reg[1:0] dcache_tlb_state ; reg[20:0] dcache_tlb_r_refill_tag ; 
    wire[20:0] dcache_tlb_io_ptw_req_bits_bits_addr = dcache_tlb_r_refill_tag ; reg[1:0] dcache_tlb_r_superpage_repl_addr ; 
    wire[1:0] dcache_tlb_waddr = dcache_tlb_r_superpage_repl_addr ; 
    reg dcache_tlb_r_sectored_hit_valid ; 
    reg dcache_tlb_r_superpage_hit_valid ; reg[1:0] dcache_tlb_r_superpage_hit_bits ; 
    reg dcache_tlb_r_vstage1_en ; 
    wire dcache_tlb_io_ptw_req_bits_bits_vstage1 = dcache_tlb_r_vstage1_en ; 
    reg dcache_tlb_r_stage2_en ; 
    wire dcache_tlb_io_ptw_req_bits_bits_stage2 = dcache_tlb_r_stage2_en ; 
    reg dcache_tlb_r_need_gpa ; 
    wire dcache_tlb_io_ptw_req_bits_bits_need_gpa = dcache_tlb_r_need_gpa ; 
    reg dcache_tlb_r_gpa_valid ; reg[32:0] dcache_tlb_r_gpa ; reg[20:0] dcache_tlb_r_gpa_vpn ; 
    reg dcache_tlb_r_gpa_is_pte ; 
    wire[1:0] dcache_tlb_io_req_bits_prv ; 
    wire dcache_tlb_priv_s = dcache_tlb_io_req_bits_prv [0]; 
    wire dcache_tlb_priv_uses_vm = dcache_tlb_io_req_bits_prv <=2'h1; 
    wire[3:0] dcache_tlb_satp_mode = dcache_tlb_priv_v  ?  dcache_tlb_io_ptw_vsatp_mode : dcache_tlb_io_ptw_ptbr_mode ; 
    wire[15:0] dcache_tlb_satp_asid = dcache_tlb_priv_v  ?  dcache_tlb_io_ptw_vsatp_asid : dcache_tlb_io_ptw_ptbr_asid ; 
    wire[43:0] dcache_tlb_satp_ppn = dcache_tlb_priv_v  ?  dcache_tlb_io_ptw_vsatp_ppn : dcache_tlb_io_ptw_ptbr_ppn ; 
    wire dcache_tlb_io_req_bits_passthrough ; 
    wire dcache_tlb_vm_enabled =( dcache_tlb_stage1_en | dcache_tlb_stage2_en )& dcache_tlb_priv_uses_vm & dcache_tlb_io_req_bits_passthrough ==1'h0; 
    reg dcache_tlb_v_entries_use_stage1 ; 
    wire dcache_tlb_vsatp_mode_mismatch = dcache_tlb_priv_v & dcache_tlb_vstage1_en != dcache_tlb_v_entries_use_stage1 & dcache_tlb_io_req_bits_passthrough ==1'h0; 
    wire[19:0] dcache_tlb_refill_ppn = dcache_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire dcache_tlb_io_sfence_valid ; 
    wire dcache_tlb_invalidate_refill = dcache_tlb_state ==2'h1|(& dcache_tlb_state )| dcache_tlb_io_sfence_valid ; 
    wire dcache_tlb__mpu_ppn_WIRE_fragmented_superpage = dcache_tlb__mpu_ppn_WIRE_1 [0]; 
    wire dcache_tlb__mpu_ppn_WIRE_c = dcache_tlb__mpu_ppn_WIRE_1 [1]; 
    wire dcache_tlb__mpu_ppn_WIRE_eff = dcache_tlb__mpu_ppn_WIRE_1 [2]; 
    wire dcache_tlb__mpu_ppn_WIRE_paa = dcache_tlb__mpu_ppn_WIRE_1 [3]; 
    wire dcache_tlb__mpu_ppn_WIRE_pal = dcache_tlb__mpu_ppn_WIRE_1 [4]; 
    wire dcache_tlb__mpu_ppn_WIRE_ppp = dcache_tlb__mpu_ppn_WIRE_1 [5]; 
    wire dcache_tlb__mpu_ppn_WIRE_pr = dcache_tlb__mpu_ppn_WIRE_1 [6]; 
    wire dcache_tlb__mpu_ppn_WIRE_px = dcache_tlb__mpu_ppn_WIRE_1 [7]; 
    wire dcache_tlb__mpu_ppn_WIRE_pw = dcache_tlb__mpu_ppn_WIRE_1 [8]; 
    wire dcache_tlb__mpu_ppn_WIRE_hr = dcache_tlb__mpu_ppn_WIRE_1 [9]; 
    wire dcache_tlb__mpu_ppn_WIRE_hx = dcache_tlb__mpu_ppn_WIRE_1 [10]; 
    wire dcache_tlb__mpu_ppn_WIRE_hw = dcache_tlb__mpu_ppn_WIRE_1 [11]; 
    wire dcache_tlb__mpu_ppn_WIRE_sr = dcache_tlb__mpu_ppn_WIRE_1 [12]; 
    wire dcache_tlb__mpu_ppn_WIRE_sx = dcache_tlb__mpu_ppn_WIRE_1 [13]; 
    wire dcache_tlb__mpu_ppn_WIRE_sw = dcache_tlb__mpu_ppn_WIRE_1 [14]; 
    wire dcache_tlb__mpu_ppn_WIRE_gf = dcache_tlb__mpu_ppn_WIRE_1 [15]; 
    wire dcache_tlb__mpu_ppn_WIRE_pf = dcache_tlb__mpu_ppn_WIRE_1 [16]; 
    wire dcache_tlb__mpu_ppn_WIRE_ae_stage2 = dcache_tlb__mpu_ppn_WIRE_1 [17]; 
    wire dcache_tlb__mpu_ppn_WIRE_ae_final = dcache_tlb__mpu_ppn_WIRE_1 [18]; 
    wire dcache_tlb__mpu_ppn_WIRE_ae_ptw = dcache_tlb__mpu_ppn_WIRE_1 [19]; 
    wire dcache_tlb__mpu_ppn_WIRE_g = dcache_tlb__mpu_ppn_WIRE_1 [20]; 
    wire dcache_tlb__mpu_ppn_WIRE_u = dcache_tlb__mpu_ppn_WIRE_1 [21]; 
    wire[19:0] dcache_tlb__mpu_ppn_WIRE_ppn = dcache_tlb__mpu_ppn_WIRE_1 [41:22];  
    wire dcache_tlb_mpu_ppn_barrier_clock;
    wire dcache_tlb_mpu_ppn_barrier_reset;
    wire[19:0] dcache_tlb_mpu_ppn_barrier_io_x_ppn;
    wire dcache_tlb_mpu_ppn_barrier_io_x_u;
    wire dcache_tlb_mpu_ppn_barrier_io_x_g;
    wire dcache_tlb_mpu_ppn_barrier_io_x_ae_ptw;
    wire dcache_tlb_mpu_ppn_barrier_io_x_ae_final;
    wire dcache_tlb_mpu_ppn_barrier_io_x_ae_stage2;
    wire dcache_tlb_mpu_ppn_barrier_io_x_pf;
    wire dcache_tlb_mpu_ppn_barrier_io_x_gf;
    wire dcache_tlb_mpu_ppn_barrier_io_x_sw;
    wire dcache_tlb_mpu_ppn_barrier_io_x_sx;
    wire dcache_tlb_mpu_ppn_barrier_io_x_sr;
    wire dcache_tlb_mpu_ppn_barrier_io_x_hw;
    wire dcache_tlb_mpu_ppn_barrier_io_x_hx;
    wire dcache_tlb_mpu_ppn_barrier_io_x_hr;
    wire dcache_tlb_mpu_ppn_barrier_io_x_pw;
    wire dcache_tlb_mpu_ppn_barrier_io_x_px;
    wire dcache_tlb_mpu_ppn_barrier_io_x_pr;
    wire dcache_tlb_mpu_ppn_barrier_io_x_ppp;
    wire dcache_tlb_mpu_ppn_barrier_io_x_pal;
    wire dcache_tlb_mpu_ppn_barrier_io_x_paa;
    wire dcache_tlb_mpu_ppn_barrier_io_x_eff;
    wire dcache_tlb_mpu_ppn_barrier_io_x_c;
    wire dcache_tlb_mpu_ppn_barrier_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_mpu_ppn_barrier_io_y_ppn;
    wire dcache_tlb_mpu_ppn_barrier_io_y_u;
    wire dcache_tlb_mpu_ppn_barrier_io_y_g;
    wire dcache_tlb_mpu_ppn_barrier_io_y_ae_ptw;
    wire dcache_tlb_mpu_ppn_barrier_io_y_ae_final;
    wire dcache_tlb_mpu_ppn_barrier_io_y_ae_stage2;
    wire dcache_tlb_mpu_ppn_barrier_io_y_pf;
    wire dcache_tlb_mpu_ppn_barrier_io_y_gf;
    wire dcache_tlb_mpu_ppn_barrier_io_y_sw;
    wire dcache_tlb_mpu_ppn_barrier_io_y_sx;
    wire dcache_tlb_mpu_ppn_barrier_io_y_sr;
    wire dcache_tlb_mpu_ppn_barrier_io_y_hw;
    wire dcache_tlb_mpu_ppn_barrier_io_y_hx;
    wire dcache_tlb_mpu_ppn_barrier_io_y_hr;
    wire dcache_tlb_mpu_ppn_barrier_io_y_pw;
    wire dcache_tlb_mpu_ppn_barrier_io_y_px;
    wire dcache_tlb_mpu_ppn_barrier_io_y_pr;
    wire dcache_tlb_mpu_ppn_barrier_io_y_ppp;
    wire dcache_tlb_mpu_ppn_barrier_io_y_pal;
    wire dcache_tlb_mpu_ppn_barrier_io_y_paa;
    wire dcache_tlb_mpu_ppn_barrier_io_y_eff;
    wire dcache_tlb_mpu_ppn_barrier_io_y_c;
    wire dcache_tlb_mpu_ppn_barrier_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_clock;
    wire dcache_tlb_entries_barrier_reset;
    wire[19:0] dcache_tlb_entries_barrier_io_x_ppn;
    wire dcache_tlb_entries_barrier_io_x_u;
    wire dcache_tlb_entries_barrier_io_x_g;
    wire dcache_tlb_entries_barrier_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_io_x_ae_final;
    wire dcache_tlb_entries_barrier_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_io_x_pf;
    wire dcache_tlb_entries_barrier_io_x_gf;
    wire dcache_tlb_entries_barrier_io_x_sw;
    wire dcache_tlb_entries_barrier_io_x_sx;
    wire dcache_tlb_entries_barrier_io_x_sr;
    wire dcache_tlb_entries_barrier_io_x_hw;
    wire dcache_tlb_entries_barrier_io_x_hx;
    wire dcache_tlb_entries_barrier_io_x_hr;
    wire dcache_tlb_entries_barrier_io_x_pw;
    wire dcache_tlb_entries_barrier_io_x_px;
    wire dcache_tlb_entries_barrier_io_x_pr;
    wire dcache_tlb_entries_barrier_io_x_ppp;
    wire dcache_tlb_entries_barrier_io_x_pal;
    wire dcache_tlb_entries_barrier_io_x_paa;
    wire dcache_tlb_entries_barrier_io_x_eff;
    wire dcache_tlb_entries_barrier_io_x_c;
    wire dcache_tlb_entries_barrier_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_io_y_ppn;
    wire dcache_tlb_entries_barrier_io_y_u;
    wire dcache_tlb_entries_barrier_io_y_g;
    wire dcache_tlb_entries_barrier_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_io_y_ae_final;
    wire dcache_tlb_entries_barrier_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_io_y_pf;
    wire dcache_tlb_entries_barrier_io_y_gf;
    wire dcache_tlb_entries_barrier_io_y_sw;
    wire dcache_tlb_entries_barrier_io_y_sx;
    wire dcache_tlb_entries_barrier_io_y_sr;
    wire dcache_tlb_entries_barrier_io_y_hw;
    wire dcache_tlb_entries_barrier_io_y_hx;
    wire dcache_tlb_entries_barrier_io_y_hr;
    wire dcache_tlb_entries_barrier_io_y_pw;
    wire dcache_tlb_entries_barrier_io_y_px;
    wire dcache_tlb_entries_barrier_io_y_pr;
    wire dcache_tlb_entries_barrier_io_y_ppp;
    wire dcache_tlb_entries_barrier_io_y_pal;
    wire dcache_tlb_entries_barrier_io_y_paa;
    wire dcache_tlb_entries_barrier_io_y_eff;
    wire dcache_tlb_entries_barrier_io_y_c;
    wire dcache_tlb_entries_barrier_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_1_clock;
    wire dcache_tlb_entries_barrier_1_reset;
    wire[19:0] dcache_tlb_entries_barrier_1_io_x_ppn;
    wire dcache_tlb_entries_barrier_1_io_x_u;
    wire dcache_tlb_entries_barrier_1_io_x_g;
    wire dcache_tlb_entries_barrier_1_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_1_io_x_ae_final;
    wire dcache_tlb_entries_barrier_1_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_1_io_x_pf;
    wire dcache_tlb_entries_barrier_1_io_x_gf;
    wire dcache_tlb_entries_barrier_1_io_x_sw;
    wire dcache_tlb_entries_barrier_1_io_x_sx;
    wire dcache_tlb_entries_barrier_1_io_x_sr;
    wire dcache_tlb_entries_barrier_1_io_x_hw;
    wire dcache_tlb_entries_barrier_1_io_x_hx;
    wire dcache_tlb_entries_barrier_1_io_x_hr;
    wire dcache_tlb_entries_barrier_1_io_x_pw;
    wire dcache_tlb_entries_barrier_1_io_x_px;
    wire dcache_tlb_entries_barrier_1_io_x_pr;
    wire dcache_tlb_entries_barrier_1_io_x_ppp;
    wire dcache_tlb_entries_barrier_1_io_x_pal;
    wire dcache_tlb_entries_barrier_1_io_x_paa;
    wire dcache_tlb_entries_barrier_1_io_x_eff;
    wire dcache_tlb_entries_barrier_1_io_x_c;
    wire dcache_tlb_entries_barrier_1_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_1_io_y_ppn;
    wire dcache_tlb_entries_barrier_1_io_y_u;
    wire dcache_tlb_entries_barrier_1_io_y_g;
    wire dcache_tlb_entries_barrier_1_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_1_io_y_ae_final;
    wire dcache_tlb_entries_barrier_1_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_1_io_y_pf;
    wire dcache_tlb_entries_barrier_1_io_y_gf;
    wire dcache_tlb_entries_barrier_1_io_y_sw;
    wire dcache_tlb_entries_barrier_1_io_y_sx;
    wire dcache_tlb_entries_barrier_1_io_y_sr;
    wire dcache_tlb_entries_barrier_1_io_y_hw;
    wire dcache_tlb_entries_barrier_1_io_y_hx;
    wire dcache_tlb_entries_barrier_1_io_y_hr;
    wire dcache_tlb_entries_barrier_1_io_y_pw;
    wire dcache_tlb_entries_barrier_1_io_y_px;
    wire dcache_tlb_entries_barrier_1_io_y_pr;
    wire dcache_tlb_entries_barrier_1_io_y_ppp;
    wire dcache_tlb_entries_barrier_1_io_y_pal;
    wire dcache_tlb_entries_barrier_1_io_y_paa;
    wire dcache_tlb_entries_barrier_1_io_y_eff;
    wire dcache_tlb_entries_barrier_1_io_y_c;
    wire dcache_tlb_entries_barrier_1_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_2_clock;
    wire dcache_tlb_entries_barrier_2_reset;
    wire[19:0] dcache_tlb_entries_barrier_2_io_x_ppn;
    wire dcache_tlb_entries_barrier_2_io_x_u;
    wire dcache_tlb_entries_barrier_2_io_x_g;
    wire dcache_tlb_entries_barrier_2_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_2_io_x_ae_final;
    wire dcache_tlb_entries_barrier_2_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_2_io_x_pf;
    wire dcache_tlb_entries_barrier_2_io_x_gf;
    wire dcache_tlb_entries_barrier_2_io_x_sw;
    wire dcache_tlb_entries_barrier_2_io_x_sx;
    wire dcache_tlb_entries_barrier_2_io_x_sr;
    wire dcache_tlb_entries_barrier_2_io_x_hw;
    wire dcache_tlb_entries_barrier_2_io_x_hx;
    wire dcache_tlb_entries_barrier_2_io_x_hr;
    wire dcache_tlb_entries_barrier_2_io_x_pw;
    wire dcache_tlb_entries_barrier_2_io_x_px;
    wire dcache_tlb_entries_barrier_2_io_x_pr;
    wire dcache_tlb_entries_barrier_2_io_x_ppp;
    wire dcache_tlb_entries_barrier_2_io_x_pal;
    wire dcache_tlb_entries_barrier_2_io_x_paa;
    wire dcache_tlb_entries_barrier_2_io_x_eff;
    wire dcache_tlb_entries_barrier_2_io_x_c;
    wire dcache_tlb_entries_barrier_2_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_2_io_y_ppn;
    wire dcache_tlb_entries_barrier_2_io_y_u;
    wire dcache_tlb_entries_barrier_2_io_y_g;
    wire dcache_tlb_entries_barrier_2_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_2_io_y_ae_final;
    wire dcache_tlb_entries_barrier_2_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_2_io_y_pf;
    wire dcache_tlb_entries_barrier_2_io_y_gf;
    wire dcache_tlb_entries_barrier_2_io_y_sw;
    wire dcache_tlb_entries_barrier_2_io_y_sx;
    wire dcache_tlb_entries_barrier_2_io_y_sr;
    wire dcache_tlb_entries_barrier_2_io_y_hw;
    wire dcache_tlb_entries_barrier_2_io_y_hx;
    wire dcache_tlb_entries_barrier_2_io_y_hr;
    wire dcache_tlb_entries_barrier_2_io_y_pw;
    wire dcache_tlb_entries_barrier_2_io_y_px;
    wire dcache_tlb_entries_barrier_2_io_y_pr;
    wire dcache_tlb_entries_barrier_2_io_y_ppp;
    wire dcache_tlb_entries_barrier_2_io_y_pal;
    wire dcache_tlb_entries_barrier_2_io_y_paa;
    wire dcache_tlb_entries_barrier_2_io_y_eff;
    wire dcache_tlb_entries_barrier_2_io_y_c;
    wire dcache_tlb_entries_barrier_2_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_3_clock;
    wire dcache_tlb_entries_barrier_3_reset;
    wire[19:0] dcache_tlb_entries_barrier_3_io_x_ppn;
    wire dcache_tlb_entries_barrier_3_io_x_u;
    wire dcache_tlb_entries_barrier_3_io_x_g;
    wire dcache_tlb_entries_barrier_3_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_3_io_x_ae_final;
    wire dcache_tlb_entries_barrier_3_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_3_io_x_pf;
    wire dcache_tlb_entries_barrier_3_io_x_gf;
    wire dcache_tlb_entries_barrier_3_io_x_sw;
    wire dcache_tlb_entries_barrier_3_io_x_sx;
    wire dcache_tlb_entries_barrier_3_io_x_sr;
    wire dcache_tlb_entries_barrier_3_io_x_hw;
    wire dcache_tlb_entries_barrier_3_io_x_hx;
    wire dcache_tlb_entries_barrier_3_io_x_hr;
    wire dcache_tlb_entries_barrier_3_io_x_pw;
    wire dcache_tlb_entries_barrier_3_io_x_px;
    wire dcache_tlb_entries_barrier_3_io_x_pr;
    wire dcache_tlb_entries_barrier_3_io_x_ppp;
    wire dcache_tlb_entries_barrier_3_io_x_pal;
    wire dcache_tlb_entries_barrier_3_io_x_paa;
    wire dcache_tlb_entries_barrier_3_io_x_eff;
    wire dcache_tlb_entries_barrier_3_io_x_c;
    wire dcache_tlb_entries_barrier_3_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_3_io_y_ppn;
    wire dcache_tlb_entries_barrier_3_io_y_u;
    wire dcache_tlb_entries_barrier_3_io_y_g;
    wire dcache_tlb_entries_barrier_3_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_3_io_y_ae_final;
    wire dcache_tlb_entries_barrier_3_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_3_io_y_pf;
    wire dcache_tlb_entries_barrier_3_io_y_gf;
    wire dcache_tlb_entries_barrier_3_io_y_sw;
    wire dcache_tlb_entries_barrier_3_io_y_sx;
    wire dcache_tlb_entries_barrier_3_io_y_sr;
    wire dcache_tlb_entries_barrier_3_io_y_hw;
    wire dcache_tlb_entries_barrier_3_io_y_hx;
    wire dcache_tlb_entries_barrier_3_io_y_hr;
    wire dcache_tlb_entries_barrier_3_io_y_pw;
    wire dcache_tlb_entries_barrier_3_io_y_px;
    wire dcache_tlb_entries_barrier_3_io_y_pr;
    wire dcache_tlb_entries_barrier_3_io_y_ppp;
    wire dcache_tlb_entries_barrier_3_io_y_pal;
    wire dcache_tlb_entries_barrier_3_io_y_paa;
    wire dcache_tlb_entries_barrier_3_io_y_eff;
    wire dcache_tlb_entries_barrier_3_io_y_c;
    wire dcache_tlb_entries_barrier_3_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_4_clock;
    wire dcache_tlb_entries_barrier_4_reset;
    wire[19:0] dcache_tlb_entries_barrier_4_io_x_ppn;
    wire dcache_tlb_entries_barrier_4_io_x_u;
    wire dcache_tlb_entries_barrier_4_io_x_g;
    wire dcache_tlb_entries_barrier_4_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_4_io_x_ae_final;
    wire dcache_tlb_entries_barrier_4_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_4_io_x_pf;
    wire dcache_tlb_entries_barrier_4_io_x_gf;
    wire dcache_tlb_entries_barrier_4_io_x_sw;
    wire dcache_tlb_entries_barrier_4_io_x_sx;
    wire dcache_tlb_entries_barrier_4_io_x_sr;
    wire dcache_tlb_entries_barrier_4_io_x_hw;
    wire dcache_tlb_entries_barrier_4_io_x_hx;
    wire dcache_tlb_entries_barrier_4_io_x_hr;
    wire dcache_tlb_entries_barrier_4_io_x_pw;
    wire dcache_tlb_entries_barrier_4_io_x_px;
    wire dcache_tlb_entries_barrier_4_io_x_pr;
    wire dcache_tlb_entries_barrier_4_io_x_ppp;
    wire dcache_tlb_entries_barrier_4_io_x_pal;
    wire dcache_tlb_entries_barrier_4_io_x_paa;
    wire dcache_tlb_entries_barrier_4_io_x_eff;
    wire dcache_tlb_entries_barrier_4_io_x_c;
    wire dcache_tlb_entries_barrier_4_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_4_io_y_ppn;
    wire dcache_tlb_entries_barrier_4_io_y_u;
    wire dcache_tlb_entries_barrier_4_io_y_g;
    wire dcache_tlb_entries_barrier_4_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_4_io_y_ae_final;
    wire dcache_tlb_entries_barrier_4_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_4_io_y_pf;
    wire dcache_tlb_entries_barrier_4_io_y_gf;
    wire dcache_tlb_entries_barrier_4_io_y_sw;
    wire dcache_tlb_entries_barrier_4_io_y_sx;
    wire dcache_tlb_entries_barrier_4_io_y_sr;
    wire dcache_tlb_entries_barrier_4_io_y_hw;
    wire dcache_tlb_entries_barrier_4_io_y_hx;
    wire dcache_tlb_entries_barrier_4_io_y_hr;
    wire dcache_tlb_entries_barrier_4_io_y_pw;
    wire dcache_tlb_entries_barrier_4_io_y_px;
    wire dcache_tlb_entries_barrier_4_io_y_pr;
    wire dcache_tlb_entries_barrier_4_io_y_ppp;
    wire dcache_tlb_entries_barrier_4_io_y_pal;
    wire dcache_tlb_entries_barrier_4_io_y_paa;
    wire dcache_tlb_entries_barrier_4_io_y_eff;
    wire dcache_tlb_entries_barrier_4_io_y_c;
    wire dcache_tlb_entries_barrier_4_io_y_fragmented_superpage;
    wire dcache_tlb_entries_barrier_5_clock;
    wire dcache_tlb_entries_barrier_5_reset;
    wire[19:0] dcache_tlb_entries_barrier_5_io_x_ppn;
    wire dcache_tlb_entries_barrier_5_io_x_u;
    wire dcache_tlb_entries_barrier_5_io_x_g;
    wire dcache_tlb_entries_barrier_5_io_x_ae_ptw;
    wire dcache_tlb_entries_barrier_5_io_x_ae_final;
    wire dcache_tlb_entries_barrier_5_io_x_ae_stage2;
    wire dcache_tlb_entries_barrier_5_io_x_pf;
    wire dcache_tlb_entries_barrier_5_io_x_gf;
    wire dcache_tlb_entries_barrier_5_io_x_sw;
    wire dcache_tlb_entries_barrier_5_io_x_sx;
    wire dcache_tlb_entries_barrier_5_io_x_sr;
    wire dcache_tlb_entries_barrier_5_io_x_hw;
    wire dcache_tlb_entries_barrier_5_io_x_hx;
    wire dcache_tlb_entries_barrier_5_io_x_hr;
    wire dcache_tlb_entries_barrier_5_io_x_pw;
    wire dcache_tlb_entries_barrier_5_io_x_px;
    wire dcache_tlb_entries_barrier_5_io_x_pr;
    wire dcache_tlb_entries_barrier_5_io_x_ppp;
    wire dcache_tlb_entries_barrier_5_io_x_pal;
    wire dcache_tlb_entries_barrier_5_io_x_paa;
    wire dcache_tlb_entries_barrier_5_io_x_eff;
    wire dcache_tlb_entries_barrier_5_io_x_c;
    wire dcache_tlb_entries_barrier_5_io_x_fragmented_superpage;
    wire[19:0] dcache_tlb_entries_barrier_5_io_y_ppn;
    wire dcache_tlb_entries_barrier_5_io_y_u;
    wire dcache_tlb_entries_barrier_5_io_y_g;
    wire dcache_tlb_entries_barrier_5_io_y_ae_ptw;
    wire dcache_tlb_entries_barrier_5_io_y_ae_final;
    wire dcache_tlb_entries_barrier_5_io_y_ae_stage2;
    wire dcache_tlb_entries_barrier_5_io_y_pf;
    wire dcache_tlb_entries_barrier_5_io_y_gf;
    wire dcache_tlb_entries_barrier_5_io_y_sw;
    wire dcache_tlb_entries_barrier_5_io_y_sx;
    wire dcache_tlb_entries_barrier_5_io_y_sr;
    wire dcache_tlb_entries_barrier_5_io_y_hw;
    wire dcache_tlb_entries_barrier_5_io_y_hx;
    wire dcache_tlb_entries_barrier_5_io_y_hr;
    wire dcache_tlb_entries_barrier_5_io_y_pw;
    wire dcache_tlb_entries_barrier_5_io_y_px;
    wire dcache_tlb_entries_barrier_5_io_y_pr;
    wire dcache_tlb_entries_barrier_5_io_y_ppp;
    wire dcache_tlb_entries_barrier_5_io_y_pal;
    wire dcache_tlb_entries_barrier_5_io_y_paa;
    wire dcache_tlb_entries_barrier_5_io_y_eff;
    wire dcache_tlb_entries_barrier_5_io_y_c;
    wire dcache_tlb_entries_barrier_5_io_y_fragmented_superpage;
    wire dcache_pma_checker_mpu_ppn_barrier_clock;
    wire dcache_pma_checker_mpu_ppn_barrier_reset;
    wire[19:0] dcache_pma_checker_mpu_ppn_barrier_io_x_ppn;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_u;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_g;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_ae_ptw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_ae_final;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_ae_stage2;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_pf;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_gf;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_sw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_sx;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_sr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_hw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_hx;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_hr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_pw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_px;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_pr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_ppp;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_pal;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_paa;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_eff;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_c;
    wire dcache_pma_checker_mpu_ppn_barrier_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_mpu_ppn_barrier_io_y_ppn;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_u;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_g;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_ae_ptw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_ae_final;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_ae_stage2;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_pf;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_gf;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_sw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_sx;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_sr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_hw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_hx;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_hr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_pw;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_px;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_pr;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_ppp;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_pal;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_paa;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_eff;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_c;
    wire dcache_pma_checker_mpu_ppn_barrier_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_clock;
    wire dcache_pma_checker_entries_barrier_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_io_x_u;
    wire dcache_pma_checker_entries_barrier_io_x_g;
    wire dcache_pma_checker_entries_barrier_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_io_x_pf;
    wire dcache_pma_checker_entries_barrier_io_x_gf;
    wire dcache_pma_checker_entries_barrier_io_x_sw;
    wire dcache_pma_checker_entries_barrier_io_x_sx;
    wire dcache_pma_checker_entries_barrier_io_x_sr;
    wire dcache_pma_checker_entries_barrier_io_x_hw;
    wire dcache_pma_checker_entries_barrier_io_x_hx;
    wire dcache_pma_checker_entries_barrier_io_x_hr;
    wire dcache_pma_checker_entries_barrier_io_x_pw;
    wire dcache_pma_checker_entries_barrier_io_x_px;
    wire dcache_pma_checker_entries_barrier_io_x_pr;
    wire dcache_pma_checker_entries_barrier_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_io_x_pal;
    wire dcache_pma_checker_entries_barrier_io_x_paa;
    wire dcache_pma_checker_entries_barrier_io_x_eff;
    wire dcache_pma_checker_entries_barrier_io_x_c;
    wire dcache_pma_checker_entries_barrier_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_io_y_u;
    wire dcache_pma_checker_entries_barrier_io_y_g;
    wire dcache_pma_checker_entries_barrier_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_io_y_pf;
    wire dcache_pma_checker_entries_barrier_io_y_gf;
    wire dcache_pma_checker_entries_barrier_io_y_sw;
    wire dcache_pma_checker_entries_barrier_io_y_sx;
    wire dcache_pma_checker_entries_barrier_io_y_sr;
    wire dcache_pma_checker_entries_barrier_io_y_hw;
    wire dcache_pma_checker_entries_barrier_io_y_hx;
    wire dcache_pma_checker_entries_barrier_io_y_hr;
    wire dcache_pma_checker_entries_barrier_io_y_pw;
    wire dcache_pma_checker_entries_barrier_io_y_px;
    wire dcache_pma_checker_entries_barrier_io_y_pr;
    wire dcache_pma_checker_entries_barrier_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_io_y_pal;
    wire dcache_pma_checker_entries_barrier_io_y_paa;
    wire dcache_pma_checker_entries_barrier_io_y_eff;
    wire dcache_pma_checker_entries_barrier_io_y_c;
    wire dcache_pma_checker_entries_barrier_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_1_clock;
    wire dcache_pma_checker_entries_barrier_1_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_1_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_1_io_x_u;
    wire dcache_pma_checker_entries_barrier_1_io_x_g;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_1_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_1_io_x_pf;
    wire dcache_pma_checker_entries_barrier_1_io_x_gf;
    wire dcache_pma_checker_entries_barrier_1_io_x_sw;
    wire dcache_pma_checker_entries_barrier_1_io_x_sx;
    wire dcache_pma_checker_entries_barrier_1_io_x_sr;
    wire dcache_pma_checker_entries_barrier_1_io_x_hw;
    wire dcache_pma_checker_entries_barrier_1_io_x_hx;
    wire dcache_pma_checker_entries_barrier_1_io_x_hr;
    wire dcache_pma_checker_entries_barrier_1_io_x_pw;
    wire dcache_pma_checker_entries_barrier_1_io_x_px;
    wire dcache_pma_checker_entries_barrier_1_io_x_pr;
    wire dcache_pma_checker_entries_barrier_1_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_1_io_x_pal;
    wire dcache_pma_checker_entries_barrier_1_io_x_paa;
    wire dcache_pma_checker_entries_barrier_1_io_x_eff;
    wire dcache_pma_checker_entries_barrier_1_io_x_c;
    wire dcache_pma_checker_entries_barrier_1_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_1_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_1_io_y_u;
    wire dcache_pma_checker_entries_barrier_1_io_y_g;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_1_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_1_io_y_pf;
    wire dcache_pma_checker_entries_barrier_1_io_y_gf;
    wire dcache_pma_checker_entries_barrier_1_io_y_sw;
    wire dcache_pma_checker_entries_barrier_1_io_y_sx;
    wire dcache_pma_checker_entries_barrier_1_io_y_sr;
    wire dcache_pma_checker_entries_barrier_1_io_y_hw;
    wire dcache_pma_checker_entries_barrier_1_io_y_hx;
    wire dcache_pma_checker_entries_barrier_1_io_y_hr;
    wire dcache_pma_checker_entries_barrier_1_io_y_pw;
    wire dcache_pma_checker_entries_barrier_1_io_y_px;
    wire dcache_pma_checker_entries_barrier_1_io_y_pr;
    wire dcache_pma_checker_entries_barrier_1_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_1_io_y_pal;
    wire dcache_pma_checker_entries_barrier_1_io_y_paa;
    wire dcache_pma_checker_entries_barrier_1_io_y_eff;
    wire dcache_pma_checker_entries_barrier_1_io_y_c;
    wire dcache_pma_checker_entries_barrier_1_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_2_clock;
    wire dcache_pma_checker_entries_barrier_2_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_2_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_2_io_x_u;
    wire dcache_pma_checker_entries_barrier_2_io_x_g;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_2_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_2_io_x_pf;
    wire dcache_pma_checker_entries_barrier_2_io_x_gf;
    wire dcache_pma_checker_entries_barrier_2_io_x_sw;
    wire dcache_pma_checker_entries_barrier_2_io_x_sx;
    wire dcache_pma_checker_entries_barrier_2_io_x_sr;
    wire dcache_pma_checker_entries_barrier_2_io_x_hw;
    wire dcache_pma_checker_entries_barrier_2_io_x_hx;
    wire dcache_pma_checker_entries_barrier_2_io_x_hr;
    wire dcache_pma_checker_entries_barrier_2_io_x_pw;
    wire dcache_pma_checker_entries_barrier_2_io_x_px;
    wire dcache_pma_checker_entries_barrier_2_io_x_pr;
    wire dcache_pma_checker_entries_barrier_2_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_2_io_x_pal;
    wire dcache_pma_checker_entries_barrier_2_io_x_paa;
    wire dcache_pma_checker_entries_barrier_2_io_x_eff;
    wire dcache_pma_checker_entries_barrier_2_io_x_c;
    wire dcache_pma_checker_entries_barrier_2_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_2_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_2_io_y_u;
    wire dcache_pma_checker_entries_barrier_2_io_y_g;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_2_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_2_io_y_pf;
    wire dcache_pma_checker_entries_barrier_2_io_y_gf;
    wire dcache_pma_checker_entries_barrier_2_io_y_sw;
    wire dcache_pma_checker_entries_barrier_2_io_y_sx;
    wire dcache_pma_checker_entries_barrier_2_io_y_sr;
    wire dcache_pma_checker_entries_barrier_2_io_y_hw;
    wire dcache_pma_checker_entries_barrier_2_io_y_hx;
    wire dcache_pma_checker_entries_barrier_2_io_y_hr;
    wire dcache_pma_checker_entries_barrier_2_io_y_pw;
    wire dcache_pma_checker_entries_barrier_2_io_y_px;
    wire dcache_pma_checker_entries_barrier_2_io_y_pr;
    wire dcache_pma_checker_entries_barrier_2_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_2_io_y_pal;
    wire dcache_pma_checker_entries_barrier_2_io_y_paa;
    wire dcache_pma_checker_entries_barrier_2_io_y_eff;
    wire dcache_pma_checker_entries_barrier_2_io_y_c;
    wire dcache_pma_checker_entries_barrier_2_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_3_clock;
    wire dcache_pma_checker_entries_barrier_3_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_3_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_3_io_x_u;
    wire dcache_pma_checker_entries_barrier_3_io_x_g;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_3_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_3_io_x_pf;
    wire dcache_pma_checker_entries_barrier_3_io_x_gf;
    wire dcache_pma_checker_entries_barrier_3_io_x_sw;
    wire dcache_pma_checker_entries_barrier_3_io_x_sx;
    wire dcache_pma_checker_entries_barrier_3_io_x_sr;
    wire dcache_pma_checker_entries_barrier_3_io_x_hw;
    wire dcache_pma_checker_entries_barrier_3_io_x_hx;
    wire dcache_pma_checker_entries_barrier_3_io_x_hr;
    wire dcache_pma_checker_entries_barrier_3_io_x_pw;
    wire dcache_pma_checker_entries_barrier_3_io_x_px;
    wire dcache_pma_checker_entries_barrier_3_io_x_pr;
    wire dcache_pma_checker_entries_barrier_3_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_3_io_x_pal;
    wire dcache_pma_checker_entries_barrier_3_io_x_paa;
    wire dcache_pma_checker_entries_barrier_3_io_x_eff;
    wire dcache_pma_checker_entries_barrier_3_io_x_c;
    wire dcache_pma_checker_entries_barrier_3_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_3_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_3_io_y_u;
    wire dcache_pma_checker_entries_barrier_3_io_y_g;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_3_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_3_io_y_pf;
    wire dcache_pma_checker_entries_barrier_3_io_y_gf;
    wire dcache_pma_checker_entries_barrier_3_io_y_sw;
    wire dcache_pma_checker_entries_barrier_3_io_y_sx;
    wire dcache_pma_checker_entries_barrier_3_io_y_sr;
    wire dcache_pma_checker_entries_barrier_3_io_y_hw;
    wire dcache_pma_checker_entries_barrier_3_io_y_hx;
    wire dcache_pma_checker_entries_barrier_3_io_y_hr;
    wire dcache_pma_checker_entries_barrier_3_io_y_pw;
    wire dcache_pma_checker_entries_barrier_3_io_y_px;
    wire dcache_pma_checker_entries_barrier_3_io_y_pr;
    wire dcache_pma_checker_entries_barrier_3_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_3_io_y_pal;
    wire dcache_pma_checker_entries_barrier_3_io_y_paa;
    wire dcache_pma_checker_entries_barrier_3_io_y_eff;
    wire dcache_pma_checker_entries_barrier_3_io_y_c;
    wire dcache_pma_checker_entries_barrier_3_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_4_clock;
    wire dcache_pma_checker_entries_barrier_4_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_4_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_4_io_x_u;
    wire dcache_pma_checker_entries_barrier_4_io_x_g;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_4_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_4_io_x_pf;
    wire dcache_pma_checker_entries_barrier_4_io_x_gf;
    wire dcache_pma_checker_entries_barrier_4_io_x_sw;
    wire dcache_pma_checker_entries_barrier_4_io_x_sx;
    wire dcache_pma_checker_entries_barrier_4_io_x_sr;
    wire dcache_pma_checker_entries_barrier_4_io_x_hw;
    wire dcache_pma_checker_entries_barrier_4_io_x_hx;
    wire dcache_pma_checker_entries_barrier_4_io_x_hr;
    wire dcache_pma_checker_entries_barrier_4_io_x_pw;
    wire dcache_pma_checker_entries_barrier_4_io_x_px;
    wire dcache_pma_checker_entries_barrier_4_io_x_pr;
    wire dcache_pma_checker_entries_barrier_4_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_4_io_x_pal;
    wire dcache_pma_checker_entries_barrier_4_io_x_paa;
    wire dcache_pma_checker_entries_barrier_4_io_x_eff;
    wire dcache_pma_checker_entries_barrier_4_io_x_c;
    wire dcache_pma_checker_entries_barrier_4_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_4_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_4_io_y_u;
    wire dcache_pma_checker_entries_barrier_4_io_y_g;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_4_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_4_io_y_pf;
    wire dcache_pma_checker_entries_barrier_4_io_y_gf;
    wire dcache_pma_checker_entries_barrier_4_io_y_sw;
    wire dcache_pma_checker_entries_barrier_4_io_y_sx;
    wire dcache_pma_checker_entries_barrier_4_io_y_sr;
    wire dcache_pma_checker_entries_barrier_4_io_y_hw;
    wire dcache_pma_checker_entries_barrier_4_io_y_hx;
    wire dcache_pma_checker_entries_barrier_4_io_y_hr;
    wire dcache_pma_checker_entries_barrier_4_io_y_pw;
    wire dcache_pma_checker_entries_barrier_4_io_y_px;
    wire dcache_pma_checker_entries_barrier_4_io_y_pr;
    wire dcache_pma_checker_entries_barrier_4_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_4_io_y_pal;
    wire dcache_pma_checker_entries_barrier_4_io_y_paa;
    wire dcache_pma_checker_entries_barrier_4_io_y_eff;
    wire dcache_pma_checker_entries_barrier_4_io_y_c;
    wire dcache_pma_checker_entries_barrier_4_io_y_fragmented_superpage;
    wire dcache_pma_checker_entries_barrier_5_clock;
    wire dcache_pma_checker_entries_barrier_5_reset;
    wire[19:0] dcache_pma_checker_entries_barrier_5_io_x_ppn;
    wire dcache_pma_checker_entries_barrier_5_io_x_u;
    wire dcache_pma_checker_entries_barrier_5_io_x_g;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_ptw;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_final;
    wire dcache_pma_checker_entries_barrier_5_io_x_ae_stage2;
    wire dcache_pma_checker_entries_barrier_5_io_x_pf;
    wire dcache_pma_checker_entries_barrier_5_io_x_gf;
    wire dcache_pma_checker_entries_barrier_5_io_x_sw;
    wire dcache_pma_checker_entries_barrier_5_io_x_sx;
    wire dcache_pma_checker_entries_barrier_5_io_x_sr;
    wire dcache_pma_checker_entries_barrier_5_io_x_hw;
    wire dcache_pma_checker_entries_barrier_5_io_x_hx;
    wire dcache_pma_checker_entries_barrier_5_io_x_hr;
    wire dcache_pma_checker_entries_barrier_5_io_x_pw;
    wire dcache_pma_checker_entries_barrier_5_io_x_px;
    wire dcache_pma_checker_entries_barrier_5_io_x_pr;
    wire dcache_pma_checker_entries_barrier_5_io_x_ppp;
    wire dcache_pma_checker_entries_barrier_5_io_x_pal;
    wire dcache_pma_checker_entries_barrier_5_io_x_paa;
    wire dcache_pma_checker_entries_barrier_5_io_x_eff;
    wire dcache_pma_checker_entries_barrier_5_io_x_c;
    wire dcache_pma_checker_entries_barrier_5_io_x_fragmented_superpage;
    wire[19:0] dcache_pma_checker_entries_barrier_5_io_y_ppn;
    wire dcache_pma_checker_entries_barrier_5_io_y_u;
    wire dcache_pma_checker_entries_barrier_5_io_y_g;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_ptw;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_final;
    wire dcache_pma_checker_entries_barrier_5_io_y_ae_stage2;
    wire dcache_pma_checker_entries_barrier_5_io_y_pf;
    wire dcache_pma_checker_entries_barrier_5_io_y_gf;
    wire dcache_pma_checker_entries_barrier_5_io_y_sw;
    wire dcache_pma_checker_entries_barrier_5_io_y_sx;
    wire dcache_pma_checker_entries_barrier_5_io_y_sr;
    wire dcache_pma_checker_entries_barrier_5_io_y_hw;
    wire dcache_pma_checker_entries_barrier_5_io_y_hx;
    wire dcache_pma_checker_entries_barrier_5_io_y_hr;
    wire dcache_pma_checker_entries_barrier_5_io_y_pw;
    wire dcache_pma_checker_entries_barrier_5_io_y_px;
    wire dcache_pma_checker_entries_barrier_5_io_y_pr;
    wire dcache_pma_checker_entries_barrier_5_io_y_ppp;
    wire dcache_pma_checker_entries_barrier_5_io_y_pal;
    wire dcache_pma_checker_entries_barrier_5_io_y_paa;
    wire dcache_pma_checker_entries_barrier_5_io_y_eff;
    wire dcache_pma_checker_entries_barrier_5_io_y_c;
    wire dcache_pma_checker_entries_barrier_5_io_y_fragmented_superpage;

    assign  dcache_tlb_mpu_ppn_barrier_io_y_ppn = dcache_tlb_mpu_ppn_barrier_io_x_ppn ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_u = dcache_tlb_mpu_ppn_barrier_io_x_u ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_g = dcache_tlb_mpu_ppn_barrier_io_x_g ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_ae_ptw = dcache_tlb_mpu_ppn_barrier_io_x_ae_ptw ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_ae_final = dcache_tlb_mpu_ppn_barrier_io_x_ae_final ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_ae_stage2 = dcache_tlb_mpu_ppn_barrier_io_x_ae_stage2 ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_pf = dcache_tlb_mpu_ppn_barrier_io_x_pf ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_gf = dcache_tlb_mpu_ppn_barrier_io_x_gf ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_sw = dcache_tlb_mpu_ppn_barrier_io_x_sw ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_sx = dcache_tlb_mpu_ppn_barrier_io_x_sx ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_sr = dcache_tlb_mpu_ppn_barrier_io_x_sr ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_hw = dcache_tlb_mpu_ppn_barrier_io_x_hw ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_hx = dcache_tlb_mpu_ppn_barrier_io_x_hx ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_hr = dcache_tlb_mpu_ppn_barrier_io_x_hr ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_pw = dcache_tlb_mpu_ppn_barrier_io_x_pw ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_px = dcache_tlb_mpu_ppn_barrier_io_x_px ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_pr = dcache_tlb_mpu_ppn_barrier_io_x_pr ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_ppp = dcache_tlb_mpu_ppn_barrier_io_x_ppp ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_pal = dcache_tlb_mpu_ppn_barrier_io_x_pal ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_paa = dcache_tlb_mpu_ppn_barrier_io_x_paa ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_eff = dcache_tlb_mpu_ppn_barrier_io_x_eff ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_c = dcache_tlb_mpu_ppn_barrier_io_x_c ; 
  assign  dcache_tlb_mpu_ppn_barrier_io_y_fragmented_superpage = dcache_tlb_mpu_ppn_barrier_io_x_fragmented_superpage ;
     
    wire[21:0] dcache_tlb_mpu_ppn = dcache_tlb_do_refill  ? {2'h0, dcache_tlb_refill_ppn }: dcache_tlb_vm_enabled  ? {2'h0, dcache__tlb_mpu_ppn_barrier_io_y_ppn }: dcache_tlb_io_req_bits_vaddr [33:12]; 
    wire[33:0] dcache_tlb_mpu_physaddr ={ dcache_tlb_mpu_ppn , dcache_tlb_io_req_bits_vaddr [11:0]}; 
    wire[2:0] dcache_tlb_mpu_priv ={ dcache_tlb_io_ptw_status_debug , dcache_tlb_io_req_bits_prv }; 
    wire[1:0] dcache_tlb_io_req_bits_size ;  
    wire dcache_tlb_pmp_clock;
    wire dcache_tlb_pmp_reset;
    wire[1:0] dcache_tlb_pmp_io_prv;
    wire dcache_tlb_pmp_io_pmp_0_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_0_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_0_cfg_a;
    wire dcache_tlb_pmp_io_pmp_0_cfg_x;
    wire dcache_tlb_pmp_io_pmp_0_cfg_w;
    wire dcache_tlb_pmp_io_pmp_0_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_0_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_0_mask;
    wire dcache_tlb_pmp_io_pmp_1_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_1_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_1_cfg_a;
    wire dcache_tlb_pmp_io_pmp_1_cfg_x;
    wire dcache_tlb_pmp_io_pmp_1_cfg_w;
    wire dcache_tlb_pmp_io_pmp_1_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_1_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_1_mask;
    wire dcache_tlb_pmp_io_pmp_2_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_2_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_2_cfg_a;
    wire dcache_tlb_pmp_io_pmp_2_cfg_x;
    wire dcache_tlb_pmp_io_pmp_2_cfg_w;
    wire dcache_tlb_pmp_io_pmp_2_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_2_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_2_mask;
    wire dcache_tlb_pmp_io_pmp_3_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_3_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_3_cfg_a;
    wire dcache_tlb_pmp_io_pmp_3_cfg_x;
    wire dcache_tlb_pmp_io_pmp_3_cfg_w;
    wire dcache_tlb_pmp_io_pmp_3_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_3_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_3_mask;
    wire dcache_tlb_pmp_io_pmp_4_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_4_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_4_cfg_a;
    wire dcache_tlb_pmp_io_pmp_4_cfg_x;
    wire dcache_tlb_pmp_io_pmp_4_cfg_w;
    wire dcache_tlb_pmp_io_pmp_4_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_4_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_4_mask;
    wire dcache_tlb_pmp_io_pmp_5_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_5_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_5_cfg_a;
    wire dcache_tlb_pmp_io_pmp_5_cfg_x;
    wire dcache_tlb_pmp_io_pmp_5_cfg_w;
    wire dcache_tlb_pmp_io_pmp_5_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_5_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_5_mask;
    wire dcache_tlb_pmp_io_pmp_6_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_6_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_6_cfg_a;
    wire dcache_tlb_pmp_io_pmp_6_cfg_x;
    wire dcache_tlb_pmp_io_pmp_6_cfg_w;
    wire dcache_tlb_pmp_io_pmp_6_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_6_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_6_mask;
    wire dcache_tlb_pmp_io_pmp_7_cfg_l;
    wire[1:0] dcache_tlb_pmp_io_pmp_7_cfg_res;
    wire[1:0] dcache_tlb_pmp_io_pmp_7_cfg_a;
    wire dcache_tlb_pmp_io_pmp_7_cfg_x;
    wire dcache_tlb_pmp_io_pmp_7_cfg_w;
    wire dcache_tlb_pmp_io_pmp_7_cfg_r;
    wire[29:0] dcache_tlb_pmp_io_pmp_7_addr;
    wire[31:0] dcache_tlb_pmp_io_pmp_7_mask;
    wire[31:0] dcache_tlb_pmp_io_addr;
    wire[1:0] dcache_tlb_pmp_io_size;
    wire dcache_tlb_pmp_io_r;
    wire dcache_tlb_pmp_io_w;
    wire dcache_tlb_pmp_io_x;
    wire dcache_pma_checker_pmp_clock;
    wire dcache_pma_checker_pmp_reset;
    wire[1:0] dcache_pma_checker_pmp_io_prv;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_0_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_0_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_0_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_0_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_0_mask;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_1_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_1_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_1_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_1_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_1_mask;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_2_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_2_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_2_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_2_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_2_mask;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_3_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_3_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_3_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_3_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_3_mask;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_4_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_4_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_4_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_4_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_4_mask;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_5_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_5_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_5_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_5_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_5_mask;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_6_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_6_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_6_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_6_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_6_mask;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_l;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_7_cfg_res;
    wire[1:0] dcache_pma_checker_pmp_io_pmp_7_cfg_a;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_x;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_w;
    wire dcache_pma_checker_pmp_io_pmp_7_cfg_r;
    wire[29:0] dcache_pma_checker_pmp_io_pmp_7_addr;
    wire[31:0] dcache_pma_checker_pmp_io_pmp_7_mask;
    wire[31:0] dcache_pma_checker_pmp_io_addr;
    wire[1:0] dcache_pma_checker_pmp_io_size;
    wire dcache_pma_checker_pmp_io_r;
    wire dcache_pma_checker_pmp_io_w;
    wire dcache_pma_checker_pmp_io_x;

    wire dcache_tlb_pmp_res_cur_cfg_l = dcache_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_cfg_res = dcache_tlb_pmp_io_pmp_7_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_cfg_a = dcache_tlb_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_addr = dcache_tlb_pmp_io_pmp_7_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_mask = dcache_tlb_pmp_io_pmp_7_mask ; 
    wire dcache_tlb_pmp_res_cur_1_cfg_l = dcache_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_1_cfg_res = dcache_tlb_pmp_io_pmp_6_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_1_cfg_a = dcache_tlb_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_1_addr = dcache_tlb_pmp_io_pmp_6_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_1_mask = dcache_tlb_pmp_io_pmp_6_mask ; 
    wire dcache_tlb_pmp_res_cur_2_cfg_l = dcache_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_2_cfg_res = dcache_tlb_pmp_io_pmp_5_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_2_cfg_a = dcache_tlb_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_2_addr = dcache_tlb_pmp_io_pmp_5_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_2_mask = dcache_tlb_pmp_io_pmp_5_mask ; 
    wire dcache_tlb_pmp_res_cur_3_cfg_l = dcache_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_3_cfg_res = dcache_tlb_pmp_io_pmp_4_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_3_cfg_a = dcache_tlb_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_3_addr = dcache_tlb_pmp_io_pmp_4_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_3_mask = dcache_tlb_pmp_io_pmp_4_mask ; 
    wire dcache_tlb_pmp_res_cur_4_cfg_l = dcache_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_4_cfg_res = dcache_tlb_pmp_io_pmp_3_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_4_cfg_a = dcache_tlb_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_4_addr = dcache_tlb_pmp_io_pmp_3_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_4_mask = dcache_tlb_pmp_io_pmp_3_mask ; 
    wire dcache_tlb_pmp_res_cur_5_cfg_l = dcache_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_5_cfg_res = dcache_tlb_pmp_io_pmp_2_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_5_cfg_a = dcache_tlb_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_5_addr = dcache_tlb_pmp_io_pmp_2_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_5_mask = dcache_tlb_pmp_io_pmp_2_mask ; 
    wire dcache_tlb_pmp_res_cur_6_cfg_l = dcache_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_6_cfg_res = dcache_tlb_pmp_io_pmp_1_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_6_cfg_a = dcache_tlb_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_6_addr = dcache_tlb_pmp_io_pmp_1_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_6_mask = dcache_tlb_pmp_io_pmp_1_mask ; 
    wire dcache_tlb_pmp_res_cur_7_cfg_l = dcache_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cur_7_cfg_res = dcache_tlb_pmp_io_pmp_0_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cur_7_cfg_a = dcache_tlb_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_res_cur_7_addr = dcache_tlb_pmp_io_pmp_0_addr ; 
    wire[31:0] dcache_tlb_pmp_res_cur_7_mask = dcache_tlb_pmp_io_pmp_0_mask ; 
    wire[1:0] dcache_tlb_pmp__pmp0_WIRE_cfg_res =2'h0; 
    wire[1:0] dcache_tlb_pmp__pmp0_WIRE_cfg_a =2'h0; 
    wire[29:0] dcache_tlb_pmp__pmp0_WIRE_addr =30'h0; 
    wire[31:0] dcache_tlb_pmp__pmp0_WIRE_mask =32'h0; 
    wire dcache_tlb_pmp__pmp0_WIRE_cfg_l =1'h0; 
    wire dcache_tlb_pmp__pmp0_WIRE_cfg_x =1'h0; 
    wire dcache_tlb_pmp__pmp0_WIRE_cfg_w =1'h0; 
    wire dcache_tlb_pmp__pmp0_WIRE_cfg_r =1'h0; 
    wire dcache_tlb_pmp_default_0 = dcache_tlb_pmp_io_prv >2'h1; 
    wire dcache_tlb_pmp_pmp0_cfg_x = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_pmp0_cfg_w = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_pmp0_cfg_r = dcache_tlb_pmp_default_0 ; 
    wire dcache_tlb_pmp_pmp0_cfg_l = dcache_tlb_pmp__pmp0_WIRE_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_pmp0_cfg_res = dcache_tlb_pmp__pmp0_WIRE_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_pmp0_cfg_a = dcache_tlb_pmp__pmp0_WIRE_cfg_a ; 
    wire[29:0] dcache_tlb_pmp_pmp0_addr = dcache_tlb_pmp__pmp0_WIRE_addr ; 
    wire[31:0] dcache_tlb_pmp_pmp0_mask = dcache_tlb_pmp__pmp0_WIRE_mask ; 
    wire[5:0] dcache_tlb_pmp__GEN =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask = dcache_tlb_pmp_io_pmp_7_mask |{29'h0,~( dcache_tlb_pmp__GEN [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_0 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_0 [31:3])&~( dcache_tlb_pmp_io_pmp_7_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_1 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_1 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_2 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_3 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_3 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_4 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_4 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_5 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_2 [2:0]))< dcache_tlb_pmp__GEN_5 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_6 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_1 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_6 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_7 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_1 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_7 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_8 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_1 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_8 [2:0]; 
    wire dcache_tlb_pmp_res_hit = dcache_tlb_pmp_io_pmp_7_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch & dcache_tlb_pmp_res_hit_lsbMatch : dcache_tlb_pmp_io_pmp_7_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess | dcache_tlb_pmp_res_hit_msbsEqual & dcache_tlb_pmp_res_hit_lsbsLess )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_1 | dcache_tlb_pmp_res_hit_msbsEqual_1 & dcache_tlb_pmp_res_hit_lsbsLess_1 ); 
    wire dcache_tlb_pmp_res_ignore = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_7_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_9 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask =~( dcache_tlb_pmp__GEN_9 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_10 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_11 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_10 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_11 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_12 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_13 =~(~{ dcache_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_12 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_13 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned =( dcache_tlb_pmp_res_aligned_straddlesLowerBound | dcache_tlb_pmp_res_aligned_straddlesUpperBound )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned =( dcache_tlb_pmp_res_aligned_lsbMask &~( dcache_tlb_pmp_io_pmp_7_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned = dcache_tlb_pmp_io_pmp_7_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned : dcache_tlb_pmp_res_aligned_rangeAligned ; 
    wire[1:0] dcache_tlb_pmp_res_hi ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_1 ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_2 ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_3 ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_4 ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_5 ={ dcache_tlb_pmp_io_pmp_7_cfg_x , dcache_tlb_pmp_io_pmp_7_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_cfg_r = dcache_tlb_pmp_res_aligned &( dcache_tlb_pmp_io_pmp_7_cfg_r | dcache_tlb_pmp_res_ignore ); 
    wire dcache_tlb_pmp_res_cur_cfg_w = dcache_tlb_pmp_res_aligned &( dcache_tlb_pmp_io_pmp_7_cfg_w | dcache_tlb_pmp_res_ignore ); 
    wire dcache_tlb_pmp_res_cur_cfg_x = dcache_tlb_pmp_res_aligned &( dcache_tlb_pmp_io_pmp_7_cfg_x | dcache_tlb_pmp_res_ignore ); 
    wire[5:0] dcache_tlb_pmp__GEN_14 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_1 = dcache_tlb_pmp_io_pmp_6_mask |{29'h0,~( dcache_tlb_pmp__GEN_14 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_15 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_1 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_15 [31:3])&~( dcache_tlb_pmp_io_pmp_6_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_16 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_1 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_16 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_1 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_17 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_18 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_2 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_18 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_19 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_2 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_19 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_20 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_2 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_17 [2:0]))< dcache_tlb_pmp__GEN_20 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_21 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_3 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_21 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_22 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_3 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_22 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_23 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_3 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_23 [2:0]; 
    wire dcache_tlb_pmp_res_hit_1 = dcache_tlb_pmp_io_pmp_6_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_1 & dcache_tlb_pmp_res_hit_lsbMatch_1 : dcache_tlb_pmp_io_pmp_6_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_2 | dcache_tlb_pmp_res_hit_msbsEqual_2 & dcache_tlb_pmp_res_hit_lsbsLess_2 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_3 | dcache_tlb_pmp_res_hit_msbsEqual_3 & dcache_tlb_pmp_res_hit_lsbsLess_3 ); 
    wire dcache_tlb_pmp_res_ignore_1 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_6_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_24 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_1 =~( dcache_tlb_pmp__GEN_24 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_25 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_26 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_1 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_25 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_26 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_27 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_28 =~(~{ dcache_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_1 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_27 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_28 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_1 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_1 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_1 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_1 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_1 =( dcache_tlb_pmp_res_aligned_lsbMask_1 &~( dcache_tlb_pmp_io_pmp_6_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_1 = dcache_tlb_pmp_io_pmp_6_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_1 : dcache_tlb_pmp_res_aligned_rangeAligned_1 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_6 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_7 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_8 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_9 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_10 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_11 ={ dcache_tlb_pmp_io_pmp_6_cfg_x , dcache_tlb_pmp_io_pmp_6_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_1_cfg_r = dcache_tlb_pmp_res_aligned_1 &( dcache_tlb_pmp_io_pmp_6_cfg_r | dcache_tlb_pmp_res_ignore_1 ); 
    wire dcache_tlb_pmp_res_cur_1_cfg_w = dcache_tlb_pmp_res_aligned_1 &( dcache_tlb_pmp_io_pmp_6_cfg_w | dcache_tlb_pmp_res_ignore_1 ); 
    wire dcache_tlb_pmp_res_cur_1_cfg_x = dcache_tlb_pmp_res_aligned_1 &( dcache_tlb_pmp_io_pmp_6_cfg_x | dcache_tlb_pmp_res_ignore_1 ); 
    wire[5:0] dcache_tlb_pmp__GEN_29 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_2 = dcache_tlb_pmp_io_pmp_5_mask |{29'h0,~( dcache_tlb_pmp__GEN_29 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_30 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_2 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_30 [31:3])&~( dcache_tlb_pmp_io_pmp_5_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_31 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_2 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_31 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_2 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_32 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_33 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_4 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_33 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_34 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_4 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_34 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_35 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_4 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_32 [2:0]))< dcache_tlb_pmp__GEN_35 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_36 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_5 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_36 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_37 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_5 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_37 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_38 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_5 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_38 [2:0]; 
    wire dcache_tlb_pmp_res_hit_2 = dcache_tlb_pmp_io_pmp_5_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_2 & dcache_tlb_pmp_res_hit_lsbMatch_2 : dcache_tlb_pmp_io_pmp_5_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_4 | dcache_tlb_pmp_res_hit_msbsEqual_4 & dcache_tlb_pmp_res_hit_lsbsLess_4 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_5 | dcache_tlb_pmp_res_hit_msbsEqual_5 & dcache_tlb_pmp_res_hit_lsbsLess_5 ); 
    wire dcache_tlb_pmp_res_ignore_2 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_5_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_39 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_2 =~( dcache_tlb_pmp__GEN_39 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_40 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_41 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_2 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_40 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_41 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_42 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_43 =~(~{ dcache_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_2 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_42 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_43 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_2 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_2 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_2 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_2 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_2 =( dcache_tlb_pmp_res_aligned_lsbMask_2 &~( dcache_tlb_pmp_io_pmp_5_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_2 = dcache_tlb_pmp_io_pmp_5_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_2 : dcache_tlb_pmp_res_aligned_rangeAligned_2 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_12 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_13 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_14 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_15 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_16 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_17 ={ dcache_tlb_pmp_io_pmp_5_cfg_x , dcache_tlb_pmp_io_pmp_5_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_2_cfg_r = dcache_tlb_pmp_res_aligned_2 &( dcache_tlb_pmp_io_pmp_5_cfg_r | dcache_tlb_pmp_res_ignore_2 ); 
    wire dcache_tlb_pmp_res_cur_2_cfg_w = dcache_tlb_pmp_res_aligned_2 &( dcache_tlb_pmp_io_pmp_5_cfg_w | dcache_tlb_pmp_res_ignore_2 ); 
    wire dcache_tlb_pmp_res_cur_2_cfg_x = dcache_tlb_pmp_res_aligned_2 &( dcache_tlb_pmp_io_pmp_5_cfg_x | dcache_tlb_pmp_res_ignore_2 ); 
    wire[5:0] dcache_tlb_pmp__GEN_44 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_3 = dcache_tlb_pmp_io_pmp_4_mask |{29'h0,~( dcache_tlb_pmp__GEN_44 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_45 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_3 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_45 [31:3])&~( dcache_tlb_pmp_io_pmp_4_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_46 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_3 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_46 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_3 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_47 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_48 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_6 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_48 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_49 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_6 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_49 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_50 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_6 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_47 [2:0]))< dcache_tlb_pmp__GEN_50 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_51 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_7 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_51 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_52 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_7 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_52 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_53 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_7 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_53 [2:0]; 
    wire dcache_tlb_pmp_res_hit_3 = dcache_tlb_pmp_io_pmp_4_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_3 & dcache_tlb_pmp_res_hit_lsbMatch_3 : dcache_tlb_pmp_io_pmp_4_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_6 | dcache_tlb_pmp_res_hit_msbsEqual_6 & dcache_tlb_pmp_res_hit_lsbsLess_6 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_7 | dcache_tlb_pmp_res_hit_msbsEqual_7 & dcache_tlb_pmp_res_hit_lsbsLess_7 ); 
    wire dcache_tlb_pmp_res_ignore_3 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_4_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_54 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_3 =~( dcache_tlb_pmp__GEN_54 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_55 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_56 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_3 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_55 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_56 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_57 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_58 =~(~{ dcache_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_3 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_57 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_58 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_3 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_3 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_3 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_3 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_3 =( dcache_tlb_pmp_res_aligned_lsbMask_3 &~( dcache_tlb_pmp_io_pmp_4_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_3 = dcache_tlb_pmp_io_pmp_4_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_3 : dcache_tlb_pmp_res_aligned_rangeAligned_3 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_18 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_19 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_20 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_21 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_22 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_23 ={ dcache_tlb_pmp_io_pmp_4_cfg_x , dcache_tlb_pmp_io_pmp_4_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_3_cfg_r = dcache_tlb_pmp_res_aligned_3 &( dcache_tlb_pmp_io_pmp_4_cfg_r | dcache_tlb_pmp_res_ignore_3 ); 
    wire dcache_tlb_pmp_res_cur_3_cfg_w = dcache_tlb_pmp_res_aligned_3 &( dcache_tlb_pmp_io_pmp_4_cfg_w | dcache_tlb_pmp_res_ignore_3 ); 
    wire dcache_tlb_pmp_res_cur_3_cfg_x = dcache_tlb_pmp_res_aligned_3 &( dcache_tlb_pmp_io_pmp_4_cfg_x | dcache_tlb_pmp_res_ignore_3 ); 
    wire[5:0] dcache_tlb_pmp__GEN_59 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_4 = dcache_tlb_pmp_io_pmp_3_mask |{29'h0,~( dcache_tlb_pmp__GEN_59 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_60 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_4 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_60 [31:3])&~( dcache_tlb_pmp_io_pmp_3_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_61 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_4 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_61 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_4 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_62 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_63 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_8 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_63 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_64 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_8 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_64 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_65 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_8 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_62 [2:0]))< dcache_tlb_pmp__GEN_65 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_66 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_9 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_66 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_67 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_9 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_67 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_68 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_9 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_68 [2:0]; 
    wire dcache_tlb_pmp_res_hit_4 = dcache_tlb_pmp_io_pmp_3_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_4 & dcache_tlb_pmp_res_hit_lsbMatch_4 : dcache_tlb_pmp_io_pmp_3_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_8 | dcache_tlb_pmp_res_hit_msbsEqual_8 & dcache_tlb_pmp_res_hit_lsbsLess_8 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_9 | dcache_tlb_pmp_res_hit_msbsEqual_9 & dcache_tlb_pmp_res_hit_lsbsLess_9 ); 
    wire dcache_tlb_pmp_res_ignore_4 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_3_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_69 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_4 =~( dcache_tlb_pmp__GEN_69 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_70 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_71 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_4 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_70 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_71 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_72 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_73 =~(~{ dcache_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_4 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_72 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_73 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_4 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_4 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_4 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_4 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_4 =( dcache_tlb_pmp_res_aligned_lsbMask_4 &~( dcache_tlb_pmp_io_pmp_3_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_4 = dcache_tlb_pmp_io_pmp_3_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_4 : dcache_tlb_pmp_res_aligned_rangeAligned_4 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_24 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_25 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_26 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_27 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_28 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_29 ={ dcache_tlb_pmp_io_pmp_3_cfg_x , dcache_tlb_pmp_io_pmp_3_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_4_cfg_r = dcache_tlb_pmp_res_aligned_4 &( dcache_tlb_pmp_io_pmp_3_cfg_r | dcache_tlb_pmp_res_ignore_4 ); 
    wire dcache_tlb_pmp_res_cur_4_cfg_w = dcache_tlb_pmp_res_aligned_4 &( dcache_tlb_pmp_io_pmp_3_cfg_w | dcache_tlb_pmp_res_ignore_4 ); 
    wire dcache_tlb_pmp_res_cur_4_cfg_x = dcache_tlb_pmp_res_aligned_4 &( dcache_tlb_pmp_io_pmp_3_cfg_x | dcache_tlb_pmp_res_ignore_4 ); 
    wire[5:0] dcache_tlb_pmp__GEN_74 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_5 = dcache_tlb_pmp_io_pmp_2_mask |{29'h0,~( dcache_tlb_pmp__GEN_74 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_75 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_5 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_75 [31:3])&~( dcache_tlb_pmp_io_pmp_2_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_76 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_5 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_76 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_5 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_77 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_78 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_10 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_78 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_79 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_10 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_79 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_80 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_10 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_77 [2:0]))< dcache_tlb_pmp__GEN_80 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_81 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_11 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_81 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_82 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_11 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_82 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_83 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_11 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_83 [2:0]; 
    wire dcache_tlb_pmp_res_hit_5 = dcache_tlb_pmp_io_pmp_2_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_5 & dcache_tlb_pmp_res_hit_lsbMatch_5 : dcache_tlb_pmp_io_pmp_2_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_10 | dcache_tlb_pmp_res_hit_msbsEqual_10 & dcache_tlb_pmp_res_hit_lsbsLess_10 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_11 | dcache_tlb_pmp_res_hit_msbsEqual_11 & dcache_tlb_pmp_res_hit_lsbsLess_11 ); 
    wire dcache_tlb_pmp_res_ignore_5 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_2_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_84 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_5 =~( dcache_tlb_pmp__GEN_84 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_85 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_86 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_5 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_85 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_86 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_87 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_88 =~(~{ dcache_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_5 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_87 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_88 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_5 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_5 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_5 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_5 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_5 =( dcache_tlb_pmp_res_aligned_lsbMask_5 &~( dcache_tlb_pmp_io_pmp_2_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_5 = dcache_tlb_pmp_io_pmp_2_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_5 : dcache_tlb_pmp_res_aligned_rangeAligned_5 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_30 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_31 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_32 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_33 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_34 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_35 ={ dcache_tlb_pmp_io_pmp_2_cfg_x , dcache_tlb_pmp_io_pmp_2_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_5_cfg_r = dcache_tlb_pmp_res_aligned_5 &( dcache_tlb_pmp_io_pmp_2_cfg_r | dcache_tlb_pmp_res_ignore_5 ); 
    wire dcache_tlb_pmp_res_cur_5_cfg_w = dcache_tlb_pmp_res_aligned_5 &( dcache_tlb_pmp_io_pmp_2_cfg_w | dcache_tlb_pmp_res_ignore_5 ); 
    wire dcache_tlb_pmp_res_cur_5_cfg_x = dcache_tlb_pmp_res_aligned_5 &( dcache_tlb_pmp_io_pmp_2_cfg_x | dcache_tlb_pmp_res_ignore_5 ); 
    wire[5:0] dcache_tlb_pmp__GEN_89 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_6 = dcache_tlb_pmp_io_pmp_1_mask |{29'h0,~( dcache_tlb_pmp__GEN_89 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_90 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_6 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_90 [31:3])&~( dcache_tlb_pmp_io_pmp_1_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_91 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_6 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_91 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_6 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_92 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_93 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_12 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_93 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_94 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_12 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_94 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_95 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_12 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_92 [2:0]))< dcache_tlb_pmp__GEN_95 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_96 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_13 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_96 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_97 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_13 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_97 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_98 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_13 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_98 [2:0]; 
    wire dcache_tlb_pmp_res_hit_6 = dcache_tlb_pmp_io_pmp_1_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_6 & dcache_tlb_pmp_res_hit_lsbMatch_6 : dcache_tlb_pmp_io_pmp_1_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_12 | dcache_tlb_pmp_res_hit_msbsEqual_12 & dcache_tlb_pmp_res_hit_lsbsLess_12 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_13 | dcache_tlb_pmp_res_hit_msbsEqual_13 & dcache_tlb_pmp_res_hit_lsbsLess_13 ); 
    wire dcache_tlb_pmp_res_ignore_6 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_1_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_99 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_6 =~( dcache_tlb_pmp__GEN_99 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_100 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_101 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_6 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_100 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_101 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_102 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_103 =~(~{ dcache_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_6 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_102 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_103 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_6 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_6 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_6 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_6 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_6 =( dcache_tlb_pmp_res_aligned_lsbMask_6 &~( dcache_tlb_pmp_io_pmp_1_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_6 = dcache_tlb_pmp_io_pmp_1_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_6 : dcache_tlb_pmp_res_aligned_rangeAligned_6 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_36 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_37 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_38 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_39 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_40 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_41 ={ dcache_tlb_pmp_io_pmp_1_cfg_x , dcache_tlb_pmp_io_pmp_1_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_6_cfg_r = dcache_tlb_pmp_res_aligned_6 &( dcache_tlb_pmp_io_pmp_1_cfg_r | dcache_tlb_pmp_res_ignore_6 ); 
    wire dcache_tlb_pmp_res_cur_6_cfg_w = dcache_tlb_pmp_res_aligned_6 &( dcache_tlb_pmp_io_pmp_1_cfg_w | dcache_tlb_pmp_res_ignore_6 ); 
    wire dcache_tlb_pmp_res_cur_6_cfg_x = dcache_tlb_pmp_res_aligned_6 &( dcache_tlb_pmp_io_pmp_1_cfg_x | dcache_tlb_pmp_res_ignore_6 ); 
    wire[5:0] dcache_tlb_pmp__GEN_104 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp_res_hit_lsbMask_7 = dcache_tlb_pmp_io_pmp_0_mask |{29'h0,~( dcache_tlb_pmp__GEN_104 [2:0])}; 
    wire[31:0] dcache_tlb_pmp__GEN_105 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbMatch_7 =(( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_105 [31:3])&~( dcache_tlb_pmp_io_pmp_0_mask [31:3]))==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_106 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbMatch_7 =(( dcache_tlb_pmp_io_addr [2:0]^ dcache_tlb_pmp__GEN_106 [2:0])&~( dcache_tlb_pmp_res_hit_lsbMask_7 [2:0]))==3'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_107 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[31:0] dcache_tlb_pmp__GEN_108 =~(~{ dcache_tlb_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_14 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_108 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_109 =~(~{ dcache_tlb_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_14 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_109 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_110 =~(~{ dcache_tlb_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_14 =( dcache_tlb_pmp_io_addr [2:0]|~( dcache_tlb_pmp__GEN_107 [2:0]))< dcache_tlb_pmp__GEN_110 [2:0]; 
    wire[31:0] dcache_tlb_pmp__GEN_111 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsLess_15 = dcache_tlb_pmp_io_addr [31:3]< dcache_tlb_pmp__GEN_111 [31:3]; 
    wire[31:0] dcache_tlb_pmp__GEN_112 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_msbsEqual_15 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_112 [31:3])==29'h0; 
    wire[31:0] dcache_tlb_pmp__GEN_113 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_hit_lsbsLess_15 = dcache_tlb_pmp_io_addr [2:0]< dcache_tlb_pmp__GEN_113 [2:0]; 
    wire dcache_tlb_pmp_res_hit_7 = dcache_tlb_pmp_io_pmp_0_cfg_a [1] ?  dcache_tlb_pmp_res_hit_msbMatch_7 & dcache_tlb_pmp_res_hit_lsbMatch_7 : dcache_tlb_pmp_io_pmp_0_cfg_a [0]&( dcache_tlb_pmp_res_hit_msbsLess_14 | dcache_tlb_pmp_res_hit_msbsEqual_14 & dcache_tlb_pmp_res_hit_lsbsLess_14 )==1'h0&( dcache_tlb_pmp_res_hit_msbsLess_15 | dcache_tlb_pmp_res_hit_msbsEqual_15 & dcache_tlb_pmp_res_hit_lsbsLess_15 ); 
    wire dcache_tlb_pmp_res_ignore_7 = dcache_tlb_pmp_default_0 & dcache_tlb_pmp_io_pmp_0_cfg_l ==1'h0; 
    wire[5:0] dcache_tlb_pmp__GEN_114 =6'h7<< dcache_tlb_pmp_io_size ; 
    wire[2:0] dcache_tlb_pmp_res_aligned_lsbMask_7 =~( dcache_tlb_pmp__GEN_114 [2:0]); 
    wire[31:0] dcache_tlb_pmp__GEN_115 =~(~{ dcache_tlb_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_116 =~(~{ dcache_tlb_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesLowerBound_7 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_115 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_116 [2:0]&~( dcache_tlb_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_tlb_pmp__GEN_117 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_tlb_pmp__GEN_118 =~(~{ dcache_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_tlb_pmp_res_aligned_straddlesUpperBound_7 =( dcache_tlb_pmp_io_addr [31:3]^ dcache_tlb_pmp__GEN_117 [31:3])==29'h0&(|( dcache_tlb_pmp__GEN_118 [2:0]&( dcache_tlb_pmp_io_addr [2:0]| dcache_tlb_pmp_res_aligned_lsbMask_7 ))); 
    wire dcache_tlb_pmp_res_aligned_rangeAligned_7 =( dcache_tlb_pmp_res_aligned_straddlesLowerBound_7 | dcache_tlb_pmp_res_aligned_straddlesUpperBound_7 )==1'h0; 
    wire dcache_tlb_pmp_res_aligned_pow2Aligned_7 =( dcache_tlb_pmp_res_aligned_lsbMask_7 &~( dcache_tlb_pmp_io_pmp_0_mask [2:0]))==3'h0; 
    wire dcache_tlb_pmp_res_aligned_7 = dcache_tlb_pmp_io_pmp_0_cfg_a [1] ?  dcache_tlb_pmp_res_aligned_pow2Aligned_7 : dcache_tlb_pmp_res_aligned_rangeAligned_7 ; 
    wire[1:0] dcache_tlb_pmp_res_hi_42 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_43 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_44 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_45 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_46 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_tlb_pmp_res_hi_47 ={ dcache_tlb_pmp_io_pmp_0_cfg_x , dcache_tlb_pmp_io_pmp_0_cfg_w }; 
    wire dcache_tlb_pmp_res_cur_7_cfg_r = dcache_tlb_pmp_res_aligned_7 &( dcache_tlb_pmp_io_pmp_0_cfg_r | dcache_tlb_pmp_res_ignore_7 ); 
    wire dcache_tlb_pmp_res_cur_7_cfg_w = dcache_tlb_pmp_res_aligned_7 &( dcache_tlb_pmp_io_pmp_0_cfg_w | dcache_tlb_pmp_res_ignore_7 ); 
    wire dcache_tlb_pmp_res_cur_7_cfg_x = dcache_tlb_pmp_res_aligned_7 &( dcache_tlb_pmp_io_pmp_0_cfg_x | dcache_tlb_pmp_res_ignore_7 ); 
    wire dcache_tlb_pmp_res_cfg_l = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_l : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_l : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_l : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_l : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_l : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_l : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_l : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_l : dcache_tlb_pmp_pmp0_cfg_l ; 
    wire[1:0] dcache_tlb_pmp_res_cfg_res = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_res : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_res : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_res : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_res : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_res : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_res : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_res : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_res : dcache_tlb_pmp_pmp0_cfg_res ; 
    wire[1:0] dcache_tlb_pmp_res_cfg_a = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_a : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_a : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_a : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_a : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_a : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_a : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_a : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_a : dcache_tlb_pmp_pmp0_cfg_a ; 
    wire dcache_tlb_pmp_res_cfg_x = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_x : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_x : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_x : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_x : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_x : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_x : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_x : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_x : dcache_tlb_pmp_pmp0_cfg_x ; 
    wire dcache_tlb_pmp_res_cfg_w = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_w : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_w : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_w : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_w : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_w : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_w : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_w : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_w : dcache_tlb_pmp_pmp0_cfg_w ; 
    wire dcache_tlb_pmp_res_cfg_r = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_cfg_r : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_cfg_r : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_cfg_r : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_cfg_r : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_cfg_r : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_cfg_r : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_cfg_r : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_cfg_r : dcache_tlb_pmp_pmp0_cfg_r ; 
    wire[29:0] dcache_tlb_pmp_res_addr = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_addr : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_addr : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_addr : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_addr : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_addr : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_addr : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_addr : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_addr : dcache_tlb_pmp_pmp0_addr ; 
    wire[31:0] dcache_tlb_pmp_res_mask = dcache_tlb_pmp_res_hit_7  ?  dcache_tlb_pmp_res_cur_7_mask : dcache_tlb_pmp_res_hit_6  ?  dcache_tlb_pmp_res_cur_6_mask : dcache_tlb_pmp_res_hit_5  ?  dcache_tlb_pmp_res_cur_5_mask : dcache_tlb_pmp_res_hit_4  ?  dcache_tlb_pmp_res_cur_4_mask : dcache_tlb_pmp_res_hit_3  ?  dcache_tlb_pmp_res_cur_3_mask : dcache_tlb_pmp_res_hit_2  ?  dcache_tlb_pmp_res_cur_2_mask : dcache_tlb_pmp_res_hit_1  ?  dcache_tlb_pmp_res_cur_1_mask : dcache_tlb_pmp_res_hit  ?  dcache_tlb_pmp_res_cur_mask : dcache_tlb_pmp_pmp0_mask ; 
  assign  dcache_tlb_pmp_io_r = dcache_tlb_pmp_res_cfg_r ; 
  assign  dcache_tlb_pmp_io_w = dcache_tlb_pmp_res_cfg_w ; 
  assign  dcache_tlb_pmp_io_x = dcache_tlb_pmp_res_cfg_x ;
     
  assign  dcache__tlb_mpu_physaddr_31to0 = dcache_tlb_mpu_physaddr [31:0]; 
  assign  dcache__tlb_mpu_priv_1to0 = dcache_tlb_mpu_priv [1:0]; 
    wire dcache_tlb__legal_address_WIRE_0 =({1'h0, dcache_tlb_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_1 =({1'h0, dcache_tlb_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_2 =({1'h0, dcache_tlb_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_3 =({1'h0, dcache_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_4 =({1'h0, dcache_tlb_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_5 =({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire dcache_tlb__legal_address_WIRE_6 =({1'h0, dcache_tlb_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0; 
    wire dcache_tlb_legal_address = dcache_tlb__legal_address_WIRE_0 | dcache_tlb__legal_address_WIRE_1 | dcache_tlb__legal_address_WIRE_2 | dcache_tlb__legal_address_WIRE_3 | dcache_tlb__legal_address_WIRE_4 | dcache_tlb__legal_address_WIRE_5 | dcache_tlb__legal_address_WIRE_6 ; 
    wire dcache_tlb__cacheable_WIRE =({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'h80000000)==35'h0|1'h0; 
    wire dcache_tlb_cacheable = dcache_tlb_legal_address & dcache_tlb__cacheable_WIRE ; 
    wire dcache_tlb_newEntry_c = dcache_tlb_cacheable ; 
    wire dcache_tlb_homogeneous =({1'h0, dcache_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0|1'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire dcache_tlb_deny_access_to_debug = dcache_tlb_mpu_priv <=3'h3&({1'h0, dcache_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire dcache_tlb_prot_r = dcache_tlb_legal_address & dcache_tlb_deny_access_to_debug ==1'h0& dcache__tlb_pmp_io_r ; 
    wire dcache_tlb_newEntry_pr = dcache_tlb_prot_r ; 
    wire dcache_tlb__prot_w_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_tlb_prot_w = dcache_tlb_legal_address & dcache_tlb__prot_w_WIRE & dcache_tlb_deny_access_to_debug ==1'h0& dcache__tlb_pmp_io_w ; 
    wire dcache_tlb_newEntry_pw = dcache_tlb_prot_w ; 
    wire dcache_tlb__prot_pp_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_tlb_prot_pp = dcache_tlb_legal_address & dcache_tlb__prot_pp_WIRE ; 
    wire dcache_tlb_newEntry_ppp = dcache_tlb_prot_pp ; 
    wire dcache_tlb__prot_al_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire dcache_tlb_prot_al = dcache_tlb_legal_address & dcache_tlb__prot_al_WIRE ; 
    wire dcache_tlb_newEntry_pal = dcache_tlb_prot_al ; 
    wire dcache_tlb__prot_aa_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire dcache_tlb_prot_aa = dcache_tlb_legal_address & dcache_tlb__prot_aa_WIRE ; 
    wire dcache_tlb_newEntry_paa = dcache_tlb_prot_aa ; 
    wire dcache_tlb__prot_x_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hCA000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_tlb_prot_x = dcache_tlb_legal_address & dcache_tlb__prot_x_WIRE & dcache_tlb_deny_access_to_debug ==1'h0& dcache__tlb_pmp_io_x ; 
    wire dcache_tlb_newEntry_px = dcache_tlb_prot_x ; 
    wire dcache_tlb__prot_eff_WIRE =({1'h0, dcache_tlb_mpu_physaddr }&35'hCA012000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|1'h0; 
    wire dcache_tlb_prot_eff = dcache_tlb_legal_address & dcache_tlb__prot_eff_WIRE ; 
    wire dcache_tlb_newEntry_eff = dcache_tlb_prot_eff ; 
    wire[20:0] dcache__GEN_0 = dcache_tlb_sectored_entries_0_0_tag_vpn ^ dcache_tlb_vpn ; 
    wire dcache_tlb_sector_hits_0 =( dcache_tlb_sectored_entries_0_0_valid_0 | dcache_tlb_sectored_entries_0_0_valid_1 | dcache_tlb_sectored_entries_0_0_valid_2 | dcache_tlb_sectored_entries_0_0_valid_3 )& dcache__GEN_0 [20:2]==19'h0& dcache_tlb_sectored_entries_0_0_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_superpage_hits_0 = dcache_tlb_superpage_entries_0_valid_0 &( dcache_tlb_superpage_entries_0_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_0_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_superpage_hits_1 = dcache_tlb_superpage_entries_1_valid_0 &( dcache_tlb_superpage_entries_1_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_1_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_superpage_hits_2 = dcache_tlb_superpage_entries_2_valid_0 &( dcache_tlb_superpage_entries_2_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_2_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_superpage_hits_3 = dcache_tlb_superpage_entries_3_valid_0 &( dcache_tlb_superpage_entries_3_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_3_tag_v == dcache_tlb_priv_v ; 
    wire[1:0] dcache_tlb_hitsVec_idx = dcache_tlb_vpn [1:0]; 
    wire[20:0] dcache__GEN_1 = dcache_tlb_sectored_entries_0_0_tag_vpn ^ dcache_tlb_vpn ; 
    reg dcache_casez_tmp ; 
  always @(*)
         begin 
             casez ( dcache_tlb_hitsVec_idx )
              2 'b00: 
                  dcache_casez_tmp  = dcache_tlb_sectored_entries_0_0_valid_0 ;
              2 'b01: 
                  dcache_casez_tmp  = dcache_tlb_sectored_entries_0_0_valid_1 ;
              2 'b10: 
                  dcache_casez_tmp  = dcache_tlb_sectored_entries_0_0_valid_2 ;
              default : 
                  dcache_casez_tmp  = dcache_tlb_sectored_entries_0_0_valid_3 ;endcase
         end
    wire dcache_tlb_hitsVec_0 = dcache_tlb_vm_enabled & dcache_casez_tmp & dcache__GEN_1 [20:2]==19'h0& dcache_tlb_sectored_entries_0_0_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_hitsVec_1 = dcache_tlb_vm_enabled & dcache_tlb_superpage_entries_0_valid_0 &( dcache_tlb_superpage_entries_0_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_0_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_hitsVec_2 = dcache_tlb_vm_enabled & dcache_tlb_superpage_entries_1_valid_0 &( dcache_tlb_superpage_entries_1_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_1_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_hitsVec_3 = dcache_tlb_vm_enabled & dcache_tlb_superpage_entries_2_valid_0 &( dcache_tlb_superpage_entries_2_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_2_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_hitsVec_4 = dcache_tlb_vm_enabled & dcache_tlb_superpage_entries_3_valid_0 &( dcache_tlb_superpage_entries_3_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_superpage_entries_3_tag_v == dcache_tlb_priv_v ; 
    wire dcache_tlb_hitsVec_5 = dcache_tlb_vm_enabled & dcache_tlb_special_entry_valid_0 &( dcache_tlb_special_entry_tag_vpn ^ dcache_tlb_vpn )==21'h0& dcache_tlb_special_entry_tag_v == dcache_tlb_priv_v ; 
    wire[1:0] dcache_tlb_real_hits_lo_hi ={ dcache_tlb_hitsVec_2 , dcache_tlb_hitsVec_1 }; 
    wire[2:0] dcache_tlb_real_hits_lo ={ dcache_tlb_real_hits_lo_hi , dcache_tlb_hitsVec_0 }; 
    wire[1:0] dcache_tlb_real_hits_hi_hi ={ dcache_tlb_hitsVec_5 , dcache_tlb_hitsVec_4 }; 
    wire[2:0] dcache_tlb_real_hits_hi ={ dcache_tlb_real_hits_hi_hi , dcache_tlb_hitsVec_3 }; 
    wire[5:0] dcache_tlb_real_hits ={ dcache_tlb_real_hits_hi , dcache_tlb_real_hits_lo }; 
    wire[6:0] dcache_tlb_hits ={ dcache_tlb_vm_enabled ==1'h0, dcache_tlb_real_hits }; 
    wire dcache_tlb_refill_v = dcache_tlb_r_vstage1_en | dcache_tlb_r_stage2_en ; 
    wire[19:0] dcache_tlb_newEntry_ppn = dcache_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire dcache_tlb_newEntry_g = dcache_tlb_io_ptw_resp_bits_pte_g & dcache_tlb_io_ptw_resp_bits_pte_v ; 
    wire dcache_tlb_newEntry_ae_stage2 = dcache_tlb_io_ptw_resp_bits_ae_final & dcache_tlb_io_ptw_resp_bits_gpa_is_pte & dcache_tlb_r_stage2_en ; 
    wire dcache_tlb_newEntry_sr = dcache_tlb_io_ptw_resp_bits_pte_v &( dcache_tlb_io_ptw_resp_bits_pte_r | dcache_tlb_io_ptw_resp_bits_pte_x & dcache_tlb_io_ptw_resp_bits_pte_w ==1'h0)& dcache_tlb_io_ptw_resp_bits_pte_a & dcache_tlb_io_ptw_resp_bits_pte_r ; 
    wire dcache_tlb_newEntry_sw = dcache_tlb_io_ptw_resp_bits_pte_v &( dcache_tlb_io_ptw_resp_bits_pte_r | dcache_tlb_io_ptw_resp_bits_pte_x & dcache_tlb_io_ptw_resp_bits_pte_w ==1'h0)& dcache_tlb_io_ptw_resp_bits_pte_a & dcache_tlb_io_ptw_resp_bits_pte_w & dcache_tlb_io_ptw_resp_bits_pte_d ; 
    wire dcache_tlb_newEntry_sx = dcache_tlb_io_ptw_resp_bits_pte_v &( dcache_tlb_io_ptw_resp_bits_pte_r | dcache_tlb_io_ptw_resp_bits_pte_x & dcache_tlb_io_ptw_resp_bits_pte_w ==1'h0)& dcache_tlb_io_ptw_resp_bits_pte_a & dcache_tlb_io_ptw_resp_bits_pte_x ; 
    wire dcache__GEN_2 = dcache_tlb_io_ptw_resp_bits_homogeneous ==1'h0&1'h1; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_lo_hi ={ dcache_tlb_special_entry_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_special_entry_data_0_lo_lo ={ dcache_tlb_special_entry_data_0_lo_lo_hi , dcache_tlb_special_entry_data_0_lo_lo_lo }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_hi_lo ={ dcache_tlb_special_entry_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_special_entry_data_0_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_special_entry_data_0_lo_hi_hi ={ dcache_tlb_special_entry_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_special_entry_data_0_lo_hi ={ dcache_tlb_special_entry_data_0_lo_hi_hi , dcache_tlb_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_special_entry_data_0_lo ={ dcache_tlb_special_entry_data_0_lo_hi , dcache_tlb_special_entry_data_0_lo_lo }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_lo_lo ={ dcache_tlb_special_entry_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_lo_hi ={ dcache_tlb_special_entry_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_special_entry_data_0_hi_lo ={ dcache_tlb_special_entry_data_0_hi_lo_hi , dcache_tlb_special_entry_data_0_hi_lo_lo }; 
    wire[1:0] dcache_tlb_special_entry_data_0_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_special_entry_data_0_hi_hi_lo ={ dcache_tlb_special_entry_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_special_entry_data_0_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_special_entry_data_0_hi_hi_hi ={ dcache_tlb_special_entry_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_special_entry_data_0_hi_hi ={ dcache_tlb_special_entry_data_0_hi_hi_hi , dcache_tlb_special_entry_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_special_entry_data_0_hi ={ dcache_tlb_special_entry_data_0_hi_hi , dcache_tlb_special_entry_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_3 ={ dcache_tlb_special_entry_data_0_hi , dcache_tlb_special_entry_data_0_lo }; 
    wire dcache__GEN_4 = dcache_tlb_do_refill &~ dcache__GEN_2 ; 
    wire dcache__GEN_5 = dcache_tlb_io_ptw_resp_bits_level <2'h2; 
    wire dcache__GEN_6 = dcache__GEN_4 & dcache__GEN_5 ; 
    wire dcache__GEN_7 = dcache_tlb_r_superpage_repl_addr ==2'h0; 
    wire[1:0] dcache__GEN_8 ={1'h0, dcache_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_0_data_0_lo_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_lo_hi , dcache_tlb_superpage_entries_0_data_0_lo_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_0_data_0_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_lo_hi_hi , dcache_tlb_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_0_data_0_lo ={ dcache_tlb_superpage_entries_0_data_0_lo_hi , dcache_tlb_superpage_entries_0_data_0_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_0_data_0_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_lo_hi , dcache_tlb_superpage_entries_0_data_0_hi_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_superpage_entries_0_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_0_data_0_hi_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi_hi , dcache_tlb_superpage_entries_0_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_0_data_0_hi ={ dcache_tlb_superpage_entries_0_data_0_hi_hi , dcache_tlb_superpage_entries_0_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_9 ={ dcache_tlb_superpage_entries_0_data_0_hi , dcache_tlb_superpage_entries_0_data_0_lo }; 
    wire dcache__GEN_10 = dcache_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_11 = dcache_tlb_r_superpage_repl_addr ==2'h1; 
    wire[1:0] dcache__GEN_12 ={1'h0, dcache_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_1_data_0_lo_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_lo_hi , dcache_tlb_superpage_entries_1_data_0_lo_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_1_data_0_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_lo_hi_hi , dcache_tlb_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_1_data_0_lo ={ dcache_tlb_superpage_entries_1_data_0_lo_hi , dcache_tlb_superpage_entries_1_data_0_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_1_data_0_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_lo_hi , dcache_tlb_superpage_entries_1_data_0_hi_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_superpage_entries_1_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_1_data_0_hi_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi_hi , dcache_tlb_superpage_entries_1_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_1_data_0_hi ={ dcache_tlb_superpage_entries_1_data_0_hi_hi , dcache_tlb_superpage_entries_1_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_13 ={ dcache_tlb_superpage_entries_1_data_0_hi , dcache_tlb_superpage_entries_1_data_0_lo }; 
    wire dcache__GEN_14 = dcache_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_15 = dcache_tlb_r_superpage_repl_addr ==2'h2; 
    wire[1:0] dcache__GEN_16 ={1'h0, dcache_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_2_data_0_lo_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_lo_hi , dcache_tlb_superpage_entries_2_data_0_lo_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_2_data_0_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_lo_hi_hi , dcache_tlb_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_2_data_0_lo ={ dcache_tlb_superpage_entries_2_data_0_lo_hi , dcache_tlb_superpage_entries_2_data_0_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_2_data_0_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_lo_hi , dcache_tlb_superpage_entries_2_data_0_hi_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_superpage_entries_2_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_2_data_0_hi_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi_hi , dcache_tlb_superpage_entries_2_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_2_data_0_hi ={ dcache_tlb_superpage_entries_2_data_0_hi_hi , dcache_tlb_superpage_entries_2_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_17 ={ dcache_tlb_superpage_entries_2_data_0_hi , dcache_tlb_superpage_entries_2_data_0_lo }; 
    wire dcache__GEN_18 = dcache_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_19 =& dcache_tlb_r_superpage_repl_addr ; 
    wire[1:0] dcache__GEN_20 ={1'h0, dcache_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_superpage_entries_3_data_0_lo_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_lo_hi , dcache_tlb_superpage_entries_3_data_0_lo_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_lo_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_superpage_entries_3_data_0_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_lo_hi_hi , dcache_tlb_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] dcache_tlb_superpage_entries_3_data_0_lo ={ dcache_tlb_superpage_entries_3_data_0_lo_hi , dcache_tlb_superpage_entries_3_data_0_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_lo_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_superpage_entries_3_data_0_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_lo_hi , dcache_tlb_superpage_entries_3_data_0_hi_lo_lo }; 
    wire[1:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_lo ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_superpage_entries_3_data_0_hi_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_superpage_entries_3_data_0_hi_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi_hi , dcache_tlb_superpage_entries_3_data_0_hi_hi_lo }; 
    wire[30:0] dcache_tlb_superpage_entries_3_data_0_hi ={ dcache_tlb_superpage_entries_3_data_0_hi_hi , dcache_tlb_superpage_entries_3_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_21 ={ dcache_tlb_superpage_entries_3_data_0_hi , dcache_tlb_superpage_entries_3_data_0_lo }; 
    wire dcache__GEN_22 = dcache_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_23 = dcache__GEN_4 &~ dcache__GEN_5 ; 
    wire dcache__GEN_24 = dcache_tlb_r_sectored_hit_valid ==1'h0; 
    wire[1:0] dcache_tlb_idx = dcache_tlb_r_refill_tag [1:0]; 
    wire dcache__GEN_25 = dcache_tlb_idx ==2'h0; 
    wire dcache__GEN_26 = dcache_tlb_idx ==2'h1; 
    wire dcache__GEN_27 = dcache_tlb_idx ==2'h2; 
    wire dcache__GEN_28 =& dcache_tlb_idx ; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_lo ={ dcache_tlb_newEntry_c , dcache_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_hi_hi ={ dcache_tlb_newEntry_pal , dcache_tlb_newEntry_paa }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_lo_hi_hi , dcache_tlb_newEntry_eff }; 
    wire[4:0] dcache_tlb_sectored_entries_0_0_data_lo_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_lo_hi , dcache_tlb_sectored_entries_0_0_data_lo_lo_lo }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_lo_hi ={ dcache_tlb_newEntry_px , dcache_tlb_newEntry_pr }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_lo_hi , dcache_tlb_newEntry_ppp }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_hi_hi ={ dcache_tlb_newEntry_hx , dcache_tlb_newEntry_hr }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_lo_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_hi_hi , dcache_tlb_newEntry_pw }; 
    wire[5:0] dcache_tlb_sectored_entries_0_0_data_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_lo_hi_hi , dcache_tlb_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] dcache_tlb_sectored_entries_0_0_data_lo ={ dcache_tlb_sectored_entries_0_0_data_lo_hi , dcache_tlb_sectored_entries_0_0_data_lo_lo }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_lo_hi ={ dcache_tlb_newEntry_sx , dcache_tlb_newEntry_sr }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_lo_hi , dcache_tlb_newEntry_hw }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_hi_hi ={ dcache_tlb_newEntry_pf , dcache_tlb_newEntry_gf }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_lo_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_hi_hi , dcache_tlb_newEntry_sw }; 
    wire[5:0] dcache_tlb_sectored_entries_0_0_data_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_lo_hi , dcache_tlb_sectored_entries_0_0_data_hi_lo_lo }; 
    wire[1:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_lo_hi ={ dcache_tlb_newEntry_ae_ptw , dcache_tlb_newEntry_ae_final }; 
    wire[2:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_lo ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_lo_hi , dcache_tlb_newEntry_ae_stage2 }; 
    wire[20:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_hi_hi ={ dcache_tlb_newEntry_ppn , dcache_tlb_newEntry_u }; 
    wire[21:0] dcache_tlb_sectored_entries_0_0_data_hi_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_hi_hi , dcache_tlb_newEntry_g }; 
    wire[24:0] dcache_tlb_sectored_entries_0_0_data_hi_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi_hi , dcache_tlb_sectored_entries_0_0_data_hi_hi_lo }; 
    wire[30:0] dcache_tlb_sectored_entries_0_0_data_hi ={ dcache_tlb_sectored_entries_0_0_data_hi_hi , dcache_tlb_sectored_entries_0_0_data_hi_lo }; 
    wire[41:0] dcache__GEN_29 ={ dcache_tlb_sectored_entries_0_0_data_hi , dcache_tlb_sectored_entries_0_0_data_lo }; 
    wire dcache__GEN_30 = dcache_tlb_idx ==2'h0; 
    wire dcache__GEN_31 = dcache_tlb_idx ==2'h1; 
    wire dcache__GEN_32 = dcache_tlb_idx ==2'h2; 
    wire dcache__GEN_33 =& dcache_tlb_idx ; reg[41:0] dcache_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( dcache_tlb_vpn [1:0])
              2 'b00: 
                  dcache_casez_tmp_0  = dcache_tlb_sectored_entries_0_0_data_0 ;
              2 'b01: 
                  dcache_casez_tmp_0  = dcache_tlb_sectored_entries_0_0_data_1 ;
              2 'b10: 
                  dcache_casez_tmp_0  = dcache_tlb_sectored_entries_0_0_data_2 ;
              default : 
                  dcache_casez_tmp_0  = dcache_tlb_sectored_entries_0_0_data_3 ;endcase
         end
    wire[41:0] dcache_tlb__entries_WIRE_1 = dcache_casez_tmp_0 ; 
    wire dcache_tlb__entries_WIRE_fragmented_superpage = dcache_tlb__entries_WIRE_1 [0]; 
    wire dcache_tlb__entries_WIRE_c = dcache_tlb__entries_WIRE_1 [1]; 
    wire dcache_tlb__entries_WIRE_eff = dcache_tlb__entries_WIRE_1 [2]; 
    wire dcache_tlb__entries_WIRE_paa = dcache_tlb__entries_WIRE_1 [3]; 
    wire dcache_tlb__entries_WIRE_pal = dcache_tlb__entries_WIRE_1 [4]; 
    wire dcache_tlb__entries_WIRE_ppp = dcache_tlb__entries_WIRE_1 [5]; 
    wire dcache_tlb__entries_WIRE_pr = dcache_tlb__entries_WIRE_1 [6]; 
    wire dcache_tlb__entries_WIRE_px = dcache_tlb__entries_WIRE_1 [7]; 
    wire dcache_tlb__entries_WIRE_pw = dcache_tlb__entries_WIRE_1 [8]; 
    wire dcache_tlb__entries_WIRE_hr = dcache_tlb__entries_WIRE_1 [9]; 
    wire dcache_tlb__entries_WIRE_hx = dcache_tlb__entries_WIRE_1 [10]; 
    wire dcache_tlb__entries_WIRE_hw = dcache_tlb__entries_WIRE_1 [11]; 
    wire dcache_tlb__entries_WIRE_sr = dcache_tlb__entries_WIRE_1 [12]; 
    wire dcache_tlb__entries_WIRE_sx = dcache_tlb__entries_WIRE_1 [13]; 
    wire dcache_tlb__entries_WIRE_sw = dcache_tlb__entries_WIRE_1 [14]; 
    wire dcache_tlb__entries_WIRE_gf = dcache_tlb__entries_WIRE_1 [15]; 
    wire dcache_tlb__entries_WIRE_pf = dcache_tlb__entries_WIRE_1 [16]; 
    wire dcache_tlb__entries_WIRE_ae_stage2 = dcache_tlb__entries_WIRE_1 [17]; 
    wire dcache_tlb__entries_WIRE_ae_final = dcache_tlb__entries_WIRE_1 [18]; 
    wire dcache_tlb__entries_WIRE_ae_ptw = dcache_tlb__entries_WIRE_1 [19]; 
    wire dcache_tlb__entries_WIRE_g = dcache_tlb__entries_WIRE_1 [20]; 
    wire dcache_tlb__entries_WIRE_u = dcache_tlb__entries_WIRE_1 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_ppn = dcache_tlb__entries_WIRE_1 [41:22];  
    
    assign  dcache_tlb_entries_barrier_io_y_ppn = dcache_tlb_entries_barrier_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_io_y_u = dcache_tlb_entries_barrier_io_x_u ; 
  assign  dcache_tlb_entries_barrier_io_y_g = dcache_tlb_entries_barrier_io_x_g ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_ptw = dcache_tlb_entries_barrier_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_final = dcache_tlb_entries_barrier_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_io_y_ae_stage2 = dcache_tlb_entries_barrier_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_io_y_pf = dcache_tlb_entries_barrier_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_io_y_gf = dcache_tlb_entries_barrier_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_io_y_sw = dcache_tlb_entries_barrier_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_io_y_sx = dcache_tlb_entries_barrier_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_io_y_sr = dcache_tlb_entries_barrier_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_io_y_hw = dcache_tlb_entries_barrier_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_io_y_hx = dcache_tlb_entries_barrier_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_io_y_hr = dcache_tlb_entries_barrier_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_io_y_pw = dcache_tlb_entries_barrier_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_io_y_px = dcache_tlb_entries_barrier_io_x_px ; 
  assign  dcache_tlb_entries_barrier_io_y_pr = dcache_tlb_entries_barrier_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_io_y_ppp = dcache_tlb_entries_barrier_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_io_y_pal = dcache_tlb_entries_barrier_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_io_y_paa = dcache_tlb_entries_barrier_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_io_y_eff = dcache_tlb_entries_barrier_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_io_y_c = dcache_tlb_entries_barrier_io_x_c ; 
  assign  dcache_tlb_entries_barrier_io_y_fragmented_superpage = dcache_tlb_entries_barrier_io_x_fragmented_superpage ;
     
    wire dcache_tlb__entries_WIRE_2_fragmented_superpage = dcache_tlb__entries_WIRE_3 [0]; 
    wire dcache_tlb__entries_WIRE_2_c = dcache_tlb__entries_WIRE_3 [1]; 
    wire dcache_tlb__entries_WIRE_2_eff = dcache_tlb__entries_WIRE_3 [2]; 
    wire dcache_tlb__entries_WIRE_2_paa = dcache_tlb__entries_WIRE_3 [3]; 
    wire dcache_tlb__entries_WIRE_2_pal = dcache_tlb__entries_WIRE_3 [4]; 
    wire dcache_tlb__entries_WIRE_2_ppp = dcache_tlb__entries_WIRE_3 [5]; 
    wire dcache_tlb__entries_WIRE_2_pr = dcache_tlb__entries_WIRE_3 [6]; 
    wire dcache_tlb__entries_WIRE_2_px = dcache_tlb__entries_WIRE_3 [7]; 
    wire dcache_tlb__entries_WIRE_2_pw = dcache_tlb__entries_WIRE_3 [8]; 
    wire dcache_tlb__entries_WIRE_2_hr = dcache_tlb__entries_WIRE_3 [9]; 
    wire dcache_tlb__entries_WIRE_2_hx = dcache_tlb__entries_WIRE_3 [10]; 
    wire dcache_tlb__entries_WIRE_2_hw = dcache_tlb__entries_WIRE_3 [11]; 
    wire dcache_tlb__entries_WIRE_2_sr = dcache_tlb__entries_WIRE_3 [12]; 
    wire dcache_tlb__entries_WIRE_2_sx = dcache_tlb__entries_WIRE_3 [13]; 
    wire dcache_tlb__entries_WIRE_2_sw = dcache_tlb__entries_WIRE_3 [14]; 
    wire dcache_tlb__entries_WIRE_2_gf = dcache_tlb__entries_WIRE_3 [15]; 
    wire dcache_tlb__entries_WIRE_2_pf = dcache_tlb__entries_WIRE_3 [16]; 
    wire dcache_tlb__entries_WIRE_2_ae_stage2 = dcache_tlb__entries_WIRE_3 [17]; 
    wire dcache_tlb__entries_WIRE_2_ae_final = dcache_tlb__entries_WIRE_3 [18]; 
    wire dcache_tlb__entries_WIRE_2_ae_ptw = dcache_tlb__entries_WIRE_3 [19]; 
    wire dcache_tlb__entries_WIRE_2_g = dcache_tlb__entries_WIRE_3 [20]; 
    wire dcache_tlb__entries_WIRE_2_u = dcache_tlb__entries_WIRE_3 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_2_ppn = dcache_tlb__entries_WIRE_3 [41:22];  
    
    assign  dcache_tlb_entries_barrier_1_io_y_ppn = dcache_tlb_entries_barrier_1_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_1_io_y_u = dcache_tlb_entries_barrier_1_io_x_u ; 
  assign  dcache_tlb_entries_barrier_1_io_y_g = dcache_tlb_entries_barrier_1_io_x_g ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_ptw = dcache_tlb_entries_barrier_1_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_final = dcache_tlb_entries_barrier_1_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ae_stage2 = dcache_tlb_entries_barrier_1_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pf = dcache_tlb_entries_barrier_1_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_1_io_y_gf = dcache_tlb_entries_barrier_1_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sw = dcache_tlb_entries_barrier_1_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sx = dcache_tlb_entries_barrier_1_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_1_io_y_sr = dcache_tlb_entries_barrier_1_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hw = dcache_tlb_entries_barrier_1_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hx = dcache_tlb_entries_barrier_1_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_1_io_y_hr = dcache_tlb_entries_barrier_1_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pw = dcache_tlb_entries_barrier_1_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_1_io_y_px = dcache_tlb_entries_barrier_1_io_x_px ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pr = dcache_tlb_entries_barrier_1_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_1_io_y_ppp = dcache_tlb_entries_barrier_1_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_1_io_y_pal = dcache_tlb_entries_barrier_1_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_1_io_y_paa = dcache_tlb_entries_barrier_1_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_1_io_y_eff = dcache_tlb_entries_barrier_1_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_1_io_y_c = dcache_tlb_entries_barrier_1_io_x_c ; 
  assign  dcache_tlb_entries_barrier_1_io_y_fragmented_superpage = dcache_tlb_entries_barrier_1_io_x_fragmented_superpage ;
     
    wire dcache_tlb__entries_WIRE_4_fragmented_superpage = dcache_tlb__entries_WIRE_5 [0]; 
    wire dcache_tlb__entries_WIRE_4_c = dcache_tlb__entries_WIRE_5 [1]; 
    wire dcache_tlb__entries_WIRE_4_eff = dcache_tlb__entries_WIRE_5 [2]; 
    wire dcache_tlb__entries_WIRE_4_paa = dcache_tlb__entries_WIRE_5 [3]; 
    wire dcache_tlb__entries_WIRE_4_pal = dcache_tlb__entries_WIRE_5 [4]; 
    wire dcache_tlb__entries_WIRE_4_ppp = dcache_tlb__entries_WIRE_5 [5]; 
    wire dcache_tlb__entries_WIRE_4_pr = dcache_tlb__entries_WIRE_5 [6]; 
    wire dcache_tlb__entries_WIRE_4_px = dcache_tlb__entries_WIRE_5 [7]; 
    wire dcache_tlb__entries_WIRE_4_pw = dcache_tlb__entries_WIRE_5 [8]; 
    wire dcache_tlb__entries_WIRE_4_hr = dcache_tlb__entries_WIRE_5 [9]; 
    wire dcache_tlb__entries_WIRE_4_hx = dcache_tlb__entries_WIRE_5 [10]; 
    wire dcache_tlb__entries_WIRE_4_hw = dcache_tlb__entries_WIRE_5 [11]; 
    wire dcache_tlb__entries_WIRE_4_sr = dcache_tlb__entries_WIRE_5 [12]; 
    wire dcache_tlb__entries_WIRE_4_sx = dcache_tlb__entries_WIRE_5 [13]; 
    wire dcache_tlb__entries_WIRE_4_sw = dcache_tlb__entries_WIRE_5 [14]; 
    wire dcache_tlb__entries_WIRE_4_gf = dcache_tlb__entries_WIRE_5 [15]; 
    wire dcache_tlb__entries_WIRE_4_pf = dcache_tlb__entries_WIRE_5 [16]; 
    wire dcache_tlb__entries_WIRE_4_ae_stage2 = dcache_tlb__entries_WIRE_5 [17]; 
    wire dcache_tlb__entries_WIRE_4_ae_final = dcache_tlb__entries_WIRE_5 [18]; 
    wire dcache_tlb__entries_WIRE_4_ae_ptw = dcache_tlb__entries_WIRE_5 [19]; 
    wire dcache_tlb__entries_WIRE_4_g = dcache_tlb__entries_WIRE_5 [20]; 
    wire dcache_tlb__entries_WIRE_4_u = dcache_tlb__entries_WIRE_5 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_4_ppn = dcache_tlb__entries_WIRE_5 [41:22];  
    
    assign  dcache_tlb_entries_barrier_2_io_y_ppn = dcache_tlb_entries_barrier_2_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_2_io_y_u = dcache_tlb_entries_barrier_2_io_x_u ; 
  assign  dcache_tlb_entries_barrier_2_io_y_g = dcache_tlb_entries_barrier_2_io_x_g ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_ptw = dcache_tlb_entries_barrier_2_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_final = dcache_tlb_entries_barrier_2_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ae_stage2 = dcache_tlb_entries_barrier_2_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pf = dcache_tlb_entries_barrier_2_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_2_io_y_gf = dcache_tlb_entries_barrier_2_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sw = dcache_tlb_entries_barrier_2_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sx = dcache_tlb_entries_barrier_2_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_2_io_y_sr = dcache_tlb_entries_barrier_2_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hw = dcache_tlb_entries_barrier_2_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hx = dcache_tlb_entries_barrier_2_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_2_io_y_hr = dcache_tlb_entries_barrier_2_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pw = dcache_tlb_entries_barrier_2_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_2_io_y_px = dcache_tlb_entries_barrier_2_io_x_px ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pr = dcache_tlb_entries_barrier_2_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_2_io_y_ppp = dcache_tlb_entries_barrier_2_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_2_io_y_pal = dcache_tlb_entries_barrier_2_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_2_io_y_paa = dcache_tlb_entries_barrier_2_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_2_io_y_eff = dcache_tlb_entries_barrier_2_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_2_io_y_c = dcache_tlb_entries_barrier_2_io_x_c ; 
  assign  dcache_tlb_entries_barrier_2_io_y_fragmented_superpage = dcache_tlb_entries_barrier_2_io_x_fragmented_superpage ;
     
    wire dcache_tlb__entries_WIRE_6_fragmented_superpage = dcache_tlb__entries_WIRE_7 [0]; 
    wire dcache_tlb__entries_WIRE_6_c = dcache_tlb__entries_WIRE_7 [1]; 
    wire dcache_tlb__entries_WIRE_6_eff = dcache_tlb__entries_WIRE_7 [2]; 
    wire dcache_tlb__entries_WIRE_6_paa = dcache_tlb__entries_WIRE_7 [3]; 
    wire dcache_tlb__entries_WIRE_6_pal = dcache_tlb__entries_WIRE_7 [4]; 
    wire dcache_tlb__entries_WIRE_6_ppp = dcache_tlb__entries_WIRE_7 [5]; 
    wire dcache_tlb__entries_WIRE_6_pr = dcache_tlb__entries_WIRE_7 [6]; 
    wire dcache_tlb__entries_WIRE_6_px = dcache_tlb__entries_WIRE_7 [7]; 
    wire dcache_tlb__entries_WIRE_6_pw = dcache_tlb__entries_WIRE_7 [8]; 
    wire dcache_tlb__entries_WIRE_6_hr = dcache_tlb__entries_WIRE_7 [9]; 
    wire dcache_tlb__entries_WIRE_6_hx = dcache_tlb__entries_WIRE_7 [10]; 
    wire dcache_tlb__entries_WIRE_6_hw = dcache_tlb__entries_WIRE_7 [11]; 
    wire dcache_tlb__entries_WIRE_6_sr = dcache_tlb__entries_WIRE_7 [12]; 
    wire dcache_tlb__entries_WIRE_6_sx = dcache_tlb__entries_WIRE_7 [13]; 
    wire dcache_tlb__entries_WIRE_6_sw = dcache_tlb__entries_WIRE_7 [14]; 
    wire dcache_tlb__entries_WIRE_6_gf = dcache_tlb__entries_WIRE_7 [15]; 
    wire dcache_tlb__entries_WIRE_6_pf = dcache_tlb__entries_WIRE_7 [16]; 
    wire dcache_tlb__entries_WIRE_6_ae_stage2 = dcache_tlb__entries_WIRE_7 [17]; 
    wire dcache_tlb__entries_WIRE_6_ae_final = dcache_tlb__entries_WIRE_7 [18]; 
    wire dcache_tlb__entries_WIRE_6_ae_ptw = dcache_tlb__entries_WIRE_7 [19]; 
    wire dcache_tlb__entries_WIRE_6_g = dcache_tlb__entries_WIRE_7 [20]; 
    wire dcache_tlb__entries_WIRE_6_u = dcache_tlb__entries_WIRE_7 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_6_ppn = dcache_tlb__entries_WIRE_7 [41:22];  
    
    assign  dcache_tlb_entries_barrier_3_io_y_ppn = dcache_tlb_entries_barrier_3_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_3_io_y_u = dcache_tlb_entries_barrier_3_io_x_u ; 
  assign  dcache_tlb_entries_barrier_3_io_y_g = dcache_tlb_entries_barrier_3_io_x_g ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_ptw = dcache_tlb_entries_barrier_3_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_final = dcache_tlb_entries_barrier_3_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ae_stage2 = dcache_tlb_entries_barrier_3_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pf = dcache_tlb_entries_barrier_3_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_3_io_y_gf = dcache_tlb_entries_barrier_3_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sw = dcache_tlb_entries_barrier_3_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sx = dcache_tlb_entries_barrier_3_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_3_io_y_sr = dcache_tlb_entries_barrier_3_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hw = dcache_tlb_entries_barrier_3_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hx = dcache_tlb_entries_barrier_3_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_3_io_y_hr = dcache_tlb_entries_barrier_3_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pw = dcache_tlb_entries_barrier_3_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_3_io_y_px = dcache_tlb_entries_barrier_3_io_x_px ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pr = dcache_tlb_entries_barrier_3_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_3_io_y_ppp = dcache_tlb_entries_barrier_3_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_3_io_y_pal = dcache_tlb_entries_barrier_3_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_3_io_y_paa = dcache_tlb_entries_barrier_3_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_3_io_y_eff = dcache_tlb_entries_barrier_3_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_3_io_y_c = dcache_tlb_entries_barrier_3_io_x_c ; 
  assign  dcache_tlb_entries_barrier_3_io_y_fragmented_superpage = dcache_tlb_entries_barrier_3_io_x_fragmented_superpage ;
     
    wire dcache_tlb__entries_WIRE_8_fragmented_superpage = dcache_tlb__entries_WIRE_9 [0]; 
    wire dcache_tlb__entries_WIRE_8_c = dcache_tlb__entries_WIRE_9 [1]; 
    wire dcache_tlb__entries_WIRE_8_eff = dcache_tlb__entries_WIRE_9 [2]; 
    wire dcache_tlb__entries_WIRE_8_paa = dcache_tlb__entries_WIRE_9 [3]; 
    wire dcache_tlb__entries_WIRE_8_pal = dcache_tlb__entries_WIRE_9 [4]; 
    wire dcache_tlb__entries_WIRE_8_ppp = dcache_tlb__entries_WIRE_9 [5]; 
    wire dcache_tlb__entries_WIRE_8_pr = dcache_tlb__entries_WIRE_9 [6]; 
    wire dcache_tlb__entries_WIRE_8_px = dcache_tlb__entries_WIRE_9 [7]; 
    wire dcache_tlb__entries_WIRE_8_pw = dcache_tlb__entries_WIRE_9 [8]; 
    wire dcache_tlb__entries_WIRE_8_hr = dcache_tlb__entries_WIRE_9 [9]; 
    wire dcache_tlb__entries_WIRE_8_hx = dcache_tlb__entries_WIRE_9 [10]; 
    wire dcache_tlb__entries_WIRE_8_hw = dcache_tlb__entries_WIRE_9 [11]; 
    wire dcache_tlb__entries_WIRE_8_sr = dcache_tlb__entries_WIRE_9 [12]; 
    wire dcache_tlb__entries_WIRE_8_sx = dcache_tlb__entries_WIRE_9 [13]; 
    wire dcache_tlb__entries_WIRE_8_sw = dcache_tlb__entries_WIRE_9 [14]; 
    wire dcache_tlb__entries_WIRE_8_gf = dcache_tlb__entries_WIRE_9 [15]; 
    wire dcache_tlb__entries_WIRE_8_pf = dcache_tlb__entries_WIRE_9 [16]; 
    wire dcache_tlb__entries_WIRE_8_ae_stage2 = dcache_tlb__entries_WIRE_9 [17]; 
    wire dcache_tlb__entries_WIRE_8_ae_final = dcache_tlb__entries_WIRE_9 [18]; 
    wire dcache_tlb__entries_WIRE_8_ae_ptw = dcache_tlb__entries_WIRE_9 [19]; 
    wire dcache_tlb__entries_WIRE_8_g = dcache_tlb__entries_WIRE_9 [20]; 
    wire dcache_tlb__entries_WIRE_8_u = dcache_tlb__entries_WIRE_9 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_8_ppn = dcache_tlb__entries_WIRE_9 [41:22];  
    
    assign  dcache_tlb_entries_barrier_4_io_y_ppn = dcache_tlb_entries_barrier_4_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_4_io_y_u = dcache_tlb_entries_barrier_4_io_x_u ; 
  assign  dcache_tlb_entries_barrier_4_io_y_g = dcache_tlb_entries_barrier_4_io_x_g ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_ptw = dcache_tlb_entries_barrier_4_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_final = dcache_tlb_entries_barrier_4_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ae_stage2 = dcache_tlb_entries_barrier_4_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pf = dcache_tlb_entries_barrier_4_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_4_io_y_gf = dcache_tlb_entries_barrier_4_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sw = dcache_tlb_entries_barrier_4_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sx = dcache_tlb_entries_barrier_4_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_4_io_y_sr = dcache_tlb_entries_barrier_4_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hw = dcache_tlb_entries_barrier_4_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hx = dcache_tlb_entries_barrier_4_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_4_io_y_hr = dcache_tlb_entries_barrier_4_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pw = dcache_tlb_entries_barrier_4_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_4_io_y_px = dcache_tlb_entries_barrier_4_io_x_px ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pr = dcache_tlb_entries_barrier_4_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_4_io_y_ppp = dcache_tlb_entries_barrier_4_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_4_io_y_pal = dcache_tlb_entries_barrier_4_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_4_io_y_paa = dcache_tlb_entries_barrier_4_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_4_io_y_eff = dcache_tlb_entries_barrier_4_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_4_io_y_c = dcache_tlb_entries_barrier_4_io_x_c ; 
  assign  dcache_tlb_entries_barrier_4_io_y_fragmented_superpage = dcache_tlb_entries_barrier_4_io_x_fragmented_superpage ;
     
    wire dcache_tlb__entries_WIRE_10_fragmented_superpage = dcache_tlb__entries_WIRE_11 [0]; 
    wire dcache_tlb__entries_WIRE_10_c = dcache_tlb__entries_WIRE_11 [1]; 
    wire dcache_tlb__entries_WIRE_10_eff = dcache_tlb__entries_WIRE_11 [2]; 
    wire dcache_tlb__entries_WIRE_10_paa = dcache_tlb__entries_WIRE_11 [3]; 
    wire dcache_tlb__entries_WIRE_10_pal = dcache_tlb__entries_WIRE_11 [4]; 
    wire dcache_tlb__entries_WIRE_10_ppp = dcache_tlb__entries_WIRE_11 [5]; 
    wire dcache_tlb__entries_WIRE_10_pr = dcache_tlb__entries_WIRE_11 [6]; 
    wire dcache_tlb__entries_WIRE_10_px = dcache_tlb__entries_WIRE_11 [7]; 
    wire dcache_tlb__entries_WIRE_10_pw = dcache_tlb__entries_WIRE_11 [8]; 
    wire dcache_tlb__entries_WIRE_10_hr = dcache_tlb__entries_WIRE_11 [9]; 
    wire dcache_tlb__entries_WIRE_10_hx = dcache_tlb__entries_WIRE_11 [10]; 
    wire dcache_tlb__entries_WIRE_10_hw = dcache_tlb__entries_WIRE_11 [11]; 
    wire dcache_tlb__entries_WIRE_10_sr = dcache_tlb__entries_WIRE_11 [12]; 
    wire dcache_tlb__entries_WIRE_10_sx = dcache_tlb__entries_WIRE_11 [13]; 
    wire dcache_tlb__entries_WIRE_10_sw = dcache_tlb__entries_WIRE_11 [14]; 
    wire dcache_tlb__entries_WIRE_10_gf = dcache_tlb__entries_WIRE_11 [15]; 
    wire dcache_tlb__entries_WIRE_10_pf = dcache_tlb__entries_WIRE_11 [16]; 
    wire dcache_tlb__entries_WIRE_10_ae_stage2 = dcache_tlb__entries_WIRE_11 [17]; 
    wire dcache_tlb__entries_WIRE_10_ae_final = dcache_tlb__entries_WIRE_11 [18]; 
    wire dcache_tlb__entries_WIRE_10_ae_ptw = dcache_tlb__entries_WIRE_11 [19]; 
    wire dcache_tlb__entries_WIRE_10_g = dcache_tlb__entries_WIRE_11 [20]; 
    wire dcache_tlb__entries_WIRE_10_u = dcache_tlb__entries_WIRE_11 [21]; 
    wire[19:0] dcache_tlb__entries_WIRE_10_ppn = dcache_tlb__entries_WIRE_11 [41:22];  
    
    assign  dcache_tlb_entries_barrier_5_io_y_ppn = dcache_tlb_entries_barrier_5_io_x_ppn ; 
  assign  dcache_tlb_entries_barrier_5_io_y_u = dcache_tlb_entries_barrier_5_io_x_u ; 
  assign  dcache_tlb_entries_barrier_5_io_y_g = dcache_tlb_entries_barrier_5_io_x_g ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_ptw = dcache_tlb_entries_barrier_5_io_x_ae_ptw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_final = dcache_tlb_entries_barrier_5_io_x_ae_final ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ae_stage2 = dcache_tlb_entries_barrier_5_io_x_ae_stage2 ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pf = dcache_tlb_entries_barrier_5_io_x_pf ; 
  assign  dcache_tlb_entries_barrier_5_io_y_gf = dcache_tlb_entries_barrier_5_io_x_gf ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sw = dcache_tlb_entries_barrier_5_io_x_sw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sx = dcache_tlb_entries_barrier_5_io_x_sx ; 
  assign  dcache_tlb_entries_barrier_5_io_y_sr = dcache_tlb_entries_barrier_5_io_x_sr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hw = dcache_tlb_entries_barrier_5_io_x_hw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hx = dcache_tlb_entries_barrier_5_io_x_hx ; 
  assign  dcache_tlb_entries_barrier_5_io_y_hr = dcache_tlb_entries_barrier_5_io_x_hr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pw = dcache_tlb_entries_barrier_5_io_x_pw ; 
  assign  dcache_tlb_entries_barrier_5_io_y_px = dcache_tlb_entries_barrier_5_io_x_px ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pr = dcache_tlb_entries_barrier_5_io_x_pr ; 
  assign  dcache_tlb_entries_barrier_5_io_y_ppp = dcache_tlb_entries_barrier_5_io_x_ppp ; 
  assign  dcache_tlb_entries_barrier_5_io_y_pal = dcache_tlb_entries_barrier_5_io_x_pal ; 
  assign  dcache_tlb_entries_barrier_5_io_y_paa = dcache_tlb_entries_barrier_5_io_x_paa ; 
  assign  dcache_tlb_entries_barrier_5_io_y_eff = dcache_tlb_entries_barrier_5_io_x_eff ; 
  assign  dcache_tlb_entries_barrier_5_io_y_c = dcache_tlb_entries_barrier_5_io_x_c ; 
  assign  dcache_tlb_entries_barrier_5_io_y_fragmented_superpage = dcache_tlb_entries_barrier_5_io_x_fragmented_superpage ;
     
    wire[19:0] dcache_tlb_ppn =( dcache_tlb_hitsVec_0  ?  dcache__tlb_entries_barrier_io_y_ppn :20'h0)|( dcache_tlb_hitsVec_1  ?  dcache__tlb_entries_barrier_1_io_y_ppn :20'h0)|( dcache_tlb_hitsVec_2  ?  dcache__tlb_entries_barrier_2_io_y_ppn :20'h0)|( dcache_tlb_hitsVec_3  ?  dcache__tlb_entries_barrier_3_io_y_ppn :20'h0)|( dcache_tlb_hitsVec_4  ?  dcache__tlb_entries_barrier_4_io_y_ppn :20'h0)|( dcache_tlb_hitsVec_5  ?  dcache__tlb_entries_barrier_5_io_y_ppn :20'h0)|( dcache_tlb_vm_enabled ==1'h0 ?  dcache_tlb_vpn [19:0]:20'h0); 
    wire[1:0] dcache_tlb_ptw_ae_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_ptw , dcache__tlb_entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] dcache_tlb_ptw_ae_array_lo ={ dcache_tlb_ptw_ae_array_lo_hi , dcache__tlb_entries_barrier_io_y_ae_ptw }; 
    wire[1:0] dcache_tlb_ptw_ae_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_ptw , dcache__tlb_entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] dcache_tlb_ptw_ae_array_hi ={ dcache_tlb_ptw_ae_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] dcache_tlb_ptw_ae_array ={1'h0,{ dcache_tlb_ptw_ae_array_hi , dcache_tlb_ptw_ae_array_lo }}; 
    wire[1:0] dcache_tlb_final_ae_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_final , dcache__tlb_entries_barrier_1_io_y_ae_final }; 
    wire[2:0] dcache_tlb_final_ae_array_lo ={ dcache_tlb_final_ae_array_lo_hi , dcache__tlb_entries_barrier_io_y_ae_final }; 
    wire[1:0] dcache_tlb_final_ae_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_final , dcache__tlb_entries_barrier_4_io_y_ae_final }; 
    wire[2:0] dcache_tlb_final_ae_array_hi ={ dcache_tlb_final_ae_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_final }; 
    wire[6:0] dcache_tlb_final_ae_array ={1'h0,{ dcache_tlb_final_ae_array_hi , dcache_tlb_final_ae_array_lo }}; 
    wire[1:0] dcache_tlb_ptw_pf_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_pf , dcache__tlb_entries_barrier_1_io_y_pf }; 
    wire[2:0] dcache_tlb_ptw_pf_array_lo ={ dcache_tlb_ptw_pf_array_lo_hi , dcache__tlb_entries_barrier_io_y_pf }; 
    wire[1:0] dcache_tlb_ptw_pf_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_pf , dcache__tlb_entries_barrier_4_io_y_pf }; 
    wire[2:0] dcache_tlb_ptw_pf_array_hi ={ dcache_tlb_ptw_pf_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_pf }; 
    wire[6:0] dcache_tlb_ptw_pf_array ={1'h0,{ dcache_tlb_ptw_pf_array_hi , dcache_tlb_ptw_pf_array_lo }}; 
    wire[1:0] dcache_tlb_ptw_gf_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_gf , dcache__tlb_entries_barrier_1_io_y_gf }; 
    wire[2:0] dcache_tlb_ptw_gf_array_lo ={ dcache_tlb_ptw_gf_array_lo_hi , dcache__tlb_entries_barrier_io_y_gf }; 
    wire[1:0] dcache_tlb_ptw_gf_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_gf , dcache__tlb_entries_barrier_4_io_y_gf }; 
    wire[2:0] dcache_tlb_ptw_gf_array_hi ={ dcache_tlb_ptw_gf_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_gf }; 
    wire[6:0] dcache_tlb_ptw_gf_array ={1'h0,{ dcache_tlb_ptw_gf_array_hi , dcache_tlb_ptw_gf_array_lo }}; 
    wire dcache_tlb_sum = dcache_tlb_priv_v  ?  dcache_tlb_io_ptw_gstatus_sum : dcache_tlb_io_ptw_status_sum ; 
    wire[1:0] dcache_tlb_priv_rw_ok_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_u , dcache__tlb_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_lo ={ dcache_tlb_priv_rw_ok_lo_hi , dcache__tlb_entries_barrier_io_y_u }; 
    wire[1:0] dcache_tlb_priv_rw_ok_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_u , dcache__tlb_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_hi ={ dcache_tlb_priv_rw_ok_hi_hi , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[1:0] dcache_tlb_priv_rw_ok_lo_hi_1 ={ dcache__tlb_entries_barrier_2_io_y_u , dcache__tlb_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_lo_1 ={ dcache_tlb_priv_rw_ok_lo_hi_1 , dcache__tlb_entries_barrier_io_y_u }; 
    wire[1:0] dcache_tlb_priv_rw_ok_hi_hi_1 ={ dcache__tlb_entries_barrier_5_io_y_u , dcache__tlb_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_tlb_priv_rw_ok_hi_1 ={ dcache_tlb_priv_rw_ok_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_tlb_priv_rw_ok =( dcache_tlb_priv_s ==1'h0| dcache_tlb_sum  ? { dcache_tlb_priv_rw_ok_hi , dcache_tlb_priv_rw_ok_lo }:6'h0)|( dcache_tlb_priv_s  ? ~{ dcache_tlb_priv_rw_ok_hi_1 , dcache_tlb_priv_rw_ok_lo_1 }:6'h0); 
    wire[1:0] dcache_tlb_priv_x_ok_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_u , dcache__tlb_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_lo ={ dcache_tlb_priv_x_ok_lo_hi , dcache__tlb_entries_barrier_io_y_u }; 
    wire[1:0] dcache_tlb_priv_x_ok_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_u , dcache__tlb_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_hi ={ dcache_tlb_priv_x_ok_hi_hi , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[1:0] dcache_tlb_priv_x_ok_lo_hi_1 ={ dcache__tlb_entries_barrier_2_io_y_u , dcache__tlb_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_lo_1 ={ dcache_tlb_priv_x_ok_lo_hi_1 , dcache__tlb_entries_barrier_io_y_u }; 
    wire[1:0] dcache_tlb_priv_x_ok_hi_hi_1 ={ dcache__tlb_entries_barrier_5_io_y_u , dcache__tlb_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_tlb_priv_x_ok_hi_1 ={ dcache_tlb_priv_x_ok_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_tlb_priv_x_ok = dcache_tlb_priv_s  ? ~{ dcache_tlb_priv_x_ok_hi , dcache_tlb_priv_x_ok_lo }:{ dcache_tlb_priv_x_ok_hi_1 , dcache_tlb_priv_x_ok_lo_1 }; 
    wire[1:0] dcache_tlb_stage1_bypass_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_ae_stage2 , dcache__tlb_entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] dcache_tlb_stage1_bypass_lo ={ dcache_tlb_stage1_bypass_lo_hi , dcache__tlb_entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] dcache_tlb_stage1_bypass_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_ae_stage2 , dcache__tlb_entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] dcache_tlb_stage1_bypass_hi ={ dcache_tlb_stage1_bypass_hi_hi , dcache__tlb_entries_barrier_3_io_y_ae_stage2 }; 
    wire dcache_tlb_mxr = dcache_tlb_io_ptw_status_mxr |( dcache_tlb_priv_v  ?  dcache_tlb_io_ptw_gstatus_mxr :1'h0); 
    wire[1:0] dcache_tlb_r_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_sr , dcache__tlb_entries_barrier_1_io_y_sr }; 
    wire[2:0] dcache_tlb_r_array_lo ={ dcache_tlb_r_array_lo_hi , dcache__tlb_entries_barrier_io_y_sr }; 
    wire[1:0] dcache_tlb_r_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_sr , dcache__tlb_entries_barrier_4_io_y_sr }; 
    wire[2:0] dcache_tlb_r_array_hi ={ dcache_tlb_r_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sr }; 
    wire[1:0] dcache_tlb_r_array_lo_hi_1 ={ dcache__tlb_entries_barrier_2_io_y_sx , dcache__tlb_entries_barrier_1_io_y_sx }; 
    wire[2:0] dcache_tlb_r_array_lo_1 ={ dcache_tlb_r_array_lo_hi_1 , dcache__tlb_entries_barrier_io_y_sx }; 
    wire[1:0] dcache_tlb_r_array_hi_hi_1 ={ dcache__tlb_entries_barrier_5_io_y_sx , dcache__tlb_entries_barrier_4_io_y_sx }; 
    wire[2:0] dcache_tlb_r_array_hi_1 ={ dcache_tlb_r_array_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_tlb_r_array ={1'h1, dcache_tlb_priv_rw_ok &({ dcache_tlb_r_array_hi , dcache_tlb_r_array_lo }|( dcache_tlb_mxr  ? { dcache_tlb_r_array_hi_1 , dcache_tlb_r_array_lo_1 }:6'h0))| dcache_tlb_stage1_bypass }; 
    wire[1:0] dcache_tlb_w_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_sw , dcache__tlb_entries_barrier_1_io_y_sw }; 
    wire[2:0] dcache_tlb_w_array_lo ={ dcache_tlb_w_array_lo_hi , dcache__tlb_entries_barrier_io_y_sw }; 
    wire[1:0] dcache_tlb_w_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_sw , dcache__tlb_entries_barrier_4_io_y_sw }; 
    wire[2:0] dcache_tlb_w_array_hi ={ dcache_tlb_w_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sw }; 
    wire[6:0] dcache_tlb_w_array ={1'h1, dcache_tlb_priv_rw_ok &{ dcache_tlb_w_array_hi , dcache_tlb_w_array_lo }| dcache_tlb_stage1_bypass }; 
    wire[1:0] dcache_tlb_x_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_sx , dcache__tlb_entries_barrier_1_io_y_sx }; 
    wire[2:0] dcache_tlb_x_array_lo ={ dcache_tlb_x_array_lo_hi , dcache__tlb_entries_barrier_io_y_sx }; 
    wire[1:0] dcache_tlb_x_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_sx , dcache__tlb_entries_barrier_4_io_y_sx }; 
    wire[2:0] dcache_tlb_x_array_hi ={ dcache_tlb_x_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_tlb_x_array ={1'h1, dcache_tlb_priv_x_ok &{ dcache_tlb_x_array_hi , dcache_tlb_x_array_lo }| dcache_tlb_stage1_bypass }; 
    wire[5:0] dcache_tlb_stage2_bypass = dcache_tlb_stage2_en ==1'h0 ? 6'h3F:6'h0; 
    wire[1:0] dcache_tlb_hr_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_hr , dcache__tlb_entries_barrier_1_io_y_hr }; 
    wire[2:0] dcache_tlb_hr_array_lo ={ dcache_tlb_hr_array_lo_hi , dcache__tlb_entries_barrier_io_y_hr }; 
    wire[1:0] dcache_tlb_hr_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_hr , dcache__tlb_entries_barrier_4_io_y_hr }; 
    wire[2:0] dcache_tlb_hr_array_hi ={ dcache_tlb_hr_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hr }; 
    wire[1:0] dcache_tlb_hr_array_lo_hi_1 ={ dcache__tlb_entries_barrier_2_io_y_hx , dcache__tlb_entries_barrier_1_io_y_hx }; 
    wire[2:0] dcache_tlb_hr_array_lo_1 ={ dcache_tlb_hr_array_lo_hi_1 , dcache__tlb_entries_barrier_io_y_hx }; 
    wire[1:0] dcache_tlb_hr_array_hi_hi_1 ={ dcache__tlb_entries_barrier_5_io_y_hx , dcache__tlb_entries_barrier_4_io_y_hx }; 
    wire[2:0] dcache_tlb_hr_array_hi_1 ={ dcache_tlb_hr_array_hi_hi_1 , dcache__tlb_entries_barrier_3_io_y_hx }; 
    wire[6:0] dcache_tlb_hr_array ={1'h1,{ dcache_tlb_hr_array_hi , dcache_tlb_hr_array_lo }|( dcache_tlb_io_ptw_status_mxr  ? { dcache_tlb_hr_array_hi_1 , dcache_tlb_hr_array_lo_1 }:6'h0)| dcache_tlb_stage2_bypass }; 
    wire[1:0] dcache_tlb_hw_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_hw , dcache__tlb_entries_barrier_1_io_y_hw }; 
    wire[2:0] dcache_tlb_hw_array_lo ={ dcache_tlb_hw_array_lo_hi , dcache__tlb_entries_barrier_io_y_hw }; 
    wire[1:0] dcache_tlb_hw_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_hw , dcache__tlb_entries_barrier_4_io_y_hw }; 
    wire[2:0] dcache_tlb_hw_array_hi ={ dcache_tlb_hw_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hw }; 
    wire[6:0] dcache_tlb_hw_array ={1'h1,{ dcache_tlb_hw_array_hi , dcache_tlb_hw_array_lo }| dcache_tlb_stage2_bypass }; 
    wire[1:0] dcache_tlb_hx_array_lo_hi ={ dcache__tlb_entries_barrier_2_io_y_hx , dcache__tlb_entries_barrier_1_io_y_hx }; 
    wire[2:0] dcache_tlb_hx_array_lo ={ dcache_tlb_hx_array_lo_hi , dcache__tlb_entries_barrier_io_y_hx }; 
    wire[1:0] dcache_tlb_hx_array_hi_hi ={ dcache__tlb_entries_barrier_5_io_y_hx , dcache__tlb_entries_barrier_4_io_y_hx }; 
    wire[2:0] dcache_tlb_hx_array_hi ={ dcache_tlb_hx_array_hi_hi , dcache__tlb_entries_barrier_3_io_y_hx }; 
    wire[6:0] dcache_tlb_hx_array ={1'h1,{ dcache_tlb_hx_array_hi , dcache_tlb_hx_array_lo }| dcache_tlb_stage2_bypass }; 
    wire[1:0] dcache_tlb_pr_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pr , dcache__tlb_entries_barrier_io_y_pr }; 
    wire[1:0] dcache_tlb_pr_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pr , dcache__tlb_entries_barrier_3_io_y_pr }; 
    wire[2:0] dcache_tlb_pr_array_hi ={ dcache_tlb_pr_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pr }; 
    wire[6:0] dcache_tlb_pr_array ={ dcache_tlb_prot_r  ? 2'h3:2'h0,{ dcache_tlb_pr_array_hi , dcache_tlb_pr_array_lo }}&~( dcache_tlb_ptw_ae_array | dcache_tlb_final_ae_array ); 
    wire[1:0] dcache_tlb_pw_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pw , dcache__tlb_entries_barrier_io_y_pw }; 
    wire[1:0] dcache_tlb_pw_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pw , dcache__tlb_entries_barrier_3_io_y_pw }; 
    wire[2:0] dcache_tlb_pw_array_hi ={ dcache_tlb_pw_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pw }; 
    wire[6:0] dcache_tlb_pw_array ={ dcache_tlb_prot_w  ? 2'h3:2'h0,{ dcache_tlb_pw_array_hi , dcache_tlb_pw_array_lo }}&~( dcache_tlb_ptw_ae_array | dcache_tlb_final_ae_array ); 
    wire[1:0] dcache_tlb_px_array_lo ={ dcache__tlb_entries_barrier_1_io_y_px , dcache__tlb_entries_barrier_io_y_px }; 
    wire[1:0] dcache_tlb_px_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_px , dcache__tlb_entries_barrier_3_io_y_px }; 
    wire[2:0] dcache_tlb_px_array_hi ={ dcache_tlb_px_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_px }; 
    wire[6:0] dcache_tlb_px_array ={ dcache_tlb_prot_x  ? 2'h3:2'h0,{ dcache_tlb_px_array_hi , dcache_tlb_px_array_lo }}&~( dcache_tlb_ptw_ae_array | dcache_tlb_final_ae_array ); 
    wire[1:0] dcache_tlb_eff_array_lo ={ dcache__tlb_entries_barrier_1_io_y_eff , dcache__tlb_entries_barrier_io_y_eff }; 
    wire[1:0] dcache_tlb_eff_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_eff , dcache__tlb_entries_barrier_3_io_y_eff }; 
    wire[2:0] dcache_tlb_eff_array_hi ={ dcache_tlb_eff_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_eff }; 
    wire[6:0] dcache_tlb_eff_array ={ dcache_tlb_prot_eff  ? 2'h3:2'h0,{ dcache_tlb_eff_array_hi , dcache_tlb_eff_array_lo }}; 
    wire[1:0] dcache_tlb_c_array_lo ={ dcache__tlb_entries_barrier_1_io_y_c , dcache__tlb_entries_barrier_io_y_c }; 
    wire[1:0] dcache_tlb_c_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_c , dcache__tlb_entries_barrier_3_io_y_c }; 
    wire[2:0] dcache_tlb_c_array_hi ={ dcache_tlb_c_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_tlb_c_array ={ dcache_tlb_cacheable  ? 2'h3:2'h0,{ dcache_tlb_c_array_hi , dcache_tlb_c_array_lo }}; 
    wire[6:0] dcache_tlb_lrscAllowed = dcache_tlb_c_array ; 
    wire[1:0] dcache_tlb_ppp_array_lo ={ dcache__tlb_entries_barrier_1_io_y_ppp , dcache__tlb_entries_barrier_io_y_ppp }; 
    wire[1:0] dcache_tlb_ppp_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_ppp , dcache__tlb_entries_barrier_3_io_y_ppp }; 
    wire[2:0] dcache_tlb_ppp_array_hi ={ dcache_tlb_ppp_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_ppp }; 
    wire[6:0] dcache_tlb_ppp_array ={ dcache_tlb_prot_pp  ? 2'h3:2'h0,{ dcache_tlb_ppp_array_hi , dcache_tlb_ppp_array_lo }}; 
    wire[1:0] dcache_tlb_paa_array_lo ={ dcache__tlb_entries_barrier_1_io_y_paa , dcache__tlb_entries_barrier_io_y_paa }; 
    wire[1:0] dcache_tlb_paa_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_paa , dcache__tlb_entries_barrier_3_io_y_paa }; 
    wire[2:0] dcache_tlb_paa_array_hi ={ dcache_tlb_paa_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_paa }; 
    wire[6:0] dcache_tlb_paa_array ={ dcache_tlb_prot_aa  ? 2'h3:2'h0,{ dcache_tlb_paa_array_hi , dcache_tlb_paa_array_lo }}; 
    wire[1:0] dcache_tlb_pal_array_lo ={ dcache__tlb_entries_barrier_1_io_y_pal , dcache__tlb_entries_barrier_io_y_pal }; 
    wire[1:0] dcache_tlb_pal_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_pal , dcache__tlb_entries_barrier_3_io_y_pal }; 
    wire[2:0] dcache_tlb_pal_array_hi ={ dcache_tlb_pal_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_pal }; 
    wire[6:0] dcache_tlb_pal_array ={ dcache_tlb_prot_al  ? 2'h3:2'h0,{ dcache_tlb_pal_array_hi , dcache_tlb_pal_array_lo }}; 
    wire[6:0] dcache_tlb_ppp_array_if_cached = dcache_tlb_ppp_array | dcache_tlb_c_array ; 
    wire[6:0] dcache_tlb_paa_array_if_cached = dcache_tlb_paa_array | dcache_tlb_c_array ; 
    wire[6:0] dcache_tlb_pal_array_if_cached = dcache_tlb_pal_array | dcache_tlb_c_array ; 
    wire[1:0] dcache_tlb_prefetchable_array_lo ={ dcache__tlb_entries_barrier_1_io_y_c , dcache__tlb_entries_barrier_io_y_c }; 
    wire[1:0] dcache_tlb_prefetchable_array_hi_hi ={ dcache__tlb_entries_barrier_4_io_y_c , dcache__tlb_entries_barrier_3_io_y_c }; 
    wire[2:0] dcache_tlb_prefetchable_array_hi ={ dcache_tlb_prefetchable_array_hi_hi , dcache__tlb_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_tlb_prefetchable_array ={{ dcache_tlb_cacheable & dcache_tlb_homogeneous ,1'h0},{ dcache_tlb_prefetchable_array_hi , dcache_tlb_prefetchable_array_lo }}; 
    wire[4:0] dcache__GEN_34 ={1'h0,4'h1<< dcache_tlb_io_req_bits_size }-5'h1; 
    wire dcache_tlb_misaligned =|( dcache_tlb_io_req_bits_vaddr &{30'h0, dcache__GEN_34 [3:0]}); 
    wire[4:0] dcache_tlb_io_req_bits_cmd ; 
    wire dcache_tlb_cmd_lrsc =( dcache_tlb_io_req_bits_cmd ==5'h6| dcache_tlb_io_req_bits_cmd ==5'h7)&1'h1; 
    wire dcache_tlb_cmd_amo_logical =( dcache_tlb_io_req_bits_cmd ==5'h4| dcache_tlb_io_req_bits_cmd ==5'h9| dcache_tlb_io_req_bits_cmd ==5'hA| dcache_tlb_io_req_bits_cmd ==5'hB)&1'h1; 
    wire dcache_tlb_cmd_amo_arithmetic =( dcache_tlb_io_req_bits_cmd ==5'h8| dcache_tlb_io_req_bits_cmd ==5'hC| dcache_tlb_io_req_bits_cmd ==5'hD| dcache_tlb_io_req_bits_cmd ==5'hE| dcache_tlb_io_req_bits_cmd ==5'hF)&1'h1; 
    wire dcache_tlb_cmd_put_partial = dcache_tlb_io_req_bits_cmd ==5'h11; 
    wire dcache_tlb_cmd_read = dcache_tlb_io_req_bits_cmd ==5'h0| dcache_tlb_io_req_bits_cmd ==5'h10| dcache_tlb_io_req_bits_cmd ==5'h6| dcache_tlb_io_req_bits_cmd ==5'h7| dcache_tlb_io_req_bits_cmd ==5'h4| dcache_tlb_io_req_bits_cmd ==5'h9| dcache_tlb_io_req_bits_cmd ==5'hA| dcache_tlb_io_req_bits_cmd ==5'hB| dcache_tlb_io_req_bits_cmd ==5'h8| dcache_tlb_io_req_bits_cmd ==5'hC| dcache_tlb_io_req_bits_cmd ==5'hD| dcache_tlb_io_req_bits_cmd ==5'hE| dcache_tlb_io_req_bits_cmd ==5'hF; 
    wire dcache_tlb_cmd_write = dcache_tlb_io_req_bits_cmd ==5'h1| dcache_tlb_io_req_bits_cmd ==5'h11| dcache_tlb_io_req_bits_cmd ==5'h7| dcache_tlb_io_req_bits_cmd ==5'h4| dcache_tlb_io_req_bits_cmd ==5'h9| dcache_tlb_io_req_bits_cmd ==5'hA| dcache_tlb_io_req_bits_cmd ==5'hB| dcache_tlb_io_req_bits_cmd ==5'h8| dcache_tlb_io_req_bits_cmd ==5'hC| dcache_tlb_io_req_bits_cmd ==5'hD| dcache_tlb_io_req_bits_cmd ==5'hE| dcache_tlb_io_req_bits_cmd ==5'hF; 
    wire dcache_tlb_cmd_write_perms = dcache_tlb_cmd_write | dcache_tlb_io_req_bits_cmd ==5'h5| dcache_tlb_io_req_bits_cmd ==5'h17; 
    wire[6:0] dcache_tlb_ae_array =( dcache_tlb_misaligned  ?  dcache_tlb_eff_array :7'h0)|( dcache_tlb_cmd_lrsc  ? ~ dcache_tlb_lrscAllowed :7'h0); 
    wire[6:0] dcache_tlb_ae_ld_array = dcache_tlb_cmd_read  ?  dcache_tlb_ae_array |~ dcache_tlb_pr_array :7'h0; 
    wire[6:0] dcache_tlb_ae_st_array =( dcache_tlb_cmd_write_perms  ?  dcache_tlb_ae_array |~ dcache_tlb_pw_array :7'h0)|( dcache_tlb_cmd_put_partial  ? ~ dcache_tlb_ppp_array_if_cached :7'h0)|( dcache_tlb_cmd_amo_logical  ? ~ dcache_tlb_pal_array_if_cached :7'h0)|( dcache_tlb_cmd_amo_arithmetic  ? ~ dcache_tlb_paa_array_if_cached :7'h0); 
    wire[6:0] dcache_tlb_must_alloc_array =( dcache_tlb_cmd_put_partial  ? ~ dcache_tlb_ppp_array :7'h0)|( dcache_tlb_cmd_amo_logical  ? ~ dcache_tlb_pal_array :7'h0)|( dcache_tlb_cmd_amo_arithmetic  ? ~ dcache_tlb_paa_array :7'h0)|( dcache_tlb_cmd_lrsc  ? 7'h7F:7'h0); 
    wire[6:0] dcache_tlb_pf_ld_array = dcache_tlb_cmd_read  ? (~( dcache_tlb_cmd_readx  ?  dcache_tlb_x_array : dcache_tlb_r_array )&~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array :7'h0; 
    wire[6:0] dcache_tlb_pf_st_array = dcache_tlb_cmd_write_perms  ? (~ dcache_tlb_w_array &~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array :7'h0; 
    wire[6:0] dcache_tlb_pf_inst_array =(~ dcache_tlb_x_array &~ dcache_tlb_ptw_ae_array | dcache_tlb_ptw_pf_array )&~ dcache_tlb_ptw_gf_array ; 
    wire[6:0] dcache_tlb_gf_ld_array = dcache_tlb_priv_v & dcache_tlb_cmd_read  ? (~( dcache_tlb_cmd_readx  ?  dcache_tlb_hx_array : dcache_tlb_hr_array )| dcache_tlb_ptw_gf_array )&~ dcache_tlb_ptw_ae_array :7'h0; 
    wire[6:0] dcache_tlb_gf_st_array = dcache_tlb_priv_v & dcache_tlb_cmd_write_perms  ? (~ dcache_tlb_hw_array | dcache_tlb_ptw_gf_array )&~ dcache_tlb_ptw_ae_array :7'h0; 
    wire[6:0] dcache_tlb_gf_inst_array = dcache_tlb_priv_v  ? (~ dcache_tlb_hx_array | dcache_tlb_ptw_gf_array )&~ dcache_tlb_ptw_ae_array :7'h0; 
    wire[6:0] dcache_tlb_gpa_hits_need_gpa_mask = dcache_tlb_gf_ld_array | dcache_tlb_gf_st_array ; 
    wire[5:0] dcache_tlb_gpa_hits_hit_mask ={1'h0, dcache_tlb_r_gpa_valid & dcache_tlb_r_gpa_vpn == dcache_tlb_vpn  ? 5'h1F:5'h0}|( dcache_tlb_vstage1_en ==1'h0 ? 6'h3F:6'h0); 
    wire[5:0] dcache_tlb_gpa_hits = dcache_tlb_gpa_hits_hit_mask |~( dcache_tlb_gpa_hits_need_gpa_mask [5:0]); 
    wire dcache_tlb_tlb_hit_if_not_gpa_miss =| dcache_tlb_real_hits ; 
    wire dcache_tlb_tlb_hit =|( dcache_tlb_real_hits & dcache_tlb_gpa_hits ); 
    wire dcache_tlb_tlb_miss = dcache_tlb_vm_enabled & dcache_tlb_vsatp_mode_mismatch ==1'h0& dcache_tlb_tlb_hit ==1'h0; reg[2:0] dcache_tlb_state_reg_1 ; 
    wire dcache_tlb_io_req_valid ; 
    wire dcache__GEN_35 = dcache_tlb_io_req_valid & dcache_tlb_vm_enabled ; 
    wire dcache__GEN_36 = dcache_tlb_superpage_hits_0 | dcache_tlb_superpage_hits_1 | dcache_tlb_superpage_hits_2 | dcache_tlb_superpage_hits_3 ; 
    wire[1:0] dcache_tlb_lo ={ dcache_tlb_superpage_hits_1 , dcache_tlb_superpage_hits_0 }; 
    wire[1:0] dcache_tlb_hi ={ dcache_tlb_superpage_hits_3 , dcache_tlb_superpage_hits_2 }; 
    wire[3:0] dcache__GEN_37 ={ dcache_tlb_hi , dcache_tlb_lo }; 
    wire[1:0] dcache_tlb_hi_1 = dcache__GEN_37 [3:2]; 
    wire[1:0] dcache_tlb_lo_1 = dcache__GEN_37 [1:0]; 
    wire[1:0] dcache__GEN_38 = dcache_tlb_hi_1 | dcache_tlb_lo_1 ; 
    wire[1:0] dcache_tlb_state_reg_touch_way_sized ={| dcache_tlb_hi_1 , dcache__GEN_38 [1]}; 
    wire dcache_tlb_state_reg_set_left_older = dcache_tlb_state_reg_touch_way_sized [1]==1'h0; 
    wire dcache_tlb_state_reg_left_subtree_state = dcache_tlb_state_reg_1 [1]; 
    wire dcache_tlb_state_reg_right_subtree_state = dcache_tlb_state_reg_1 [0]; 
    wire[1:0] dcache_tlb_state_reg_hi ={ dcache_tlb_state_reg_set_left_older , dcache_tlb_state_reg_set_left_older  ?  dcache_tlb_state_reg_left_subtree_state : dcache_tlb_state_reg_touch_way_sized [0]==1'h0}; 
    wire[2:0] dcache__GEN_39 ={ dcache_tlb_state_reg_hi , dcache_tlb_state_reg_set_left_older  ?  dcache_tlb_state_reg_touch_way_sized [0]==1'h0: dcache_tlb_state_reg_right_subtree_state }; 
    wire[2:0] dcache__tlb_real_hits_2to0 = dcache_tlb_real_hits [2:0]; 
    wire dcache_tlb_multipleHits_leftOne = dcache__tlb_real_hits_2to0 [0]; 
    wire[1:0] dcache__tlb_real_hits_2to0_2to1 = dcache__tlb_real_hits_2to0 [2:1]; 
    wire dcache_tlb_multipleHits_leftOne_1 = dcache__tlb_real_hits_2to0_2to1 [0]; 
    wire dcache_tlb_multipleHits_rightOne = dcache__tlb_real_hits_2to0_2to1 [1]; 
    wire dcache_tlb_multipleHits_rightOne_1 = dcache_tlb_multipleHits_leftOne_1 | dcache_tlb_multipleHits_rightOne ; 
    wire dcache_tlb_multipleHits_rightTwo = dcache_tlb_multipleHits_leftOne_1 & dcache_tlb_multipleHits_rightOne |1'h0; 
    wire dcache_tlb_multipleHits_leftOne_2 = dcache_tlb_multipleHits_leftOne | dcache_tlb_multipleHits_rightOne_1 ; 
    wire dcache_tlb_multipleHits_leftTwo = dcache_tlb_multipleHits_rightTwo |1'h0| dcache_tlb_multipleHits_leftOne & dcache_tlb_multipleHits_rightOne_1 ; 
    wire[2:0] dcache__tlb_real_hits_5to3 = dcache_tlb_real_hits [5:3]; 
    wire dcache_tlb_multipleHits_leftOne_3 = dcache__tlb_real_hits_5to3 [0]; 
    wire[1:0] dcache__tlb_real_hits_5to3_2to1 = dcache__tlb_real_hits_5to3 [2:1]; 
    wire dcache_tlb_multipleHits_leftOne_4 = dcache__tlb_real_hits_5to3_2to1 [0]; 
    wire dcache_tlb_multipleHits_rightOne_2 = dcache__tlb_real_hits_5to3_2to1 [1]; 
    wire dcache_tlb_multipleHits_rightOne_3 = dcache_tlb_multipleHits_leftOne_4 | dcache_tlb_multipleHits_rightOne_2 ; 
    wire dcache_tlb_multipleHits_rightTwo_1 = dcache_tlb_multipleHits_leftOne_4 & dcache_tlb_multipleHits_rightOne_2 |1'h0; 
    wire dcache_tlb_multipleHits_rightOne_4 = dcache_tlb_multipleHits_leftOne_3 | dcache_tlb_multipleHits_rightOne_3 ; 
    wire dcache_tlb_multipleHits_rightTwo_2 = dcache_tlb_multipleHits_rightTwo_1 |1'h0| dcache_tlb_multipleHits_leftOne_3 & dcache_tlb_multipleHits_rightOne_3 ; 
    wire dcache_tlb_multipleHits = dcache_tlb_multipleHits_leftTwo | dcache_tlb_multipleHits_rightTwo_2 | dcache_tlb_multipleHits_leftOne_2 & dcache_tlb_multipleHits_rightOne_4 ; 
    wire dcache_tlb_io_req_ready = dcache_tlb_state ==2'h0; 
    wire dcache_tlb_io_resp_pf_ld =(|( dcache_tlb_pf_ld_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_pf_st =(|( dcache_tlb_pf_st_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_pf_inst =(|( dcache_tlb_pf_inst_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_gf_ld =(|( dcache_tlb_gf_ld_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_gf_st =(|( dcache_tlb_gf_st_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_gf_inst =(|( dcache_tlb_gf_inst_array & dcache_tlb_hits ))|1'h0; 
    wire dcache_tlb_io_resp_ae_ld =|( dcache_tlb_ae_ld_array & dcache_tlb_hits ); 
    wire dcache_tlb_io_resp_ae_st =|( dcache_tlb_ae_st_array & dcache_tlb_hits ); 
    wire dcache_tlb_io_resp_ae_inst =|(~ dcache_tlb_px_array & dcache_tlb_hits ); 
    wire dcache_tlb_io_resp_ma_ld = dcache_tlb_misaligned & dcache_tlb_cmd_read ; 
    wire dcache_tlb_io_resp_ma_st = dcache_tlb_misaligned & dcache_tlb_cmd_write ; 
    wire dcache_tlb_io_resp_cacheable =|( dcache_tlb_c_array & dcache_tlb_hits ); 
    wire dcache_tlb_io_resp_must_alloc =|( dcache_tlb_must_alloc_array & dcache_tlb_hits ); 
    wire dcache_tlb_io_resp_miss = dcache_tlb_do_refill | dcache_tlb_vsatp_mode_mismatch | dcache_tlb_tlb_miss | dcache_tlb_multipleHits ; 
    wire[31:0] dcache_tlb_io_resp_paddr ={ dcache_tlb_ppn , dcache_tlb_io_req_bits_vaddr [11:0]}; 
    wire dcache_tlb_io_resp_gpa_is_pte = dcache_tlb_vstage1_en & dcache_tlb_r_gpa_is_pte ; 
    wire[21:0] dcache_tlb_io_resp_gpa_page = dcache_tlb_vstage1_en ==1'h0 ? {1'h0, dcache_tlb_vpn }:{1'h0, dcache_tlb_r_gpa [32:12]}; 
    wire[11:0] dcache_tlb_io_resp_gpa_offset = dcache_tlb_io_resp_gpa_is_pte  ?  dcache_tlb_r_gpa [11:0]: dcache_tlb_io_req_bits_vaddr [11:0]; 
    wire[33:0] dcache_tlb_io_resp_gpa ={ dcache_tlb_io_resp_gpa_page , dcache_tlb_io_resp_gpa_offset }; 
  assign  dcache_tlb_io_ptw_req_valid = dcache_tlb_state ==2'h1; 
    wire dcache_tlb_io_kill ; 
    wire dcache_tlb_io_ptw_req_bits_valid = dcache_tlb_io_kill ==1'h0; 
    wire dcache_pma_checker_newEntry_ae_ptw = dcache_pma_checker_io_ptw_resp_bits_ae_ptw ; 
    wire dcache_pma_checker_newEntry_ae_final = dcache_pma_checker_io_ptw_resp_bits_ae_final ; 
    wire dcache_pma_checker_newEntry_pf = dcache_pma_checker_io_ptw_resp_bits_pf ; 
    wire dcache_pma_checker_newEntry_gf = dcache_pma_checker_io_ptw_resp_bits_gf ; 
    wire dcache_pma_checker_newEntry_hr = dcache_pma_checker_io_ptw_resp_bits_hr ; 
    wire dcache_pma_checker_newEntry_hw = dcache_pma_checker_io_ptw_resp_bits_hw ; 
    wire dcache_pma_checker_newEntry_hx = dcache_pma_checker_io_ptw_resp_bits_hx ; 
    wire dcache_pma_checker_newEntry_u = dcache_pma_checker_io_ptw_resp_bits_pte_u ; 
    wire dcache_pma_checker_newEntry_fragmented_superpage = dcache_pma_checker_io_ptw_resp_bits_fragmented_superpage ; 
    wire[33:0] dcache_pma_checker_io_req_bits_vaddr ; 
    wire[20:0] dcache_pma_checker_vpn = dcache_pma_checker_io_req_bits_vaddr [32:12]; reg[1:0] dcache_pma_checker_sectored_entries_0_0_level ; reg[20:0] dcache_pma_checker_sectored_entries_0_0_tag_vpn ; 
    reg dcache_pma_checker_sectored_entries_0_0_tag_v ; reg[41:0] dcache_pma_checker_sectored_entries_0_0_data_0 ; reg[41:0] dcache_pma_checker_sectored_entries_0_0_data_1 ; reg[41:0] dcache_pma_checker_sectored_entries_0_0_data_2 ; reg[41:0] dcache_pma_checker_sectored_entries_0_0_data_3 ; 
    reg dcache_pma_checker_sectored_entries_0_0_valid_0 ; 
    reg dcache_pma_checker_sectored_entries_0_0_valid_1 ; 
    reg dcache_pma_checker_sectored_entries_0_0_valid_2 ; 
    reg dcache_pma_checker_sectored_entries_0_0_valid_3 ; reg[1:0] dcache_pma_checker_superpage_entries_0_level ; reg[20:0] dcache_pma_checker_superpage_entries_0_tag_vpn ; 
    reg dcache_pma_checker_superpage_entries_0_tag_v ; reg[41:0] dcache_pma_checker_superpage_entries_0_data_0 ; 
    wire[41:0] dcache_pma_checker__entries_WIRE_3 = dcache_pma_checker_superpage_entries_0_data_0 ; 
    reg dcache_pma_checker_superpage_entries_0_valid_0 ; reg[1:0] dcache_pma_checker_superpage_entries_1_level ; reg[20:0] dcache_pma_checker_superpage_entries_1_tag_vpn ; 
    reg dcache_pma_checker_superpage_entries_1_tag_v ; reg[41:0] dcache_pma_checker_superpage_entries_1_data_0 ; 
    wire[41:0] dcache_pma_checker__entries_WIRE_5 = dcache_pma_checker_superpage_entries_1_data_0 ; 
    reg dcache_pma_checker_superpage_entries_1_valid_0 ; reg[1:0] dcache_pma_checker_superpage_entries_2_level ; reg[20:0] dcache_pma_checker_superpage_entries_2_tag_vpn ; 
    reg dcache_pma_checker_superpage_entries_2_tag_v ; reg[41:0] dcache_pma_checker_superpage_entries_2_data_0 ; 
    wire[41:0] dcache_pma_checker__entries_WIRE_7 = dcache_pma_checker_superpage_entries_2_data_0 ; 
    reg dcache_pma_checker_superpage_entries_2_valid_0 ; reg[1:0] dcache_pma_checker_superpage_entries_3_level ; reg[20:0] dcache_pma_checker_superpage_entries_3_tag_vpn ; 
    reg dcache_pma_checker_superpage_entries_3_tag_v ; reg[41:0] dcache_pma_checker_superpage_entries_3_data_0 ; 
    wire[41:0] dcache_pma_checker__entries_WIRE_9 = dcache_pma_checker_superpage_entries_3_data_0 ; 
    reg dcache_pma_checker_superpage_entries_3_valid_0 ; reg[1:0] dcache_pma_checker_special_entry_level ; reg[20:0] dcache_pma_checker_special_entry_tag_vpn ; 
    reg dcache_pma_checker_special_entry_tag_v ; reg[41:0] dcache_pma_checker_special_entry_data_0 ; 
    wire[41:0] dcache_pma_checker__mpu_ppn_WIRE_1 = dcache_pma_checker_special_entry_data_0 ; 
    wire[41:0] dcache_pma_checker__entries_WIRE_11 = dcache_pma_checker_special_entry_data_0 ; 
    reg dcache_pma_checker_special_entry_valid_0 ; reg[1:0] dcache_pma_checker_state ; reg[20:0] dcache_pma_checker_r_refill_tag ; 
    wire[20:0] dcache_pma_checker_io_ptw_req_bits_bits_addr = dcache_pma_checker_r_refill_tag ; reg[1:0] dcache_pma_checker_r_superpage_repl_addr ; 
    wire[1:0] dcache_pma_checker_waddr = dcache_pma_checker_r_superpage_repl_addr ; 
    reg dcache_pma_checker_r_sectored_hit_valid ; 
    reg dcache_pma_checker_r_superpage_hit_valid ; reg[1:0] dcache_pma_checker_r_superpage_hit_bits ; 
    reg dcache_pma_checker_r_vstage1_en ; 
    wire dcache_pma_checker_io_ptw_req_bits_bits_vstage1 = dcache_pma_checker_r_vstage1_en ; 
    reg dcache_pma_checker_r_stage2_en ; 
    wire dcache_pma_checker_io_ptw_req_bits_bits_stage2 = dcache_pma_checker_r_stage2_en ; 
    reg dcache_pma_checker_r_need_gpa ; 
    wire dcache_pma_checker_io_ptw_req_bits_bits_need_gpa = dcache_pma_checker_r_need_gpa ; 
    reg dcache_pma_checker_r_gpa_valid ; reg[32:0] dcache_pma_checker_r_gpa ; reg[20:0] dcache_pma_checker_r_gpa_vpn ; 
    reg dcache_pma_checker_r_gpa_is_pte ; 
    wire[1:0] dcache_pma_checker_io_req_bits_prv ; 
    wire dcache_pma_checker_priv_s = dcache_pma_checker_io_req_bits_prv [0]; 
    wire dcache_pma_checker_priv_uses_vm = dcache_pma_checker_io_req_bits_prv <=2'h1; 
    wire[3:0] dcache_pma_checker_satp_mode = dcache_pma_checker_priv_v  ?  dcache_pma_checker_io_ptw_vsatp_mode : dcache_pma_checker_io_ptw_ptbr_mode ; 
    wire[15:0] dcache_pma_checker_satp_asid = dcache_pma_checker_priv_v  ?  dcache_pma_checker_io_ptw_vsatp_asid : dcache_pma_checker_io_ptw_ptbr_asid ; 
    wire[43:0] dcache_pma_checker_satp_ppn = dcache_pma_checker_priv_v  ?  dcache_pma_checker_io_ptw_vsatp_ppn : dcache_pma_checker_io_ptw_ptbr_ppn ; 
    wire dcache_pma_checker_vm_enabled =( dcache_pma_checker_stage1_en | dcache_pma_checker_stage2_en )& dcache_pma_checker_priv_uses_vm & dcache_pma_checker_io_req_bits_passthrough ==1'h0; 
    reg dcache_pma_checker_v_entries_use_stage1 ; 
    wire dcache_pma_checker_vsatp_mode_mismatch = dcache_pma_checker_priv_v & dcache_pma_checker_vstage1_en != dcache_pma_checker_v_entries_use_stage1 & dcache_pma_checker_io_req_bits_passthrough ==1'h0; 
    wire[19:0] dcache_pma_checker_refill_ppn = dcache_pma_checker_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire dcache_pma_checker_invalidate_refill = dcache_pma_checker_state ==2'h1|(& dcache_pma_checker_state )| dcache_pma_checker_io_sfence_valid ; 
    wire dcache_pma_checker__mpu_ppn_WIRE_fragmented_superpage = dcache_pma_checker__mpu_ppn_WIRE_1 [0]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_c = dcache_pma_checker__mpu_ppn_WIRE_1 [1]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_eff = dcache_pma_checker__mpu_ppn_WIRE_1 [2]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_paa = dcache_pma_checker__mpu_ppn_WIRE_1 [3]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_pal = dcache_pma_checker__mpu_ppn_WIRE_1 [4]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_ppp = dcache_pma_checker__mpu_ppn_WIRE_1 [5]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_pr = dcache_pma_checker__mpu_ppn_WIRE_1 [6]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_px = dcache_pma_checker__mpu_ppn_WIRE_1 [7]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_pw = dcache_pma_checker__mpu_ppn_WIRE_1 [8]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_hr = dcache_pma_checker__mpu_ppn_WIRE_1 [9]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_hx = dcache_pma_checker__mpu_ppn_WIRE_1 [10]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_hw = dcache_pma_checker__mpu_ppn_WIRE_1 [11]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_sr = dcache_pma_checker__mpu_ppn_WIRE_1 [12]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_sx = dcache_pma_checker__mpu_ppn_WIRE_1 [13]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_sw = dcache_pma_checker__mpu_ppn_WIRE_1 [14]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_gf = dcache_pma_checker__mpu_ppn_WIRE_1 [15]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_pf = dcache_pma_checker__mpu_ppn_WIRE_1 [16]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_ae_stage2 = dcache_pma_checker__mpu_ppn_WIRE_1 [17]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_ae_final = dcache_pma_checker__mpu_ppn_WIRE_1 [18]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_ae_ptw = dcache_pma_checker__mpu_ppn_WIRE_1 [19]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_g = dcache_pma_checker__mpu_ppn_WIRE_1 [20]; 
    wire dcache_pma_checker__mpu_ppn_WIRE_u = dcache_pma_checker__mpu_ppn_WIRE_1 [21]; 
    wire[19:0] dcache_pma_checker__mpu_ppn_WIRE_ppn = dcache_pma_checker__mpu_ppn_WIRE_1 [41:22];  
    
    assign  dcache_pma_checker_mpu_ppn_barrier_io_y_ppn = dcache_pma_checker_mpu_ppn_barrier_io_x_ppn ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_u = dcache_pma_checker_mpu_ppn_barrier_io_x_u ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_g = dcache_pma_checker_mpu_ppn_barrier_io_x_g ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_ae_ptw = dcache_pma_checker_mpu_ppn_barrier_io_x_ae_ptw ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_ae_final = dcache_pma_checker_mpu_ppn_barrier_io_x_ae_final ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_ae_stage2 = dcache_pma_checker_mpu_ppn_barrier_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_pf = dcache_pma_checker_mpu_ppn_barrier_io_x_pf ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_gf = dcache_pma_checker_mpu_ppn_barrier_io_x_gf ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_sw = dcache_pma_checker_mpu_ppn_barrier_io_x_sw ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_sx = dcache_pma_checker_mpu_ppn_barrier_io_x_sx ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_sr = dcache_pma_checker_mpu_ppn_barrier_io_x_sr ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_hw = dcache_pma_checker_mpu_ppn_barrier_io_x_hw ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_hx = dcache_pma_checker_mpu_ppn_barrier_io_x_hx ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_hr = dcache_pma_checker_mpu_ppn_barrier_io_x_hr ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_pw = dcache_pma_checker_mpu_ppn_barrier_io_x_pw ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_px = dcache_pma_checker_mpu_ppn_barrier_io_x_px ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_pr = dcache_pma_checker_mpu_ppn_barrier_io_x_pr ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_ppp = dcache_pma_checker_mpu_ppn_barrier_io_x_ppp ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_pal = dcache_pma_checker_mpu_ppn_barrier_io_x_pal ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_paa = dcache_pma_checker_mpu_ppn_barrier_io_x_paa ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_eff = dcache_pma_checker_mpu_ppn_barrier_io_x_eff ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_c = dcache_pma_checker_mpu_ppn_barrier_io_x_c ; 
  assign  dcache_pma_checker_mpu_ppn_barrier_io_y_fragmented_superpage = dcache_pma_checker_mpu_ppn_barrier_io_x_fragmented_superpage ;
     
    wire[21:0] dcache_pma_checker_mpu_ppn = dcache_pma_checker_do_refill  ? {2'h0, dcache_pma_checker_refill_ppn }: dcache_pma_checker_vm_enabled  ? {2'h0, dcache__pma_checker_mpu_ppn_barrier_io_y_ppn }: dcache_pma_checker_io_req_bits_vaddr [33:12]; 
    wire[33:0] dcache_pma_checker_mpu_physaddr ={ dcache_pma_checker_mpu_ppn , dcache_pma_checker_io_req_bits_vaddr [11:0]}; 
    wire[2:0] dcache_pma_checker_mpu_priv ={ dcache_pma_checker_io_ptw_status_debug , dcache_pma_checker_io_req_bits_prv }; 
    wire[1:0] dcache_pma_checker_io_req_bits_size ;  
    
    wire dcache_pma_checker_pmp_res_cur_cfg_l = dcache_pma_checker_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_cfg_res = dcache_pma_checker_pmp_io_pmp_7_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_cfg_a = dcache_pma_checker_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_addr = dcache_pma_checker_pmp_io_pmp_7_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_mask = dcache_pma_checker_pmp_io_pmp_7_mask ; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_l = dcache_pma_checker_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_1_cfg_res = dcache_pma_checker_pmp_io_pmp_6_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_1_cfg_a = dcache_pma_checker_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_1_addr = dcache_pma_checker_pmp_io_pmp_6_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_1_mask = dcache_pma_checker_pmp_io_pmp_6_mask ; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_l = dcache_pma_checker_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_2_cfg_res = dcache_pma_checker_pmp_io_pmp_5_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_2_cfg_a = dcache_pma_checker_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_2_addr = dcache_pma_checker_pmp_io_pmp_5_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_2_mask = dcache_pma_checker_pmp_io_pmp_5_mask ; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_l = dcache_pma_checker_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_3_cfg_res = dcache_pma_checker_pmp_io_pmp_4_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_3_cfg_a = dcache_pma_checker_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_3_addr = dcache_pma_checker_pmp_io_pmp_4_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_3_mask = dcache_pma_checker_pmp_io_pmp_4_mask ; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_l = dcache_pma_checker_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_4_cfg_res = dcache_pma_checker_pmp_io_pmp_3_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_4_cfg_a = dcache_pma_checker_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_4_addr = dcache_pma_checker_pmp_io_pmp_3_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_4_mask = dcache_pma_checker_pmp_io_pmp_3_mask ; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_l = dcache_pma_checker_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_5_cfg_res = dcache_pma_checker_pmp_io_pmp_2_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_5_cfg_a = dcache_pma_checker_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_5_addr = dcache_pma_checker_pmp_io_pmp_2_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_5_mask = dcache_pma_checker_pmp_io_pmp_2_mask ; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_l = dcache_pma_checker_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_6_cfg_res = dcache_pma_checker_pmp_io_pmp_1_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_6_cfg_a = dcache_pma_checker_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_6_addr = dcache_pma_checker_pmp_io_pmp_1_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_6_mask = dcache_pma_checker_pmp_io_pmp_1_mask ; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_l = dcache_pma_checker_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_7_cfg_res = dcache_pma_checker_pmp_io_pmp_0_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cur_7_cfg_a = dcache_pma_checker_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_res_cur_7_addr = dcache_pma_checker_pmp_io_pmp_0_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_cur_7_mask = dcache_pma_checker_pmp_io_pmp_0_mask ; 
    wire[1:0] dcache_pma_checker_pmp__pmp0_WIRE_cfg_res =2'h0; 
    wire[1:0] dcache_pma_checker_pmp__pmp0_WIRE_cfg_a =2'h0; 
    wire[29:0] dcache_pma_checker_pmp__pmp0_WIRE_addr =30'h0; 
    wire[31:0] dcache_pma_checker_pmp__pmp0_WIRE_mask =32'h0; 
    wire dcache_pma_checker_pmp__pmp0_WIRE_cfg_l =1'h0; 
    wire dcache_pma_checker_pmp__pmp0_WIRE_cfg_x =1'h0; 
    wire dcache_pma_checker_pmp__pmp0_WIRE_cfg_w =1'h0; 
    wire dcache_pma_checker_pmp__pmp0_WIRE_cfg_r =1'h0; 
    wire dcache_pma_checker_pmp_default_0 = dcache_pma_checker_pmp_io_prv >2'h1; 
    wire dcache_pma_checker_pmp_pmp0_cfg_x = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_pmp0_cfg_w = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_pmp0_cfg_r = dcache_pma_checker_pmp_default_0 ; 
    wire dcache_pma_checker_pmp_pmp0_cfg_l = dcache_pma_checker_pmp__pmp0_WIRE_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_pmp0_cfg_res = dcache_pma_checker_pmp__pmp0_WIRE_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_pmp0_cfg_a = dcache_pma_checker_pmp__pmp0_WIRE_cfg_a ; 
    wire[29:0] dcache_pma_checker_pmp_pmp0_addr = dcache_pma_checker_pmp__pmp0_WIRE_addr ; 
    wire[31:0] dcache_pma_checker_pmp_pmp0_mask = dcache_pma_checker_pmp__pmp0_WIRE_mask ; 
    wire[5:0] dcache_pma_checker_pmp__GEN =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask = dcache_pma_checker_pmp_io_pmp_7_mask |{29'h0,~( dcache_pma_checker_pmp__GEN [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_0 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_0 [31:3])&~( dcache_pma_checker_pmp_io_pmp_7_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_1 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_1 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_2 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_3 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_3 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_4 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_4 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_5 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_2 [2:0]))< dcache_pma_checker_pmp__GEN_5 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_6 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_1 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_6 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_7 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_1 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_7 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_8 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_1 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_8 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit = dcache_pma_checker_pmp_io_pmp_7_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch & dcache_pma_checker_pmp_res_hit_lsbMatch : dcache_pma_checker_pmp_io_pmp_7_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess | dcache_pma_checker_pmp_res_hit_msbsEqual & dcache_pma_checker_pmp_res_hit_lsbsLess )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_1 | dcache_pma_checker_pmp_res_hit_msbsEqual_1 & dcache_pma_checker_pmp_res_hit_lsbsLess_1 ); 
    wire dcache_pma_checker_pmp_res_ignore = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_7_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_9 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask =~( dcache_pma_checker_pmp__GEN_9 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_10 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_11 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_10 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_11 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_12 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_13 =~(~{ dcache_pma_checker_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_12 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_13 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned =( dcache_pma_checker_pmp_res_aligned_lsbMask &~( dcache_pma_checker_pmp_io_pmp_7_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned = dcache_pma_checker_pmp_io_pmp_7_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned : dcache_pma_checker_pmp_res_aligned_rangeAligned ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_1 ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_2 ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_3 ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_4 ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_5 ={ dcache_pma_checker_pmp_io_pmp_7_cfg_x , dcache_pma_checker_pmp_io_pmp_7_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_cfg_r = dcache_pma_checker_pmp_res_aligned &( dcache_pma_checker_pmp_io_pmp_7_cfg_r | dcache_pma_checker_pmp_res_ignore ); 
    wire dcache_pma_checker_pmp_res_cur_cfg_w = dcache_pma_checker_pmp_res_aligned &( dcache_pma_checker_pmp_io_pmp_7_cfg_w | dcache_pma_checker_pmp_res_ignore ); 
    wire dcache_pma_checker_pmp_res_cur_cfg_x = dcache_pma_checker_pmp_res_aligned &( dcache_pma_checker_pmp_io_pmp_7_cfg_x | dcache_pma_checker_pmp_res_ignore ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_14 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_1 = dcache_pma_checker_pmp_io_pmp_6_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_14 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_15 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_1 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_15 [31:3])&~( dcache_pma_checker_pmp_io_pmp_6_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_16 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_1 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_16 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_1 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_17 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_18 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_2 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_18 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_19 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_2 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_19 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_20 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_2 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_17 [2:0]))< dcache_pma_checker_pmp__GEN_20 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_21 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_3 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_21 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_22 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_3 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_22 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_23 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_3 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_23 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_1 = dcache_pma_checker_pmp_io_pmp_6_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_1 & dcache_pma_checker_pmp_res_hit_lsbMatch_1 : dcache_pma_checker_pmp_io_pmp_6_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_2 | dcache_pma_checker_pmp_res_hit_msbsEqual_2 & dcache_pma_checker_pmp_res_hit_lsbsLess_2 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_3 | dcache_pma_checker_pmp_res_hit_msbsEqual_3 & dcache_pma_checker_pmp_res_hit_lsbsLess_3 ); 
    wire dcache_pma_checker_pmp_res_ignore_1 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_6_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_24 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_1 =~( dcache_pma_checker_pmp__GEN_24 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_25 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_26 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_1 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_25 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_26 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_27 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_28 =~(~{ dcache_pma_checker_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_1 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_27 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_28 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_1 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_1 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_1 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_1 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_1 =( dcache_pma_checker_pmp_res_aligned_lsbMask_1 &~( dcache_pma_checker_pmp_io_pmp_6_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_1 = dcache_pma_checker_pmp_io_pmp_6_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_1 : dcache_pma_checker_pmp_res_aligned_rangeAligned_1 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_6 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_7 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_8 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_9 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_10 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_11 ={ dcache_pma_checker_pmp_io_pmp_6_cfg_x , dcache_pma_checker_pmp_io_pmp_6_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_r = dcache_pma_checker_pmp_res_aligned_1 &( dcache_pma_checker_pmp_io_pmp_6_cfg_r | dcache_pma_checker_pmp_res_ignore_1 ); 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_w = dcache_pma_checker_pmp_res_aligned_1 &( dcache_pma_checker_pmp_io_pmp_6_cfg_w | dcache_pma_checker_pmp_res_ignore_1 ); 
    wire dcache_pma_checker_pmp_res_cur_1_cfg_x = dcache_pma_checker_pmp_res_aligned_1 &( dcache_pma_checker_pmp_io_pmp_6_cfg_x | dcache_pma_checker_pmp_res_ignore_1 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_29 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_2 = dcache_pma_checker_pmp_io_pmp_5_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_29 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_30 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_2 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_30 [31:3])&~( dcache_pma_checker_pmp_io_pmp_5_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_31 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_2 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_31 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_2 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_32 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_33 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_4 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_33 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_34 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_4 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_34 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_35 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_4 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_32 [2:0]))< dcache_pma_checker_pmp__GEN_35 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_36 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_5 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_36 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_37 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_5 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_37 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_38 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_5 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_38 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_2 = dcache_pma_checker_pmp_io_pmp_5_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_2 & dcache_pma_checker_pmp_res_hit_lsbMatch_2 : dcache_pma_checker_pmp_io_pmp_5_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_4 | dcache_pma_checker_pmp_res_hit_msbsEqual_4 & dcache_pma_checker_pmp_res_hit_lsbsLess_4 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_5 | dcache_pma_checker_pmp_res_hit_msbsEqual_5 & dcache_pma_checker_pmp_res_hit_lsbsLess_5 ); 
    wire dcache_pma_checker_pmp_res_ignore_2 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_5_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_39 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_2 =~( dcache_pma_checker_pmp__GEN_39 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_40 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_41 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_2 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_40 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_41 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_42 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_43 =~(~{ dcache_pma_checker_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_2 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_42 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_43 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_2 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_2 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_2 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_2 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_2 =( dcache_pma_checker_pmp_res_aligned_lsbMask_2 &~( dcache_pma_checker_pmp_io_pmp_5_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_2 = dcache_pma_checker_pmp_io_pmp_5_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_2 : dcache_pma_checker_pmp_res_aligned_rangeAligned_2 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_12 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_13 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_14 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_15 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_16 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_17 ={ dcache_pma_checker_pmp_io_pmp_5_cfg_x , dcache_pma_checker_pmp_io_pmp_5_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_r = dcache_pma_checker_pmp_res_aligned_2 &( dcache_pma_checker_pmp_io_pmp_5_cfg_r | dcache_pma_checker_pmp_res_ignore_2 ); 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_w = dcache_pma_checker_pmp_res_aligned_2 &( dcache_pma_checker_pmp_io_pmp_5_cfg_w | dcache_pma_checker_pmp_res_ignore_2 ); 
    wire dcache_pma_checker_pmp_res_cur_2_cfg_x = dcache_pma_checker_pmp_res_aligned_2 &( dcache_pma_checker_pmp_io_pmp_5_cfg_x | dcache_pma_checker_pmp_res_ignore_2 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_44 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_3 = dcache_pma_checker_pmp_io_pmp_4_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_44 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_45 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_3 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_45 [31:3])&~( dcache_pma_checker_pmp_io_pmp_4_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_46 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_3 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_46 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_3 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_47 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_48 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_6 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_48 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_49 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_6 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_49 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_50 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_6 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_47 [2:0]))< dcache_pma_checker_pmp__GEN_50 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_51 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_7 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_51 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_52 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_7 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_52 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_53 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_7 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_53 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_3 = dcache_pma_checker_pmp_io_pmp_4_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_3 & dcache_pma_checker_pmp_res_hit_lsbMatch_3 : dcache_pma_checker_pmp_io_pmp_4_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_6 | dcache_pma_checker_pmp_res_hit_msbsEqual_6 & dcache_pma_checker_pmp_res_hit_lsbsLess_6 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_7 | dcache_pma_checker_pmp_res_hit_msbsEqual_7 & dcache_pma_checker_pmp_res_hit_lsbsLess_7 ); 
    wire dcache_pma_checker_pmp_res_ignore_3 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_4_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_54 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_3 =~( dcache_pma_checker_pmp__GEN_54 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_55 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_56 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_3 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_55 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_56 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_57 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_58 =~(~{ dcache_pma_checker_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_3 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_57 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_58 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_3 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_3 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_3 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_3 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_3 =( dcache_pma_checker_pmp_res_aligned_lsbMask_3 &~( dcache_pma_checker_pmp_io_pmp_4_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_3 = dcache_pma_checker_pmp_io_pmp_4_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_3 : dcache_pma_checker_pmp_res_aligned_rangeAligned_3 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_18 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_19 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_20 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_21 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_22 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_23 ={ dcache_pma_checker_pmp_io_pmp_4_cfg_x , dcache_pma_checker_pmp_io_pmp_4_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_r = dcache_pma_checker_pmp_res_aligned_3 &( dcache_pma_checker_pmp_io_pmp_4_cfg_r | dcache_pma_checker_pmp_res_ignore_3 ); 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_w = dcache_pma_checker_pmp_res_aligned_3 &( dcache_pma_checker_pmp_io_pmp_4_cfg_w | dcache_pma_checker_pmp_res_ignore_3 ); 
    wire dcache_pma_checker_pmp_res_cur_3_cfg_x = dcache_pma_checker_pmp_res_aligned_3 &( dcache_pma_checker_pmp_io_pmp_4_cfg_x | dcache_pma_checker_pmp_res_ignore_3 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_59 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_4 = dcache_pma_checker_pmp_io_pmp_3_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_59 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_60 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_4 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_60 [31:3])&~( dcache_pma_checker_pmp_io_pmp_3_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_61 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_4 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_61 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_4 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_62 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_63 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_8 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_63 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_64 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_8 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_64 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_65 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_8 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_62 [2:0]))< dcache_pma_checker_pmp__GEN_65 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_66 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_9 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_66 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_67 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_9 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_67 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_68 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_9 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_68 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_4 = dcache_pma_checker_pmp_io_pmp_3_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_4 & dcache_pma_checker_pmp_res_hit_lsbMatch_4 : dcache_pma_checker_pmp_io_pmp_3_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_8 | dcache_pma_checker_pmp_res_hit_msbsEqual_8 & dcache_pma_checker_pmp_res_hit_lsbsLess_8 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_9 | dcache_pma_checker_pmp_res_hit_msbsEqual_9 & dcache_pma_checker_pmp_res_hit_lsbsLess_9 ); 
    wire dcache_pma_checker_pmp_res_ignore_4 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_3_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_69 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_4 =~( dcache_pma_checker_pmp__GEN_69 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_70 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_71 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_4 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_70 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_71 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_72 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_73 =~(~{ dcache_pma_checker_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_4 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_72 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_73 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_4 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_4 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_4 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_4 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_4 =( dcache_pma_checker_pmp_res_aligned_lsbMask_4 &~( dcache_pma_checker_pmp_io_pmp_3_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_4 = dcache_pma_checker_pmp_io_pmp_3_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_4 : dcache_pma_checker_pmp_res_aligned_rangeAligned_4 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_24 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_25 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_26 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_27 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_28 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_29 ={ dcache_pma_checker_pmp_io_pmp_3_cfg_x , dcache_pma_checker_pmp_io_pmp_3_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_r = dcache_pma_checker_pmp_res_aligned_4 &( dcache_pma_checker_pmp_io_pmp_3_cfg_r | dcache_pma_checker_pmp_res_ignore_4 ); 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_w = dcache_pma_checker_pmp_res_aligned_4 &( dcache_pma_checker_pmp_io_pmp_3_cfg_w | dcache_pma_checker_pmp_res_ignore_4 ); 
    wire dcache_pma_checker_pmp_res_cur_4_cfg_x = dcache_pma_checker_pmp_res_aligned_4 &( dcache_pma_checker_pmp_io_pmp_3_cfg_x | dcache_pma_checker_pmp_res_ignore_4 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_74 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_5 = dcache_pma_checker_pmp_io_pmp_2_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_74 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_75 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_5 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_75 [31:3])&~( dcache_pma_checker_pmp_io_pmp_2_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_76 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_5 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_76 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_5 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_77 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_78 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_10 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_78 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_79 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_10 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_79 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_80 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_10 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_77 [2:0]))< dcache_pma_checker_pmp__GEN_80 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_81 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_11 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_81 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_82 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_11 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_82 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_83 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_11 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_83 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_5 = dcache_pma_checker_pmp_io_pmp_2_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_5 & dcache_pma_checker_pmp_res_hit_lsbMatch_5 : dcache_pma_checker_pmp_io_pmp_2_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_10 | dcache_pma_checker_pmp_res_hit_msbsEqual_10 & dcache_pma_checker_pmp_res_hit_lsbsLess_10 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_11 | dcache_pma_checker_pmp_res_hit_msbsEqual_11 & dcache_pma_checker_pmp_res_hit_lsbsLess_11 ); 
    wire dcache_pma_checker_pmp_res_ignore_5 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_2_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_84 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_5 =~( dcache_pma_checker_pmp__GEN_84 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_85 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_86 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_5 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_85 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_86 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_87 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_88 =~(~{ dcache_pma_checker_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_5 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_87 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_88 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_5 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_5 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_5 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_5 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_5 =( dcache_pma_checker_pmp_res_aligned_lsbMask_5 &~( dcache_pma_checker_pmp_io_pmp_2_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_5 = dcache_pma_checker_pmp_io_pmp_2_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_5 : dcache_pma_checker_pmp_res_aligned_rangeAligned_5 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_30 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_31 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_32 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_33 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_34 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_35 ={ dcache_pma_checker_pmp_io_pmp_2_cfg_x , dcache_pma_checker_pmp_io_pmp_2_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_r = dcache_pma_checker_pmp_res_aligned_5 &( dcache_pma_checker_pmp_io_pmp_2_cfg_r | dcache_pma_checker_pmp_res_ignore_5 ); 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_w = dcache_pma_checker_pmp_res_aligned_5 &( dcache_pma_checker_pmp_io_pmp_2_cfg_w | dcache_pma_checker_pmp_res_ignore_5 ); 
    wire dcache_pma_checker_pmp_res_cur_5_cfg_x = dcache_pma_checker_pmp_res_aligned_5 &( dcache_pma_checker_pmp_io_pmp_2_cfg_x | dcache_pma_checker_pmp_res_ignore_5 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_89 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_6 = dcache_pma_checker_pmp_io_pmp_1_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_89 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_90 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_6 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_90 [31:3])&~( dcache_pma_checker_pmp_io_pmp_1_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_91 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_6 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_91 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_6 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_92 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_93 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_12 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_93 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_94 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_12 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_94 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_95 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_12 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_92 [2:0]))< dcache_pma_checker_pmp__GEN_95 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_96 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_13 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_96 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_97 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_13 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_97 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_98 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_13 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_98 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_6 = dcache_pma_checker_pmp_io_pmp_1_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_6 & dcache_pma_checker_pmp_res_hit_lsbMatch_6 : dcache_pma_checker_pmp_io_pmp_1_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_12 | dcache_pma_checker_pmp_res_hit_msbsEqual_12 & dcache_pma_checker_pmp_res_hit_lsbsLess_12 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_13 | dcache_pma_checker_pmp_res_hit_msbsEqual_13 & dcache_pma_checker_pmp_res_hit_lsbsLess_13 ); 
    wire dcache_pma_checker_pmp_res_ignore_6 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_1_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_99 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_6 =~( dcache_pma_checker_pmp__GEN_99 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_100 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_101 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_6 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_100 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_101 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_102 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_103 =~(~{ dcache_pma_checker_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_6 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_102 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_103 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_6 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_6 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_6 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_6 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_6 =( dcache_pma_checker_pmp_res_aligned_lsbMask_6 &~( dcache_pma_checker_pmp_io_pmp_1_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_6 = dcache_pma_checker_pmp_io_pmp_1_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_6 : dcache_pma_checker_pmp_res_aligned_rangeAligned_6 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_36 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_37 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_38 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_39 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_40 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_41 ={ dcache_pma_checker_pmp_io_pmp_1_cfg_x , dcache_pma_checker_pmp_io_pmp_1_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_r = dcache_pma_checker_pmp_res_aligned_6 &( dcache_pma_checker_pmp_io_pmp_1_cfg_r | dcache_pma_checker_pmp_res_ignore_6 ); 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_w = dcache_pma_checker_pmp_res_aligned_6 &( dcache_pma_checker_pmp_io_pmp_1_cfg_w | dcache_pma_checker_pmp_res_ignore_6 ); 
    wire dcache_pma_checker_pmp_res_cur_6_cfg_x = dcache_pma_checker_pmp_res_aligned_6 &( dcache_pma_checker_pmp_io_pmp_1_cfg_x | dcache_pma_checker_pmp_res_ignore_6 ); 
    wire[5:0] dcache_pma_checker_pmp__GEN_104 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp_res_hit_lsbMask_7 = dcache_pma_checker_pmp_io_pmp_0_mask |{29'h0,~( dcache_pma_checker_pmp__GEN_104 [2:0])}; 
    wire[31:0] dcache_pma_checker_pmp__GEN_105 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbMatch_7 =(( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_105 [31:3])&~( dcache_pma_checker_pmp_io_pmp_0_mask [31:3]))==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_106 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbMatch_7 =(( dcache_pma_checker_pmp_io_addr [2:0]^ dcache_pma_checker_pmp__GEN_106 [2:0])&~( dcache_pma_checker_pmp_res_hit_lsbMask_7 [2:0]))==3'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_107 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[31:0] dcache_pma_checker_pmp__GEN_108 =~(~{ dcache_pma_checker_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_14 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_108 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_109 =~(~{ dcache_pma_checker_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_14 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_109 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_110 =~(~{ dcache_pma_checker_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_14 =( dcache_pma_checker_pmp_io_addr [2:0]|~( dcache_pma_checker_pmp__GEN_107 [2:0]))< dcache_pma_checker_pmp__GEN_110 [2:0]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_111 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsLess_15 = dcache_pma_checker_pmp_io_addr [31:3]< dcache_pma_checker_pmp__GEN_111 [31:3]; 
    wire[31:0] dcache_pma_checker_pmp__GEN_112 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_msbsEqual_15 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_112 [31:3])==29'h0; 
    wire[31:0] dcache_pma_checker_pmp__GEN_113 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_hit_lsbsLess_15 = dcache_pma_checker_pmp_io_addr [2:0]< dcache_pma_checker_pmp__GEN_113 [2:0]; 
    wire dcache_pma_checker_pmp_res_hit_7 = dcache_pma_checker_pmp_io_pmp_0_cfg_a [1] ?  dcache_pma_checker_pmp_res_hit_msbMatch_7 & dcache_pma_checker_pmp_res_hit_lsbMatch_7 : dcache_pma_checker_pmp_io_pmp_0_cfg_a [0]&( dcache_pma_checker_pmp_res_hit_msbsLess_14 | dcache_pma_checker_pmp_res_hit_msbsEqual_14 & dcache_pma_checker_pmp_res_hit_lsbsLess_14 )==1'h0&( dcache_pma_checker_pmp_res_hit_msbsLess_15 | dcache_pma_checker_pmp_res_hit_msbsEqual_15 & dcache_pma_checker_pmp_res_hit_lsbsLess_15 ); 
    wire dcache_pma_checker_pmp_res_ignore_7 = dcache_pma_checker_pmp_default_0 & dcache_pma_checker_pmp_io_pmp_0_cfg_l ==1'h0; 
    wire[5:0] dcache_pma_checker_pmp__GEN_114 =6'h7<< dcache_pma_checker_pmp_io_size ; 
    wire[2:0] dcache_pma_checker_pmp_res_aligned_lsbMask_7 =~( dcache_pma_checker_pmp__GEN_114 [2:0]); 
    wire[31:0] dcache_pma_checker_pmp__GEN_115 =~(~{ dcache_pma_checker_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_116 =~(~{ dcache_pma_checker_pmp_pmp0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_7 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_115 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_116 [2:0]&~( dcache_pma_checker_pmp_io_addr [2:0]))); 
    wire[31:0] dcache_pma_checker_pmp__GEN_117 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire[31:0] dcache_pma_checker_pmp__GEN_118 =~(~{ dcache_pma_checker_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_7 =( dcache_pma_checker_pmp_io_addr [31:3]^ dcache_pma_checker_pmp__GEN_117 [31:3])==29'h0&(|( dcache_pma_checker_pmp__GEN_118 [2:0]&( dcache_pma_checker_pmp_io_addr [2:0]| dcache_pma_checker_pmp_res_aligned_lsbMask_7 ))); 
    wire dcache_pma_checker_pmp_res_aligned_rangeAligned_7 =( dcache_pma_checker_pmp_res_aligned_straddlesLowerBound_7 | dcache_pma_checker_pmp_res_aligned_straddlesUpperBound_7 )==1'h0; 
    wire dcache_pma_checker_pmp_res_aligned_pow2Aligned_7 =( dcache_pma_checker_pmp_res_aligned_lsbMask_7 &~( dcache_pma_checker_pmp_io_pmp_0_mask [2:0]))==3'h0; 
    wire dcache_pma_checker_pmp_res_aligned_7 = dcache_pma_checker_pmp_io_pmp_0_cfg_a [1] ?  dcache_pma_checker_pmp_res_aligned_pow2Aligned_7 : dcache_pma_checker_pmp_res_aligned_rangeAligned_7 ; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_42 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_43 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_44 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_45 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_46 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] dcache_pma_checker_pmp_res_hi_47 ={ dcache_pma_checker_pmp_io_pmp_0_cfg_x , dcache_pma_checker_pmp_io_pmp_0_cfg_w }; 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_r = dcache_pma_checker_pmp_res_aligned_7 &( dcache_pma_checker_pmp_io_pmp_0_cfg_r | dcache_pma_checker_pmp_res_ignore_7 ); 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_w = dcache_pma_checker_pmp_res_aligned_7 &( dcache_pma_checker_pmp_io_pmp_0_cfg_w | dcache_pma_checker_pmp_res_ignore_7 ); 
    wire dcache_pma_checker_pmp_res_cur_7_cfg_x = dcache_pma_checker_pmp_res_aligned_7 &( dcache_pma_checker_pmp_io_pmp_0_cfg_x | dcache_pma_checker_pmp_res_ignore_7 ); 
    wire dcache_pma_checker_pmp_res_cfg_l = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_l : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_l : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_l : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_l : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_l : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_l : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_l : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_l : dcache_pma_checker_pmp_pmp0_cfg_l ; 
    wire[1:0] dcache_pma_checker_pmp_res_cfg_res = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_res : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_res : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_res : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_res : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_res : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_res : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_res : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_res : dcache_pma_checker_pmp_pmp0_cfg_res ; 
    wire[1:0] dcache_pma_checker_pmp_res_cfg_a = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_a : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_a : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_a : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_a : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_a : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_a : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_a : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_a : dcache_pma_checker_pmp_pmp0_cfg_a ; 
    wire dcache_pma_checker_pmp_res_cfg_x = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_x : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_x : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_x : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_x : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_x : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_x : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_x : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_x : dcache_pma_checker_pmp_pmp0_cfg_x ; 
    wire dcache_pma_checker_pmp_res_cfg_w = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_w : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_w : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_w : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_w : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_w : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_w : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_w : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_w : dcache_pma_checker_pmp_pmp0_cfg_w ; 
    wire dcache_pma_checker_pmp_res_cfg_r = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_cfg_r : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_cfg_r : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_cfg_r : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_cfg_r : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_cfg_r : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_cfg_r : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_cfg_r : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_cfg_r : dcache_pma_checker_pmp_pmp0_cfg_r ; 
    wire[29:0] dcache_pma_checker_pmp_res_addr = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_addr : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_addr : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_addr : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_addr : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_addr : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_addr : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_addr : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_addr : dcache_pma_checker_pmp_pmp0_addr ; 
    wire[31:0] dcache_pma_checker_pmp_res_mask = dcache_pma_checker_pmp_res_hit_7  ?  dcache_pma_checker_pmp_res_cur_7_mask : dcache_pma_checker_pmp_res_hit_6  ?  dcache_pma_checker_pmp_res_cur_6_mask : dcache_pma_checker_pmp_res_hit_5  ?  dcache_pma_checker_pmp_res_cur_5_mask : dcache_pma_checker_pmp_res_hit_4  ?  dcache_pma_checker_pmp_res_cur_4_mask : dcache_pma_checker_pmp_res_hit_3  ?  dcache_pma_checker_pmp_res_cur_3_mask : dcache_pma_checker_pmp_res_hit_2  ?  dcache_pma_checker_pmp_res_cur_2_mask : dcache_pma_checker_pmp_res_hit_1  ?  dcache_pma_checker_pmp_res_cur_1_mask : dcache_pma_checker_pmp_res_hit  ?  dcache_pma_checker_pmp_res_cur_mask : dcache_pma_checker_pmp_pmp0_mask ; 
  assign  dcache_pma_checker_pmp_io_r = dcache_pma_checker_pmp_res_cfg_r ; 
  assign  dcache_pma_checker_pmp_io_w = dcache_pma_checker_pmp_res_cfg_w ; 
  assign  dcache_pma_checker_pmp_io_x = dcache_pma_checker_pmp_res_cfg_x ;
    assign dcache_tlb_pmp_clock = dcache_tlb_clock;
    assign dcache_tlb_pmp_reset = dcache_tlb_reset;
    assign dcache_tlb_pmp_io_prv = dcache__tlb_mpu_priv_1to0;
    assign dcache_tlb_pmp_io_pmp_0_cfg_l = dcache_tlb_io_ptw_pmp_0_cfg_l;
    assign dcache_tlb_pmp_io_pmp_0_cfg_res = dcache_tlb_io_ptw_pmp_0_cfg_res;
    assign dcache_tlb_pmp_io_pmp_0_cfg_a = dcache_tlb_io_ptw_pmp_0_cfg_a;
    assign dcache_tlb_pmp_io_pmp_0_cfg_x = dcache_tlb_io_ptw_pmp_0_cfg_x;
    assign dcache_tlb_pmp_io_pmp_0_cfg_w = dcache_tlb_io_ptw_pmp_0_cfg_w;
    assign dcache_tlb_pmp_io_pmp_0_cfg_r = dcache_tlb_io_ptw_pmp_0_cfg_r;
    assign dcache_tlb_pmp_io_pmp_0_addr = dcache_tlb_io_ptw_pmp_0_addr;
    assign dcache_tlb_pmp_io_pmp_0_mask = dcache_tlb_io_ptw_pmp_0_mask;
    assign dcache_tlb_pmp_io_pmp_1_cfg_l = dcache_tlb_io_ptw_pmp_1_cfg_l;
    assign dcache_tlb_pmp_io_pmp_1_cfg_res = dcache_tlb_io_ptw_pmp_1_cfg_res;
    assign dcache_tlb_pmp_io_pmp_1_cfg_a = dcache_tlb_io_ptw_pmp_1_cfg_a;
    assign dcache_tlb_pmp_io_pmp_1_cfg_x = dcache_tlb_io_ptw_pmp_1_cfg_x;
    assign dcache_tlb_pmp_io_pmp_1_cfg_w = dcache_tlb_io_ptw_pmp_1_cfg_w;
    assign dcache_tlb_pmp_io_pmp_1_cfg_r = dcache_tlb_io_ptw_pmp_1_cfg_r;
    assign dcache_tlb_pmp_io_pmp_1_addr = dcache_tlb_io_ptw_pmp_1_addr;
    assign dcache_tlb_pmp_io_pmp_1_mask = dcache_tlb_io_ptw_pmp_1_mask;
    assign dcache_tlb_pmp_io_pmp_2_cfg_l = dcache_tlb_io_ptw_pmp_2_cfg_l;
    assign dcache_tlb_pmp_io_pmp_2_cfg_res = dcache_tlb_io_ptw_pmp_2_cfg_res;
    assign dcache_tlb_pmp_io_pmp_2_cfg_a = dcache_tlb_io_ptw_pmp_2_cfg_a;
    assign dcache_tlb_pmp_io_pmp_2_cfg_x = dcache_tlb_io_ptw_pmp_2_cfg_x;
    assign dcache_tlb_pmp_io_pmp_2_cfg_w = dcache_tlb_io_ptw_pmp_2_cfg_w;
    assign dcache_tlb_pmp_io_pmp_2_cfg_r = dcache_tlb_io_ptw_pmp_2_cfg_r;
    assign dcache_tlb_pmp_io_pmp_2_addr = dcache_tlb_io_ptw_pmp_2_addr;
    assign dcache_tlb_pmp_io_pmp_2_mask = dcache_tlb_io_ptw_pmp_2_mask;
    assign dcache_tlb_pmp_io_pmp_3_cfg_l = dcache_tlb_io_ptw_pmp_3_cfg_l;
    assign dcache_tlb_pmp_io_pmp_3_cfg_res = dcache_tlb_io_ptw_pmp_3_cfg_res;
    assign dcache_tlb_pmp_io_pmp_3_cfg_a = dcache_tlb_io_ptw_pmp_3_cfg_a;
    assign dcache_tlb_pmp_io_pmp_3_cfg_x = dcache_tlb_io_ptw_pmp_3_cfg_x;
    assign dcache_tlb_pmp_io_pmp_3_cfg_w = dcache_tlb_io_ptw_pmp_3_cfg_w;
    assign dcache_tlb_pmp_io_pmp_3_cfg_r = dcache_tlb_io_ptw_pmp_3_cfg_r;
    assign dcache_tlb_pmp_io_pmp_3_addr = dcache_tlb_io_ptw_pmp_3_addr;
    assign dcache_tlb_pmp_io_pmp_3_mask = dcache_tlb_io_ptw_pmp_3_mask;
    assign dcache_tlb_pmp_io_pmp_4_cfg_l = dcache_tlb_io_ptw_pmp_4_cfg_l;
    assign dcache_tlb_pmp_io_pmp_4_cfg_res = dcache_tlb_io_ptw_pmp_4_cfg_res;
    assign dcache_tlb_pmp_io_pmp_4_cfg_a = dcache_tlb_io_ptw_pmp_4_cfg_a;
    assign dcache_tlb_pmp_io_pmp_4_cfg_x = dcache_tlb_io_ptw_pmp_4_cfg_x;
    assign dcache_tlb_pmp_io_pmp_4_cfg_w = dcache_tlb_io_ptw_pmp_4_cfg_w;
    assign dcache_tlb_pmp_io_pmp_4_cfg_r = dcache_tlb_io_ptw_pmp_4_cfg_r;
    assign dcache_tlb_pmp_io_pmp_4_addr = dcache_tlb_io_ptw_pmp_4_addr;
    assign dcache_tlb_pmp_io_pmp_4_mask = dcache_tlb_io_ptw_pmp_4_mask;
    assign dcache_tlb_pmp_io_pmp_5_cfg_l = dcache_tlb_io_ptw_pmp_5_cfg_l;
    assign dcache_tlb_pmp_io_pmp_5_cfg_res = dcache_tlb_io_ptw_pmp_5_cfg_res;
    assign dcache_tlb_pmp_io_pmp_5_cfg_a = dcache_tlb_io_ptw_pmp_5_cfg_a;
    assign dcache_tlb_pmp_io_pmp_5_cfg_x = dcache_tlb_io_ptw_pmp_5_cfg_x;
    assign dcache_tlb_pmp_io_pmp_5_cfg_w = dcache_tlb_io_ptw_pmp_5_cfg_w;
    assign dcache_tlb_pmp_io_pmp_5_cfg_r = dcache_tlb_io_ptw_pmp_5_cfg_r;
    assign dcache_tlb_pmp_io_pmp_5_addr = dcache_tlb_io_ptw_pmp_5_addr;
    assign dcache_tlb_pmp_io_pmp_5_mask = dcache_tlb_io_ptw_pmp_5_mask;
    assign dcache_tlb_pmp_io_pmp_6_cfg_l = dcache_tlb_io_ptw_pmp_6_cfg_l;
    assign dcache_tlb_pmp_io_pmp_6_cfg_res = dcache_tlb_io_ptw_pmp_6_cfg_res;
    assign dcache_tlb_pmp_io_pmp_6_cfg_a = dcache_tlb_io_ptw_pmp_6_cfg_a;
    assign dcache_tlb_pmp_io_pmp_6_cfg_x = dcache_tlb_io_ptw_pmp_6_cfg_x;
    assign dcache_tlb_pmp_io_pmp_6_cfg_w = dcache_tlb_io_ptw_pmp_6_cfg_w;
    assign dcache_tlb_pmp_io_pmp_6_cfg_r = dcache_tlb_io_ptw_pmp_6_cfg_r;
    assign dcache_tlb_pmp_io_pmp_6_addr = dcache_tlb_io_ptw_pmp_6_addr;
    assign dcache_tlb_pmp_io_pmp_6_mask = dcache_tlb_io_ptw_pmp_6_mask;
    assign dcache_tlb_pmp_io_pmp_7_cfg_l = dcache_tlb_io_ptw_pmp_7_cfg_l;
    assign dcache_tlb_pmp_io_pmp_7_cfg_res = dcache_tlb_io_ptw_pmp_7_cfg_res;
    assign dcache_tlb_pmp_io_pmp_7_cfg_a = dcache_tlb_io_ptw_pmp_7_cfg_a;
    assign dcache_tlb_pmp_io_pmp_7_cfg_x = dcache_tlb_io_ptw_pmp_7_cfg_x;
    assign dcache_tlb_pmp_io_pmp_7_cfg_w = dcache_tlb_io_ptw_pmp_7_cfg_w;
    assign dcache_tlb_pmp_io_pmp_7_cfg_r = dcache_tlb_io_ptw_pmp_7_cfg_r;
    assign dcache_tlb_pmp_io_pmp_7_addr = dcache_tlb_io_ptw_pmp_7_addr;
    assign dcache_tlb_pmp_io_pmp_7_mask = dcache_tlb_io_ptw_pmp_7_mask;
    assign dcache_tlb_pmp_io_addr = dcache__tlb_mpu_physaddr_31to0;
    assign dcache_tlb_pmp_io_size = dcache_tlb_io_req_bits_size;
    assign dcache__tlb_pmp_io_r = dcache_tlb_pmp_io_r;
    assign dcache__tlb_pmp_io_w = dcache_tlb_pmp_io_w;
    assign dcache__tlb_pmp_io_x = dcache_tlb_pmp_io_x;
    assign dcache_pma_checker_pmp_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_pmp_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_pmp_io_prv = dcache__pma_checker_mpu_priv_1to0;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_l = dcache_pma_checker_io_ptw_pmp_0_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_res = dcache_pma_checker_io_ptw_pmp_0_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_a = dcache_pma_checker_io_ptw_pmp_0_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_x = dcache_pma_checker_io_ptw_pmp_0_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_w = dcache_pma_checker_io_ptw_pmp_0_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_0_cfg_r = dcache_pma_checker_io_ptw_pmp_0_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_0_addr = dcache_pma_checker_io_ptw_pmp_0_addr;
    assign dcache_pma_checker_pmp_io_pmp_0_mask = dcache_pma_checker_io_ptw_pmp_0_mask;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_l = dcache_pma_checker_io_ptw_pmp_1_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_res = dcache_pma_checker_io_ptw_pmp_1_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_a = dcache_pma_checker_io_ptw_pmp_1_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_x = dcache_pma_checker_io_ptw_pmp_1_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_w = dcache_pma_checker_io_ptw_pmp_1_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_1_cfg_r = dcache_pma_checker_io_ptw_pmp_1_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_1_addr = dcache_pma_checker_io_ptw_pmp_1_addr;
    assign dcache_pma_checker_pmp_io_pmp_1_mask = dcache_pma_checker_io_ptw_pmp_1_mask;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_l = dcache_pma_checker_io_ptw_pmp_2_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_res = dcache_pma_checker_io_ptw_pmp_2_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_a = dcache_pma_checker_io_ptw_pmp_2_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_x = dcache_pma_checker_io_ptw_pmp_2_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_w = dcache_pma_checker_io_ptw_pmp_2_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_2_cfg_r = dcache_pma_checker_io_ptw_pmp_2_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_2_addr = dcache_pma_checker_io_ptw_pmp_2_addr;
    assign dcache_pma_checker_pmp_io_pmp_2_mask = dcache_pma_checker_io_ptw_pmp_2_mask;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_l = dcache_pma_checker_io_ptw_pmp_3_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_res = dcache_pma_checker_io_ptw_pmp_3_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_a = dcache_pma_checker_io_ptw_pmp_3_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_x = dcache_pma_checker_io_ptw_pmp_3_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_w = dcache_pma_checker_io_ptw_pmp_3_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_3_cfg_r = dcache_pma_checker_io_ptw_pmp_3_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_3_addr = dcache_pma_checker_io_ptw_pmp_3_addr;
    assign dcache_pma_checker_pmp_io_pmp_3_mask = dcache_pma_checker_io_ptw_pmp_3_mask;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_l = dcache_pma_checker_io_ptw_pmp_4_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_res = dcache_pma_checker_io_ptw_pmp_4_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_a = dcache_pma_checker_io_ptw_pmp_4_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_x = dcache_pma_checker_io_ptw_pmp_4_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_w = dcache_pma_checker_io_ptw_pmp_4_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_4_cfg_r = dcache_pma_checker_io_ptw_pmp_4_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_4_addr = dcache_pma_checker_io_ptw_pmp_4_addr;
    assign dcache_pma_checker_pmp_io_pmp_4_mask = dcache_pma_checker_io_ptw_pmp_4_mask;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_l = dcache_pma_checker_io_ptw_pmp_5_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_res = dcache_pma_checker_io_ptw_pmp_5_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_a = dcache_pma_checker_io_ptw_pmp_5_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_x = dcache_pma_checker_io_ptw_pmp_5_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_w = dcache_pma_checker_io_ptw_pmp_5_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_5_cfg_r = dcache_pma_checker_io_ptw_pmp_5_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_5_addr = dcache_pma_checker_io_ptw_pmp_5_addr;
    assign dcache_pma_checker_pmp_io_pmp_5_mask = dcache_pma_checker_io_ptw_pmp_5_mask;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_l = dcache_pma_checker_io_ptw_pmp_6_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_res = dcache_pma_checker_io_ptw_pmp_6_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_a = dcache_pma_checker_io_ptw_pmp_6_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_x = dcache_pma_checker_io_ptw_pmp_6_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_w = dcache_pma_checker_io_ptw_pmp_6_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_6_cfg_r = dcache_pma_checker_io_ptw_pmp_6_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_6_addr = dcache_pma_checker_io_ptw_pmp_6_addr;
    assign dcache_pma_checker_pmp_io_pmp_6_mask = dcache_pma_checker_io_ptw_pmp_6_mask;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_l = dcache_pma_checker_io_ptw_pmp_7_cfg_l;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_res = dcache_pma_checker_io_ptw_pmp_7_cfg_res;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_a = dcache_pma_checker_io_ptw_pmp_7_cfg_a;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_x = dcache_pma_checker_io_ptw_pmp_7_cfg_x;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_w = dcache_pma_checker_io_ptw_pmp_7_cfg_w;
    assign dcache_pma_checker_pmp_io_pmp_7_cfg_r = dcache_pma_checker_io_ptw_pmp_7_cfg_r;
    assign dcache_pma_checker_pmp_io_pmp_7_addr = dcache_pma_checker_io_ptw_pmp_7_addr;
    assign dcache_pma_checker_pmp_io_pmp_7_mask = dcache_pma_checker_io_ptw_pmp_7_mask;
    assign dcache_pma_checker_pmp_io_addr = dcache__pma_checker_mpu_physaddr_31to0;
    assign dcache_pma_checker_pmp_io_size = dcache_pma_checker_io_req_bits_size;
    assign dcache__pma_checker_pmp_io_r = dcache_pma_checker_pmp_io_r;
    assign dcache__pma_checker_pmp_io_w = dcache_pma_checker_pmp_io_w;
    assign dcache__pma_checker_pmp_io_x = dcache_pma_checker_pmp_io_x;
     
  assign  dcache__pma_checker_mpu_physaddr_31to0 = dcache_pma_checker_mpu_physaddr [31:0]; 
  assign  dcache__pma_checker_mpu_priv_1to0 = dcache_pma_checker_mpu_priv [1:0]; 
    wire dcache_pma_checker__legal_address_WIRE_0 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_1 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_2 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_3 =({1'h0, dcache_pma_checker_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_4 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_5 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire dcache_pma_checker__legal_address_WIRE_6 =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0; 
    wire dcache_pma_checker_legal_address = dcache_pma_checker__legal_address_WIRE_0 | dcache_pma_checker__legal_address_WIRE_1 | dcache_pma_checker__legal_address_WIRE_2 | dcache_pma_checker__legal_address_WIRE_3 | dcache_pma_checker__legal_address_WIRE_4 | dcache_pma_checker__legal_address_WIRE_5 | dcache_pma_checker__legal_address_WIRE_6 ; 
    wire dcache_pma_checker__cacheable_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'h80000000)==35'h0|1'h0; 
    wire dcache_pma_checker_cacheable = dcache_pma_checker_legal_address & dcache_pma_checker__cacheable_WIRE ; 
    wire dcache_pma_checker_newEntry_c = dcache_pma_checker_cacheable ; 
    wire dcache_pma_checker_homogeneous =({1'h0, dcache_pma_checker_mpu_physaddr }&35'h7FFFFF000)==35'h0|1'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire dcache_pma_checker_deny_access_to_debug = dcache_pma_checker_mpu_priv <=3'h3&({1'h0, dcache_pma_checker_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire dcache_pma_checker_prot_r = dcache_pma_checker_legal_address & dcache_pma_checker_deny_access_to_debug ==1'h0& dcache__pma_checker_pmp_io_r ; 
    wire dcache_pma_checker_newEntry_pr = dcache_pma_checker_prot_r ; 
    wire dcache_pma_checker__prot_w_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_pma_checker_prot_w = dcache_pma_checker_legal_address & dcache_pma_checker__prot_w_WIRE & dcache_pma_checker_deny_access_to_debug ==1'h0& dcache__pma_checker_pmp_io_w ; 
    wire dcache_pma_checker_newEntry_pw = dcache_pma_checker_prot_w ; 
    wire dcache_pma_checker__prot_pp_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_pma_checker_prot_pp = dcache_pma_checker_legal_address & dcache_pma_checker__prot_pp_WIRE ; 
    wire dcache_pma_checker_newEntry_ppp = dcache_pma_checker_prot_pp ; 
    wire dcache_pma_checker__prot_al_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire dcache_pma_checker_prot_al = dcache_pma_checker_legal_address & dcache_pma_checker__prot_al_WIRE ; 
    wire dcache_pma_checker_newEntry_pal = dcache_pma_checker_prot_al ; 
    wire dcache_pma_checker__prot_aa_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire dcache_pma_checker_prot_aa = dcache_pma_checker_legal_address & dcache_pma_checker__prot_aa_WIRE ; 
    wire dcache_pma_checker_newEntry_paa = dcache_pma_checker_prot_aa ; 
    wire dcache_pma_checker__prot_x_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hCA000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire dcache_pma_checker_prot_x = dcache_pma_checker_legal_address & dcache_pma_checker__prot_x_WIRE & dcache_pma_checker_deny_access_to_debug ==1'h0& dcache__pma_checker_pmp_io_x ; 
    wire dcache_pma_checker_newEntry_px = dcache_pma_checker_prot_x ; 
    wire dcache_pma_checker__prot_eff_WIRE =({1'h0, dcache_pma_checker_mpu_physaddr }&35'hCA012000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_pma_checker_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|1'h0; 
    wire dcache_pma_checker_prot_eff = dcache_pma_checker_legal_address & dcache_pma_checker__prot_eff_WIRE ; 
    wire dcache_pma_checker_newEntry_eff = dcache_pma_checker_prot_eff ; 
    wire[20:0] dcache__GEN_40 = dcache_pma_checker_sectored_entries_0_0_tag_vpn ^ dcache_pma_checker_vpn ; 
    wire dcache_pma_checker_sector_hits_0 =( dcache_pma_checker_sectored_entries_0_0_valid_0 | dcache_pma_checker_sectored_entries_0_0_valid_1 | dcache_pma_checker_sectored_entries_0_0_valid_2 | dcache_pma_checker_sectored_entries_0_0_valid_3 )& dcache__GEN_40 [20:2]==19'h0& dcache_pma_checker_sectored_entries_0_0_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_superpage_hits_0 = dcache_pma_checker_superpage_entries_0_valid_0 &( dcache_pma_checker_superpage_entries_0_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_0_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_superpage_hits_1 = dcache_pma_checker_superpage_entries_1_valid_0 &( dcache_pma_checker_superpage_entries_1_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_1_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_superpage_hits_2 = dcache_pma_checker_superpage_entries_2_valid_0 &( dcache_pma_checker_superpage_entries_2_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_2_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_superpage_hits_3 = dcache_pma_checker_superpage_entries_3_valid_0 &( dcache_pma_checker_superpage_entries_3_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_3_tag_v == dcache_pma_checker_priv_v ; 
    wire[1:0] dcache_pma_checker_hitsVec_idx = dcache_pma_checker_vpn [1:0]; 
    wire[20:0] dcache__GEN_41 = dcache_pma_checker_sectored_entries_0_0_tag_vpn ^ dcache_pma_checker_vpn ; 
    reg dcache_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( dcache_pma_checker_hitsVec_idx )
              2 'b00: 
                  dcache_casez_tmp_1  = dcache_pma_checker_sectored_entries_0_0_valid_0 ;
              2 'b01: 
                  dcache_casez_tmp_1  = dcache_pma_checker_sectored_entries_0_0_valid_1 ;
              2 'b10: 
                  dcache_casez_tmp_1  = dcache_pma_checker_sectored_entries_0_0_valid_2 ;
              default : 
                  dcache_casez_tmp_1  = dcache_pma_checker_sectored_entries_0_0_valid_3 ;endcase
         end
    wire dcache_pma_checker_hitsVec_0 = dcache_pma_checker_vm_enabled & dcache_casez_tmp_1 & dcache__GEN_41 [20:2]==19'h0& dcache_pma_checker_sectored_entries_0_0_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_hitsVec_1 = dcache_pma_checker_vm_enabled & dcache_pma_checker_superpage_entries_0_valid_0 &( dcache_pma_checker_superpage_entries_0_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_0_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_hitsVec_2 = dcache_pma_checker_vm_enabled & dcache_pma_checker_superpage_entries_1_valid_0 &( dcache_pma_checker_superpage_entries_1_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_1_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_hitsVec_3 = dcache_pma_checker_vm_enabled & dcache_pma_checker_superpage_entries_2_valid_0 &( dcache_pma_checker_superpage_entries_2_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_2_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_hitsVec_4 = dcache_pma_checker_vm_enabled & dcache_pma_checker_superpage_entries_3_valid_0 &( dcache_pma_checker_superpage_entries_3_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_superpage_entries_3_tag_v == dcache_pma_checker_priv_v ; 
    wire dcache_pma_checker_hitsVec_5 = dcache_pma_checker_vm_enabled & dcache_pma_checker_special_entry_valid_0 &( dcache_pma_checker_special_entry_tag_vpn ^ dcache_pma_checker_vpn )==21'h0& dcache_pma_checker_special_entry_tag_v == dcache_pma_checker_priv_v ; 
    wire[1:0] dcache_pma_checker_real_hits_lo_hi ={ dcache_pma_checker_hitsVec_2 , dcache_pma_checker_hitsVec_1 }; 
    wire[2:0] dcache_pma_checker_real_hits_lo ={ dcache_pma_checker_real_hits_lo_hi , dcache_pma_checker_hitsVec_0 }; 
    wire[1:0] dcache_pma_checker_real_hits_hi_hi ={ dcache_pma_checker_hitsVec_5 , dcache_pma_checker_hitsVec_4 }; 
    wire[2:0] dcache_pma_checker_real_hits_hi ={ dcache_pma_checker_real_hits_hi_hi , dcache_pma_checker_hitsVec_3 }; 
    wire[5:0] dcache_pma_checker_real_hits ={ dcache_pma_checker_real_hits_hi , dcache_pma_checker_real_hits_lo }; 
    wire[6:0] dcache_pma_checker_hits ={ dcache_pma_checker_vm_enabled ==1'h0, dcache_pma_checker_real_hits }; 
    wire dcache_pma_checker_refill_v = dcache_pma_checker_r_vstage1_en | dcache_pma_checker_r_stage2_en ; 
    wire[19:0] dcache_pma_checker_newEntry_ppn = dcache_pma_checker_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire dcache_pma_checker_newEntry_g = dcache_pma_checker_io_ptw_resp_bits_pte_g & dcache_pma_checker_io_ptw_resp_bits_pte_v ; 
    wire dcache_pma_checker_newEntry_ae_stage2 = dcache_pma_checker_io_ptw_resp_bits_ae_final & dcache_pma_checker_io_ptw_resp_bits_gpa_is_pte & dcache_pma_checker_r_stage2_en ; 
    wire dcache_pma_checker_newEntry_sr = dcache_pma_checker_io_ptw_resp_bits_pte_v &( dcache_pma_checker_io_ptw_resp_bits_pte_r | dcache_pma_checker_io_ptw_resp_bits_pte_x & dcache_pma_checker_io_ptw_resp_bits_pte_w ==1'h0)& dcache_pma_checker_io_ptw_resp_bits_pte_a & dcache_pma_checker_io_ptw_resp_bits_pte_r ; 
    wire dcache_pma_checker_newEntry_sw = dcache_pma_checker_io_ptw_resp_bits_pte_v &( dcache_pma_checker_io_ptw_resp_bits_pte_r | dcache_pma_checker_io_ptw_resp_bits_pte_x & dcache_pma_checker_io_ptw_resp_bits_pte_w ==1'h0)& dcache_pma_checker_io_ptw_resp_bits_pte_a & dcache_pma_checker_io_ptw_resp_bits_pte_w & dcache_pma_checker_io_ptw_resp_bits_pte_d ; 
    wire dcache_pma_checker_newEntry_sx = dcache_pma_checker_io_ptw_resp_bits_pte_v &( dcache_pma_checker_io_ptw_resp_bits_pte_r | dcache_pma_checker_io_ptw_resp_bits_pte_x & dcache_pma_checker_io_ptw_resp_bits_pte_w ==1'h0)& dcache_pma_checker_io_ptw_resp_bits_pte_a & dcache_pma_checker_io_ptw_resp_bits_pte_x ; 
    wire dcache__GEN_42 = dcache_pma_checker_io_ptw_resp_bits_homogeneous ==1'h0&1'h1; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_lo_hi ={ dcache_pma_checker_special_entry_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_special_entry_data_0_lo_lo ={ dcache_pma_checker_special_entry_data_0_lo_lo_hi , dcache_pma_checker_special_entry_data_0_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_hi_lo ={ dcache_pma_checker_special_entry_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_lo_hi_hi ={ dcache_pma_checker_special_entry_data_0_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_special_entry_data_0_lo_hi ={ dcache_pma_checker_special_entry_data_0_lo_hi_hi , dcache_pma_checker_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_special_entry_data_0_lo ={ dcache_pma_checker_special_entry_data_0_lo_hi , dcache_pma_checker_special_entry_data_0_lo_lo }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_lo_lo ={ dcache_pma_checker_special_entry_data_0_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_lo_hi ={ dcache_pma_checker_special_entry_data_0_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_special_entry_data_0_hi_lo ={ dcache_pma_checker_special_entry_data_0_hi_lo_hi , dcache_pma_checker_special_entry_data_0_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_special_entry_data_0_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_special_entry_data_0_hi_hi_lo ={ dcache_pma_checker_special_entry_data_0_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_special_entry_data_0_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_special_entry_data_0_hi_hi_hi ={ dcache_pma_checker_special_entry_data_0_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_special_entry_data_0_hi_hi ={ dcache_pma_checker_special_entry_data_0_hi_hi_hi , dcache_pma_checker_special_entry_data_0_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_special_entry_data_0_hi ={ dcache_pma_checker_special_entry_data_0_hi_hi , dcache_pma_checker_special_entry_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_43 ={ dcache_pma_checker_special_entry_data_0_hi , dcache_pma_checker_special_entry_data_0_lo }; 
    wire dcache__GEN_44 = dcache_pma_checker_do_refill &~ dcache__GEN_42 ; 
    wire dcache__GEN_45 = dcache_pma_checker_io_ptw_resp_bits_level <2'h2; 
    wire dcache__GEN_46 = dcache__GEN_44 & dcache__GEN_45 ; 
    wire dcache__GEN_47 = dcache_pma_checker_r_superpage_repl_addr ==2'h0; 
    wire[1:0] dcache__GEN_48 ={1'h0, dcache_pma_checker_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_0_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_lo_hi , dcache_pma_checker_superpage_entries_0_data_0_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_0_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_0_data_0_lo ={ dcache_pma_checker_superpage_entries_0_data_0_lo_hi , dcache_pma_checker_superpage_entries_0_data_0_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo ={ dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi ={ dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_0_data_0_hi_lo ={ dcache_pma_checker_superpage_entries_0_data_0_hi_lo_hi , dcache_pma_checker_superpage_entries_0_data_0_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo ={ dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi ={ dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_superpage_entries_0_data_0_hi_hi ={ dcache_pma_checker_superpage_entries_0_data_0_hi_hi_hi , dcache_pma_checker_superpage_entries_0_data_0_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_superpage_entries_0_data_0_hi ={ dcache_pma_checker_superpage_entries_0_data_0_hi_hi , dcache_pma_checker_superpage_entries_0_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_49 ={ dcache_pma_checker_superpage_entries_0_data_0_hi , dcache_pma_checker_superpage_entries_0_data_0_lo }; 
    wire dcache__GEN_50 = dcache_pma_checker_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_51 = dcache_pma_checker_r_superpage_repl_addr ==2'h1; 
    wire[1:0] dcache__GEN_52 ={1'h0, dcache_pma_checker_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_1_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_lo_hi , dcache_pma_checker_superpage_entries_1_data_0_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_1_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_1_data_0_lo ={ dcache_pma_checker_superpage_entries_1_data_0_lo_hi , dcache_pma_checker_superpage_entries_1_data_0_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo ={ dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi ={ dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_1_data_0_hi_lo ={ dcache_pma_checker_superpage_entries_1_data_0_hi_lo_hi , dcache_pma_checker_superpage_entries_1_data_0_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo ={ dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi ={ dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_superpage_entries_1_data_0_hi_hi ={ dcache_pma_checker_superpage_entries_1_data_0_hi_hi_hi , dcache_pma_checker_superpage_entries_1_data_0_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_superpage_entries_1_data_0_hi ={ dcache_pma_checker_superpage_entries_1_data_0_hi_hi , dcache_pma_checker_superpage_entries_1_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_53 ={ dcache_pma_checker_superpage_entries_1_data_0_hi , dcache_pma_checker_superpage_entries_1_data_0_lo }; 
    wire dcache__GEN_54 = dcache_pma_checker_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_55 = dcache_pma_checker_r_superpage_repl_addr ==2'h2; 
    wire[1:0] dcache__GEN_56 ={1'h0, dcache_pma_checker_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_2_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_lo_hi , dcache_pma_checker_superpage_entries_2_data_0_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_2_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_2_data_0_lo ={ dcache_pma_checker_superpage_entries_2_data_0_lo_hi , dcache_pma_checker_superpage_entries_2_data_0_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo ={ dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi ={ dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_2_data_0_hi_lo ={ dcache_pma_checker_superpage_entries_2_data_0_hi_lo_hi , dcache_pma_checker_superpage_entries_2_data_0_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo ={ dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi ={ dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_superpage_entries_2_data_0_hi_hi ={ dcache_pma_checker_superpage_entries_2_data_0_hi_hi_hi , dcache_pma_checker_superpage_entries_2_data_0_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_superpage_entries_2_data_0_hi ={ dcache_pma_checker_superpage_entries_2_data_0_hi_hi , dcache_pma_checker_superpage_entries_2_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_57 ={ dcache_pma_checker_superpage_entries_2_data_0_hi , dcache_pma_checker_superpage_entries_2_data_0_lo }; 
    wire dcache__GEN_58 = dcache_pma_checker_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_59 =& dcache_pma_checker_r_superpage_repl_addr ; 
    wire[1:0] dcache__GEN_60 ={1'h0, dcache_pma_checker_io_ptw_resp_bits_level [0]}; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi ={ dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_superpage_entries_3_data_0_lo_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_lo_hi , dcache_pma_checker_superpage_entries_3_data_0_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_3_data_0_lo_hi ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi_hi , dcache_pma_checker_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_superpage_entries_3_data_0_lo ={ dcache_pma_checker_superpage_entries_3_data_0_lo_hi , dcache_pma_checker_superpage_entries_3_data_0_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo ={ dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi ={ dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_superpage_entries_3_data_0_hi_lo ={ dcache_pma_checker_superpage_entries_3_data_0_hi_lo_hi , dcache_pma_checker_superpage_entries_3_data_0_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo ={ dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi ={ dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_superpage_entries_3_data_0_hi_hi ={ dcache_pma_checker_superpage_entries_3_data_0_hi_hi_hi , dcache_pma_checker_superpage_entries_3_data_0_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_superpage_entries_3_data_0_hi ={ dcache_pma_checker_superpage_entries_3_data_0_hi_hi , dcache_pma_checker_superpage_entries_3_data_0_hi_lo }; 
    wire[41:0] dcache__GEN_61 ={ dcache_pma_checker_superpage_entries_3_data_0_hi , dcache_pma_checker_superpage_entries_3_data_0_lo }; 
    wire dcache__GEN_62 = dcache_pma_checker_invalidate_refill  ? 1'h0:1'h1; 
    wire dcache__GEN_63 = dcache__GEN_44 &~ dcache__GEN_45 ; 
    wire dcache__GEN_64 = dcache_pma_checker_r_sectored_hit_valid ==1'h0; 
    wire[1:0] dcache_pma_checker_idx = dcache_pma_checker_r_refill_tag [1:0]; 
    wire dcache__GEN_65 = dcache_pma_checker_idx ==2'h0; 
    wire dcache__GEN_66 = dcache_pma_checker_idx ==2'h1; 
    wire dcache__GEN_67 = dcache_pma_checker_idx ==2'h2; 
    wire dcache__GEN_68 =& dcache_pma_checker_idx ; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_lo ={ dcache_pma_checker_newEntry_c , dcache_pma_checker_newEntry_fragmented_superpage }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi_hi ={ dcache_pma_checker_newEntry_pal , dcache_pma_checker_newEntry_paa }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi ={ dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi_hi , dcache_pma_checker_newEntry_eff }; 
    wire[4:0] dcache_pma_checker_sectored_entries_0_0_data_lo_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_lo_hi , dcache_pma_checker_sectored_entries_0_0_data_lo_lo_lo }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo_hi ={ dcache_pma_checker_newEntry_px , dcache_pma_checker_newEntry_pr }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo_hi , dcache_pma_checker_newEntry_ppp }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi_hi ={ dcache_pma_checker_newEntry_hx , dcache_pma_checker_newEntry_hr }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi_hi , dcache_pma_checker_newEntry_pw }; 
    wire[5:0] dcache_pma_checker_sectored_entries_0_0_data_lo_hi ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi_hi , dcache_pma_checker_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] dcache_pma_checker_sectored_entries_0_0_data_lo ={ dcache_pma_checker_sectored_entries_0_0_data_lo_hi , dcache_pma_checker_sectored_entries_0_0_data_lo_lo }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo_hi ={ dcache_pma_checker_newEntry_sx , dcache_pma_checker_newEntry_sr }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo ={ dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo_hi , dcache_pma_checker_newEntry_hw }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi_hi ={ dcache_pma_checker_newEntry_pf , dcache_pma_checker_newEntry_gf }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi ={ dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi_hi , dcache_pma_checker_newEntry_sw }; 
    wire[5:0] dcache_pma_checker_sectored_entries_0_0_data_hi_lo ={ dcache_pma_checker_sectored_entries_0_0_data_hi_lo_hi , dcache_pma_checker_sectored_entries_0_0_data_hi_lo_lo }; 
    wire[1:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo_hi ={ dcache_pma_checker_newEntry_ae_ptw , dcache_pma_checker_newEntry_ae_final }; 
    wire[2:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo ={ dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo_hi , dcache_pma_checker_newEntry_ae_stage2 }; 
    wire[20:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi_hi ={ dcache_pma_checker_newEntry_ppn , dcache_pma_checker_newEntry_u }; 
    wire[21:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi ={ dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi_hi , dcache_pma_checker_newEntry_g }; 
    wire[24:0] dcache_pma_checker_sectored_entries_0_0_data_hi_hi ={ dcache_pma_checker_sectored_entries_0_0_data_hi_hi_hi , dcache_pma_checker_sectored_entries_0_0_data_hi_hi_lo }; 
    wire[30:0] dcache_pma_checker_sectored_entries_0_0_data_hi ={ dcache_pma_checker_sectored_entries_0_0_data_hi_hi , dcache_pma_checker_sectored_entries_0_0_data_hi_lo }; 
    wire[41:0] dcache__GEN_69 ={ dcache_pma_checker_sectored_entries_0_0_data_hi , dcache_pma_checker_sectored_entries_0_0_data_lo }; 
    wire dcache__GEN_70 = dcache_pma_checker_idx ==2'h0; 
    wire dcache__GEN_71 = dcache_pma_checker_idx ==2'h1; 
    wire dcache__GEN_72 = dcache_pma_checker_idx ==2'h2; 
    wire dcache__GEN_73 =& dcache_pma_checker_idx ; reg[41:0] dcache_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( dcache_pma_checker_vpn [1:0])
              2 'b00: 
                  dcache_casez_tmp_2  = dcache_pma_checker_sectored_entries_0_0_data_0 ;
              2 'b01: 
                  dcache_casez_tmp_2  = dcache_pma_checker_sectored_entries_0_0_data_1 ;
              2 'b10: 
                  dcache_casez_tmp_2  = dcache_pma_checker_sectored_entries_0_0_data_2 ;
              default : 
                  dcache_casez_tmp_2  = dcache_pma_checker_sectored_entries_0_0_data_3 ;endcase
         end
    wire[41:0] dcache_pma_checker__entries_WIRE_1 = dcache_casez_tmp_2 ; 
    wire dcache_pma_checker__entries_WIRE_fragmented_superpage = dcache_pma_checker__entries_WIRE_1 [0]; 
    wire dcache_pma_checker__entries_WIRE_c = dcache_pma_checker__entries_WIRE_1 [1]; 
    wire dcache_pma_checker__entries_WIRE_eff = dcache_pma_checker__entries_WIRE_1 [2]; 
    wire dcache_pma_checker__entries_WIRE_paa = dcache_pma_checker__entries_WIRE_1 [3]; 
    wire dcache_pma_checker__entries_WIRE_pal = dcache_pma_checker__entries_WIRE_1 [4]; 
    wire dcache_pma_checker__entries_WIRE_ppp = dcache_pma_checker__entries_WIRE_1 [5]; 
    wire dcache_pma_checker__entries_WIRE_pr = dcache_pma_checker__entries_WIRE_1 [6]; 
    wire dcache_pma_checker__entries_WIRE_px = dcache_pma_checker__entries_WIRE_1 [7]; 
    wire dcache_pma_checker__entries_WIRE_pw = dcache_pma_checker__entries_WIRE_1 [8]; 
    wire dcache_pma_checker__entries_WIRE_hr = dcache_pma_checker__entries_WIRE_1 [9]; 
    wire dcache_pma_checker__entries_WIRE_hx = dcache_pma_checker__entries_WIRE_1 [10]; 
    wire dcache_pma_checker__entries_WIRE_hw = dcache_pma_checker__entries_WIRE_1 [11]; 
    wire dcache_pma_checker__entries_WIRE_sr = dcache_pma_checker__entries_WIRE_1 [12]; 
    wire dcache_pma_checker__entries_WIRE_sx = dcache_pma_checker__entries_WIRE_1 [13]; 
    wire dcache_pma_checker__entries_WIRE_sw = dcache_pma_checker__entries_WIRE_1 [14]; 
    wire dcache_pma_checker__entries_WIRE_gf = dcache_pma_checker__entries_WIRE_1 [15]; 
    wire dcache_pma_checker__entries_WIRE_pf = dcache_pma_checker__entries_WIRE_1 [16]; 
    wire dcache_pma_checker__entries_WIRE_ae_stage2 = dcache_pma_checker__entries_WIRE_1 [17]; 
    wire dcache_pma_checker__entries_WIRE_ae_final = dcache_pma_checker__entries_WIRE_1 [18]; 
    wire dcache_pma_checker__entries_WIRE_ae_ptw = dcache_pma_checker__entries_WIRE_1 [19]; 
    wire dcache_pma_checker__entries_WIRE_g = dcache_pma_checker__entries_WIRE_1 [20]; 
    wire dcache_pma_checker__entries_WIRE_u = dcache_pma_checker__entries_WIRE_1 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_ppn = dcache_pma_checker__entries_WIRE_1 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_io_y_ppn = dcache_pma_checker_entries_barrier_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_io_y_u = dcache_pma_checker_entries_barrier_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_io_y_g = dcache_pma_checker_entries_barrier_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_ptw = dcache_pma_checker_entries_barrier_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_final = dcache_pma_checker_entries_barrier_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pf = dcache_pma_checker_entries_barrier_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_io_y_gf = dcache_pma_checker_entries_barrier_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sw = dcache_pma_checker_entries_barrier_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sx = dcache_pma_checker_entries_barrier_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_io_y_sr = dcache_pma_checker_entries_barrier_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hw = dcache_pma_checker_entries_barrier_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hx = dcache_pma_checker_entries_barrier_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_io_y_hr = dcache_pma_checker_entries_barrier_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pw = dcache_pma_checker_entries_barrier_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_io_y_px = dcache_pma_checker_entries_barrier_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pr = dcache_pma_checker_entries_barrier_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_io_y_ppp = dcache_pma_checker_entries_barrier_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_io_y_pal = dcache_pma_checker_entries_barrier_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_io_y_paa = dcache_pma_checker_entries_barrier_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_io_y_eff = dcache_pma_checker_entries_barrier_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_io_y_c = dcache_pma_checker_entries_barrier_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_io_x_fragmented_superpage ;
     
    wire dcache_pma_checker__entries_WIRE_2_fragmented_superpage = dcache_pma_checker__entries_WIRE_3 [0]; 
    wire dcache_pma_checker__entries_WIRE_2_c = dcache_pma_checker__entries_WIRE_3 [1]; 
    wire dcache_pma_checker__entries_WIRE_2_eff = dcache_pma_checker__entries_WIRE_3 [2]; 
    wire dcache_pma_checker__entries_WIRE_2_paa = dcache_pma_checker__entries_WIRE_3 [3]; 
    wire dcache_pma_checker__entries_WIRE_2_pal = dcache_pma_checker__entries_WIRE_3 [4]; 
    wire dcache_pma_checker__entries_WIRE_2_ppp = dcache_pma_checker__entries_WIRE_3 [5]; 
    wire dcache_pma_checker__entries_WIRE_2_pr = dcache_pma_checker__entries_WIRE_3 [6]; 
    wire dcache_pma_checker__entries_WIRE_2_px = dcache_pma_checker__entries_WIRE_3 [7]; 
    wire dcache_pma_checker__entries_WIRE_2_pw = dcache_pma_checker__entries_WIRE_3 [8]; 
    wire dcache_pma_checker__entries_WIRE_2_hr = dcache_pma_checker__entries_WIRE_3 [9]; 
    wire dcache_pma_checker__entries_WIRE_2_hx = dcache_pma_checker__entries_WIRE_3 [10]; 
    wire dcache_pma_checker__entries_WIRE_2_hw = dcache_pma_checker__entries_WIRE_3 [11]; 
    wire dcache_pma_checker__entries_WIRE_2_sr = dcache_pma_checker__entries_WIRE_3 [12]; 
    wire dcache_pma_checker__entries_WIRE_2_sx = dcache_pma_checker__entries_WIRE_3 [13]; 
    wire dcache_pma_checker__entries_WIRE_2_sw = dcache_pma_checker__entries_WIRE_3 [14]; 
    wire dcache_pma_checker__entries_WIRE_2_gf = dcache_pma_checker__entries_WIRE_3 [15]; 
    wire dcache_pma_checker__entries_WIRE_2_pf = dcache_pma_checker__entries_WIRE_3 [16]; 
    wire dcache_pma_checker__entries_WIRE_2_ae_stage2 = dcache_pma_checker__entries_WIRE_3 [17]; 
    wire dcache_pma_checker__entries_WIRE_2_ae_final = dcache_pma_checker__entries_WIRE_3 [18]; 
    wire dcache_pma_checker__entries_WIRE_2_ae_ptw = dcache_pma_checker__entries_WIRE_3 [19]; 
    wire dcache_pma_checker__entries_WIRE_2_g = dcache_pma_checker__entries_WIRE_3 [20]; 
    wire dcache_pma_checker__entries_WIRE_2_u = dcache_pma_checker__entries_WIRE_3 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_2_ppn = dcache_pma_checker__entries_WIRE_3 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_1_io_y_ppn = dcache_pma_checker_entries_barrier_1_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_u = dcache_pma_checker_entries_barrier_1_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_g = dcache_pma_checker_entries_barrier_1_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_ptw = dcache_pma_checker_entries_barrier_1_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_final = dcache_pma_checker_entries_barrier_1_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_1_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pf = dcache_pma_checker_entries_barrier_1_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_gf = dcache_pma_checker_entries_barrier_1_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sw = dcache_pma_checker_entries_barrier_1_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sx = dcache_pma_checker_entries_barrier_1_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_sr = dcache_pma_checker_entries_barrier_1_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hw = dcache_pma_checker_entries_barrier_1_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hx = dcache_pma_checker_entries_barrier_1_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_hr = dcache_pma_checker_entries_barrier_1_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pw = dcache_pma_checker_entries_barrier_1_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_px = dcache_pma_checker_entries_barrier_1_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pr = dcache_pma_checker_entries_barrier_1_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_ppp = dcache_pma_checker_entries_barrier_1_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_pal = dcache_pma_checker_entries_barrier_1_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_paa = dcache_pma_checker_entries_barrier_1_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_eff = dcache_pma_checker_entries_barrier_1_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_c = dcache_pma_checker_entries_barrier_1_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_1_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_1_io_x_fragmented_superpage ;
     
    wire dcache_pma_checker__entries_WIRE_4_fragmented_superpage = dcache_pma_checker__entries_WIRE_5 [0]; 
    wire dcache_pma_checker__entries_WIRE_4_c = dcache_pma_checker__entries_WIRE_5 [1]; 
    wire dcache_pma_checker__entries_WIRE_4_eff = dcache_pma_checker__entries_WIRE_5 [2]; 
    wire dcache_pma_checker__entries_WIRE_4_paa = dcache_pma_checker__entries_WIRE_5 [3]; 
    wire dcache_pma_checker__entries_WIRE_4_pal = dcache_pma_checker__entries_WIRE_5 [4]; 
    wire dcache_pma_checker__entries_WIRE_4_ppp = dcache_pma_checker__entries_WIRE_5 [5]; 
    wire dcache_pma_checker__entries_WIRE_4_pr = dcache_pma_checker__entries_WIRE_5 [6]; 
    wire dcache_pma_checker__entries_WIRE_4_px = dcache_pma_checker__entries_WIRE_5 [7]; 
    wire dcache_pma_checker__entries_WIRE_4_pw = dcache_pma_checker__entries_WIRE_5 [8]; 
    wire dcache_pma_checker__entries_WIRE_4_hr = dcache_pma_checker__entries_WIRE_5 [9]; 
    wire dcache_pma_checker__entries_WIRE_4_hx = dcache_pma_checker__entries_WIRE_5 [10]; 
    wire dcache_pma_checker__entries_WIRE_4_hw = dcache_pma_checker__entries_WIRE_5 [11]; 
    wire dcache_pma_checker__entries_WIRE_4_sr = dcache_pma_checker__entries_WIRE_5 [12]; 
    wire dcache_pma_checker__entries_WIRE_4_sx = dcache_pma_checker__entries_WIRE_5 [13]; 
    wire dcache_pma_checker__entries_WIRE_4_sw = dcache_pma_checker__entries_WIRE_5 [14]; 
    wire dcache_pma_checker__entries_WIRE_4_gf = dcache_pma_checker__entries_WIRE_5 [15]; 
    wire dcache_pma_checker__entries_WIRE_4_pf = dcache_pma_checker__entries_WIRE_5 [16]; 
    wire dcache_pma_checker__entries_WIRE_4_ae_stage2 = dcache_pma_checker__entries_WIRE_5 [17]; 
    wire dcache_pma_checker__entries_WIRE_4_ae_final = dcache_pma_checker__entries_WIRE_5 [18]; 
    wire dcache_pma_checker__entries_WIRE_4_ae_ptw = dcache_pma_checker__entries_WIRE_5 [19]; 
    wire dcache_pma_checker__entries_WIRE_4_g = dcache_pma_checker__entries_WIRE_5 [20]; 
    wire dcache_pma_checker__entries_WIRE_4_u = dcache_pma_checker__entries_WIRE_5 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_4_ppn = dcache_pma_checker__entries_WIRE_5 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_2_io_y_ppn = dcache_pma_checker_entries_barrier_2_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_u = dcache_pma_checker_entries_barrier_2_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_g = dcache_pma_checker_entries_barrier_2_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_ptw = dcache_pma_checker_entries_barrier_2_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_final = dcache_pma_checker_entries_barrier_2_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_2_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pf = dcache_pma_checker_entries_barrier_2_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_gf = dcache_pma_checker_entries_barrier_2_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sw = dcache_pma_checker_entries_barrier_2_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sx = dcache_pma_checker_entries_barrier_2_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_sr = dcache_pma_checker_entries_barrier_2_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hw = dcache_pma_checker_entries_barrier_2_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hx = dcache_pma_checker_entries_barrier_2_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_hr = dcache_pma_checker_entries_barrier_2_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pw = dcache_pma_checker_entries_barrier_2_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_px = dcache_pma_checker_entries_barrier_2_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pr = dcache_pma_checker_entries_barrier_2_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_ppp = dcache_pma_checker_entries_barrier_2_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_pal = dcache_pma_checker_entries_barrier_2_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_paa = dcache_pma_checker_entries_barrier_2_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_eff = dcache_pma_checker_entries_barrier_2_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_c = dcache_pma_checker_entries_barrier_2_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_2_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_2_io_x_fragmented_superpage ;
     
    wire dcache_pma_checker__entries_WIRE_6_fragmented_superpage = dcache_pma_checker__entries_WIRE_7 [0]; 
    wire dcache_pma_checker__entries_WIRE_6_c = dcache_pma_checker__entries_WIRE_7 [1]; 
    wire dcache_pma_checker__entries_WIRE_6_eff = dcache_pma_checker__entries_WIRE_7 [2]; 
    wire dcache_pma_checker__entries_WIRE_6_paa = dcache_pma_checker__entries_WIRE_7 [3]; 
    wire dcache_pma_checker__entries_WIRE_6_pal = dcache_pma_checker__entries_WIRE_7 [4]; 
    wire dcache_pma_checker__entries_WIRE_6_ppp = dcache_pma_checker__entries_WIRE_7 [5]; 
    wire dcache_pma_checker__entries_WIRE_6_pr = dcache_pma_checker__entries_WIRE_7 [6]; 
    wire dcache_pma_checker__entries_WIRE_6_px = dcache_pma_checker__entries_WIRE_7 [7]; 
    wire dcache_pma_checker__entries_WIRE_6_pw = dcache_pma_checker__entries_WIRE_7 [8]; 
    wire dcache_pma_checker__entries_WIRE_6_hr = dcache_pma_checker__entries_WIRE_7 [9]; 
    wire dcache_pma_checker__entries_WIRE_6_hx = dcache_pma_checker__entries_WIRE_7 [10]; 
    wire dcache_pma_checker__entries_WIRE_6_hw = dcache_pma_checker__entries_WIRE_7 [11]; 
    wire dcache_pma_checker__entries_WIRE_6_sr = dcache_pma_checker__entries_WIRE_7 [12]; 
    wire dcache_pma_checker__entries_WIRE_6_sx = dcache_pma_checker__entries_WIRE_7 [13]; 
    wire dcache_pma_checker__entries_WIRE_6_sw = dcache_pma_checker__entries_WIRE_7 [14]; 
    wire dcache_pma_checker__entries_WIRE_6_gf = dcache_pma_checker__entries_WIRE_7 [15]; 
    wire dcache_pma_checker__entries_WIRE_6_pf = dcache_pma_checker__entries_WIRE_7 [16]; 
    wire dcache_pma_checker__entries_WIRE_6_ae_stage2 = dcache_pma_checker__entries_WIRE_7 [17]; 
    wire dcache_pma_checker__entries_WIRE_6_ae_final = dcache_pma_checker__entries_WIRE_7 [18]; 
    wire dcache_pma_checker__entries_WIRE_6_ae_ptw = dcache_pma_checker__entries_WIRE_7 [19]; 
    wire dcache_pma_checker__entries_WIRE_6_g = dcache_pma_checker__entries_WIRE_7 [20]; 
    wire dcache_pma_checker__entries_WIRE_6_u = dcache_pma_checker__entries_WIRE_7 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_6_ppn = dcache_pma_checker__entries_WIRE_7 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_3_io_y_ppn = dcache_pma_checker_entries_barrier_3_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_u = dcache_pma_checker_entries_barrier_3_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_g = dcache_pma_checker_entries_barrier_3_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_ptw = dcache_pma_checker_entries_barrier_3_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_final = dcache_pma_checker_entries_barrier_3_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_3_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pf = dcache_pma_checker_entries_barrier_3_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_gf = dcache_pma_checker_entries_barrier_3_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sw = dcache_pma_checker_entries_barrier_3_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sx = dcache_pma_checker_entries_barrier_3_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_sr = dcache_pma_checker_entries_barrier_3_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hw = dcache_pma_checker_entries_barrier_3_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hx = dcache_pma_checker_entries_barrier_3_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_hr = dcache_pma_checker_entries_barrier_3_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pw = dcache_pma_checker_entries_barrier_3_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_px = dcache_pma_checker_entries_barrier_3_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pr = dcache_pma_checker_entries_barrier_3_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_ppp = dcache_pma_checker_entries_barrier_3_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_pal = dcache_pma_checker_entries_barrier_3_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_paa = dcache_pma_checker_entries_barrier_3_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_eff = dcache_pma_checker_entries_barrier_3_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_c = dcache_pma_checker_entries_barrier_3_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_3_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_3_io_x_fragmented_superpage ;
     
    wire dcache_pma_checker__entries_WIRE_8_fragmented_superpage = dcache_pma_checker__entries_WIRE_9 [0]; 
    wire dcache_pma_checker__entries_WIRE_8_c = dcache_pma_checker__entries_WIRE_9 [1]; 
    wire dcache_pma_checker__entries_WIRE_8_eff = dcache_pma_checker__entries_WIRE_9 [2]; 
    wire dcache_pma_checker__entries_WIRE_8_paa = dcache_pma_checker__entries_WIRE_9 [3]; 
    wire dcache_pma_checker__entries_WIRE_8_pal = dcache_pma_checker__entries_WIRE_9 [4]; 
    wire dcache_pma_checker__entries_WIRE_8_ppp = dcache_pma_checker__entries_WIRE_9 [5]; 
    wire dcache_pma_checker__entries_WIRE_8_pr = dcache_pma_checker__entries_WIRE_9 [6]; 
    wire dcache_pma_checker__entries_WIRE_8_px = dcache_pma_checker__entries_WIRE_9 [7]; 
    wire dcache_pma_checker__entries_WIRE_8_pw = dcache_pma_checker__entries_WIRE_9 [8]; 
    wire dcache_pma_checker__entries_WIRE_8_hr = dcache_pma_checker__entries_WIRE_9 [9]; 
    wire dcache_pma_checker__entries_WIRE_8_hx = dcache_pma_checker__entries_WIRE_9 [10]; 
    wire dcache_pma_checker__entries_WIRE_8_hw = dcache_pma_checker__entries_WIRE_9 [11]; 
    wire dcache_pma_checker__entries_WIRE_8_sr = dcache_pma_checker__entries_WIRE_9 [12]; 
    wire dcache_pma_checker__entries_WIRE_8_sx = dcache_pma_checker__entries_WIRE_9 [13]; 
    wire dcache_pma_checker__entries_WIRE_8_sw = dcache_pma_checker__entries_WIRE_9 [14]; 
    wire dcache_pma_checker__entries_WIRE_8_gf = dcache_pma_checker__entries_WIRE_9 [15]; 
    wire dcache_pma_checker__entries_WIRE_8_pf = dcache_pma_checker__entries_WIRE_9 [16]; 
    wire dcache_pma_checker__entries_WIRE_8_ae_stage2 = dcache_pma_checker__entries_WIRE_9 [17]; 
    wire dcache_pma_checker__entries_WIRE_8_ae_final = dcache_pma_checker__entries_WIRE_9 [18]; 
    wire dcache_pma_checker__entries_WIRE_8_ae_ptw = dcache_pma_checker__entries_WIRE_9 [19]; 
    wire dcache_pma_checker__entries_WIRE_8_g = dcache_pma_checker__entries_WIRE_9 [20]; 
    wire dcache_pma_checker__entries_WIRE_8_u = dcache_pma_checker__entries_WIRE_9 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_8_ppn = dcache_pma_checker__entries_WIRE_9 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_4_io_y_ppn = dcache_pma_checker_entries_barrier_4_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_u = dcache_pma_checker_entries_barrier_4_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_g = dcache_pma_checker_entries_barrier_4_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_ptw = dcache_pma_checker_entries_barrier_4_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_final = dcache_pma_checker_entries_barrier_4_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_4_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pf = dcache_pma_checker_entries_barrier_4_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_gf = dcache_pma_checker_entries_barrier_4_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sw = dcache_pma_checker_entries_barrier_4_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sx = dcache_pma_checker_entries_barrier_4_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_sr = dcache_pma_checker_entries_barrier_4_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hw = dcache_pma_checker_entries_barrier_4_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hx = dcache_pma_checker_entries_barrier_4_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_hr = dcache_pma_checker_entries_barrier_4_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pw = dcache_pma_checker_entries_barrier_4_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_px = dcache_pma_checker_entries_barrier_4_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pr = dcache_pma_checker_entries_barrier_4_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_ppp = dcache_pma_checker_entries_barrier_4_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_pal = dcache_pma_checker_entries_barrier_4_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_paa = dcache_pma_checker_entries_barrier_4_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_eff = dcache_pma_checker_entries_barrier_4_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_c = dcache_pma_checker_entries_barrier_4_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_4_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_4_io_x_fragmented_superpage ;
     
    wire dcache_pma_checker__entries_WIRE_10_fragmented_superpage = dcache_pma_checker__entries_WIRE_11 [0]; 
    wire dcache_pma_checker__entries_WIRE_10_c = dcache_pma_checker__entries_WIRE_11 [1]; 
    wire dcache_pma_checker__entries_WIRE_10_eff = dcache_pma_checker__entries_WIRE_11 [2]; 
    wire dcache_pma_checker__entries_WIRE_10_paa = dcache_pma_checker__entries_WIRE_11 [3]; 
    wire dcache_pma_checker__entries_WIRE_10_pal = dcache_pma_checker__entries_WIRE_11 [4]; 
    wire dcache_pma_checker__entries_WIRE_10_ppp = dcache_pma_checker__entries_WIRE_11 [5]; 
    wire dcache_pma_checker__entries_WIRE_10_pr = dcache_pma_checker__entries_WIRE_11 [6]; 
    wire dcache_pma_checker__entries_WIRE_10_px = dcache_pma_checker__entries_WIRE_11 [7]; 
    wire dcache_pma_checker__entries_WIRE_10_pw = dcache_pma_checker__entries_WIRE_11 [8]; 
    wire dcache_pma_checker__entries_WIRE_10_hr = dcache_pma_checker__entries_WIRE_11 [9]; 
    wire dcache_pma_checker__entries_WIRE_10_hx = dcache_pma_checker__entries_WIRE_11 [10]; 
    wire dcache_pma_checker__entries_WIRE_10_hw = dcache_pma_checker__entries_WIRE_11 [11]; 
    wire dcache_pma_checker__entries_WIRE_10_sr = dcache_pma_checker__entries_WIRE_11 [12]; 
    wire dcache_pma_checker__entries_WIRE_10_sx = dcache_pma_checker__entries_WIRE_11 [13]; 
    wire dcache_pma_checker__entries_WIRE_10_sw = dcache_pma_checker__entries_WIRE_11 [14]; 
    wire dcache_pma_checker__entries_WIRE_10_gf = dcache_pma_checker__entries_WIRE_11 [15]; 
    wire dcache_pma_checker__entries_WIRE_10_pf = dcache_pma_checker__entries_WIRE_11 [16]; 
    wire dcache_pma_checker__entries_WIRE_10_ae_stage2 = dcache_pma_checker__entries_WIRE_11 [17]; 
    wire dcache_pma_checker__entries_WIRE_10_ae_final = dcache_pma_checker__entries_WIRE_11 [18]; 
    wire dcache_pma_checker__entries_WIRE_10_ae_ptw = dcache_pma_checker__entries_WIRE_11 [19]; 
    wire dcache_pma_checker__entries_WIRE_10_g = dcache_pma_checker__entries_WIRE_11 [20]; 
    wire dcache_pma_checker__entries_WIRE_10_u = dcache_pma_checker__entries_WIRE_11 [21]; 
    wire[19:0] dcache_pma_checker__entries_WIRE_10_ppn = dcache_pma_checker__entries_WIRE_11 [41:22];  
    
    assign  dcache_pma_checker_entries_barrier_5_io_y_ppn = dcache_pma_checker_entries_barrier_5_io_x_ppn ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_u = dcache_pma_checker_entries_barrier_5_io_x_u ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_g = dcache_pma_checker_entries_barrier_5_io_x_g ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_ptw = dcache_pma_checker_entries_barrier_5_io_x_ae_ptw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_final = dcache_pma_checker_entries_barrier_5_io_x_ae_final ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_5_io_x_ae_stage2 ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pf = dcache_pma_checker_entries_barrier_5_io_x_pf ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_gf = dcache_pma_checker_entries_barrier_5_io_x_gf ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sw = dcache_pma_checker_entries_barrier_5_io_x_sw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sx = dcache_pma_checker_entries_barrier_5_io_x_sx ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_sr = dcache_pma_checker_entries_barrier_5_io_x_sr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hw = dcache_pma_checker_entries_barrier_5_io_x_hw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hx = dcache_pma_checker_entries_barrier_5_io_x_hx ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_hr = dcache_pma_checker_entries_barrier_5_io_x_hr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pw = dcache_pma_checker_entries_barrier_5_io_x_pw ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_px = dcache_pma_checker_entries_barrier_5_io_x_px ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pr = dcache_pma_checker_entries_barrier_5_io_x_pr ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_ppp = dcache_pma_checker_entries_barrier_5_io_x_ppp ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_pal = dcache_pma_checker_entries_barrier_5_io_x_pal ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_paa = dcache_pma_checker_entries_barrier_5_io_x_paa ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_eff = dcache_pma_checker_entries_barrier_5_io_x_eff ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_c = dcache_pma_checker_entries_barrier_5_io_x_c ; 
  assign  dcache_pma_checker_entries_barrier_5_io_y_fragmented_superpage = dcache_pma_checker_entries_barrier_5_io_x_fragmented_superpage ;
    assign dcache_tlb_mpu_ppn_barrier_clock = dcache_tlb_clock;
    assign dcache_tlb_mpu_ppn_barrier_reset = dcache_tlb_reset;
    assign dcache_tlb_mpu_ppn_barrier_io_x_ppn = dcache_tlb__mpu_ppn_WIRE_ppn;
    assign dcache_tlb_mpu_ppn_barrier_io_x_u = dcache_tlb__mpu_ppn_WIRE_u;
    assign dcache_tlb_mpu_ppn_barrier_io_x_g = dcache_tlb__mpu_ppn_WIRE_g;
    assign dcache_tlb_mpu_ppn_barrier_io_x_ae_ptw = dcache_tlb__mpu_ppn_WIRE_ae_ptw;
    assign dcache_tlb_mpu_ppn_barrier_io_x_ae_final = dcache_tlb__mpu_ppn_WIRE_ae_final;
    assign dcache_tlb_mpu_ppn_barrier_io_x_ae_stage2 = dcache_tlb__mpu_ppn_WIRE_ae_stage2;
    assign dcache_tlb_mpu_ppn_barrier_io_x_pf = dcache_tlb__mpu_ppn_WIRE_pf;
    assign dcache_tlb_mpu_ppn_barrier_io_x_gf = dcache_tlb__mpu_ppn_WIRE_gf;
    assign dcache_tlb_mpu_ppn_barrier_io_x_sw = dcache_tlb__mpu_ppn_WIRE_sw;
    assign dcache_tlb_mpu_ppn_barrier_io_x_sx = dcache_tlb__mpu_ppn_WIRE_sx;
    assign dcache_tlb_mpu_ppn_barrier_io_x_sr = dcache_tlb__mpu_ppn_WIRE_sr;
    assign dcache_tlb_mpu_ppn_barrier_io_x_hw = dcache_tlb__mpu_ppn_WIRE_hw;
    assign dcache_tlb_mpu_ppn_barrier_io_x_hx = dcache_tlb__mpu_ppn_WIRE_hx;
    assign dcache_tlb_mpu_ppn_barrier_io_x_hr = dcache_tlb__mpu_ppn_WIRE_hr;
    assign dcache_tlb_mpu_ppn_barrier_io_x_pw = dcache_tlb__mpu_ppn_WIRE_pw;
    assign dcache_tlb_mpu_ppn_barrier_io_x_px = dcache_tlb__mpu_ppn_WIRE_px;
    assign dcache_tlb_mpu_ppn_barrier_io_x_pr = dcache_tlb__mpu_ppn_WIRE_pr;
    assign dcache_tlb_mpu_ppn_barrier_io_x_ppp = dcache_tlb__mpu_ppn_WIRE_ppp;
    assign dcache_tlb_mpu_ppn_barrier_io_x_pal = dcache_tlb__mpu_ppn_WIRE_pal;
    assign dcache_tlb_mpu_ppn_barrier_io_x_paa = dcache_tlb__mpu_ppn_WIRE_paa;
    assign dcache_tlb_mpu_ppn_barrier_io_x_eff = dcache_tlb__mpu_ppn_WIRE_eff;
    assign dcache_tlb_mpu_ppn_barrier_io_x_c = dcache_tlb__mpu_ppn_WIRE_c;
    assign dcache_tlb_mpu_ppn_barrier_io_x_fragmented_superpage = dcache_tlb__mpu_ppn_WIRE_fragmented_superpage;
    assign dcache__tlb_mpu_ppn_barrier_io_y_ppn = dcache_tlb_mpu_ppn_barrier_io_y_ppn;
    assign dcache_tlb_entries_barrier_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_io_x_ppn = dcache_tlb__entries_WIRE_ppn;
    assign dcache_tlb_entries_barrier_io_x_u = dcache_tlb__entries_WIRE_u;
    assign dcache_tlb_entries_barrier_io_x_g = dcache_tlb__entries_WIRE_g;
    assign dcache_tlb_entries_barrier_io_x_ae_ptw = dcache_tlb__entries_WIRE_ae_ptw;
    assign dcache_tlb_entries_barrier_io_x_ae_final = dcache_tlb__entries_WIRE_ae_final;
    assign dcache_tlb_entries_barrier_io_x_ae_stage2 = dcache_tlb__entries_WIRE_ae_stage2;
    assign dcache_tlb_entries_barrier_io_x_pf = dcache_tlb__entries_WIRE_pf;
    assign dcache_tlb_entries_barrier_io_x_gf = dcache_tlb__entries_WIRE_gf;
    assign dcache_tlb_entries_barrier_io_x_sw = dcache_tlb__entries_WIRE_sw;
    assign dcache_tlb_entries_barrier_io_x_sx = dcache_tlb__entries_WIRE_sx;
    assign dcache_tlb_entries_barrier_io_x_sr = dcache_tlb__entries_WIRE_sr;
    assign dcache_tlb_entries_barrier_io_x_hw = dcache_tlb__entries_WIRE_hw;
    assign dcache_tlb_entries_barrier_io_x_hx = dcache_tlb__entries_WIRE_hx;
    assign dcache_tlb_entries_barrier_io_x_hr = dcache_tlb__entries_WIRE_hr;
    assign dcache_tlb_entries_barrier_io_x_pw = dcache_tlb__entries_WIRE_pw;
    assign dcache_tlb_entries_barrier_io_x_px = dcache_tlb__entries_WIRE_px;
    assign dcache_tlb_entries_barrier_io_x_pr = dcache_tlb__entries_WIRE_pr;
    assign dcache_tlb_entries_barrier_io_x_ppp = dcache_tlb__entries_WIRE_ppp;
    assign dcache_tlb_entries_barrier_io_x_pal = dcache_tlb__entries_WIRE_pal;
    assign dcache_tlb_entries_barrier_io_x_paa = dcache_tlb__entries_WIRE_paa;
    assign dcache_tlb_entries_barrier_io_x_eff = dcache_tlb__entries_WIRE_eff;
    assign dcache_tlb_entries_barrier_io_x_c = dcache_tlb__entries_WIRE_c;
    assign dcache_tlb_entries_barrier_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_fragmented_superpage;
    assign dcache__tlb_entries_barrier_io_y_ppn = dcache_tlb_entries_barrier_io_y_ppn;
    assign dcache__tlb_entries_barrier_io_y_u = dcache_tlb_entries_barrier_io_y_u;
    assign dcache__tlb_entries_barrier_io_y_ae_ptw = dcache_tlb_entries_barrier_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_io_y_ae_final = dcache_tlb_entries_barrier_io_y_ae_final;
    assign dcache__tlb_entries_barrier_io_y_ae_stage2 = dcache_tlb_entries_barrier_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_io_y_pf = dcache_tlb_entries_barrier_io_y_pf;
    assign dcache__tlb_entries_barrier_io_y_gf = dcache_tlb_entries_barrier_io_y_gf;
    assign dcache__tlb_entries_barrier_io_y_sw = dcache_tlb_entries_barrier_io_y_sw;
    assign dcache__tlb_entries_barrier_io_y_sx = dcache_tlb_entries_barrier_io_y_sx;
    assign dcache__tlb_entries_barrier_io_y_sr = dcache_tlb_entries_barrier_io_y_sr;
    assign dcache__tlb_entries_barrier_io_y_hw = dcache_tlb_entries_barrier_io_y_hw;
    assign dcache__tlb_entries_barrier_io_y_hx = dcache_tlb_entries_barrier_io_y_hx;
    assign dcache__tlb_entries_barrier_io_y_hr = dcache_tlb_entries_barrier_io_y_hr;
    assign dcache__tlb_entries_barrier_io_y_pw = dcache_tlb_entries_barrier_io_y_pw;
    assign dcache__tlb_entries_barrier_io_y_px = dcache_tlb_entries_barrier_io_y_px;
    assign dcache__tlb_entries_barrier_io_y_pr = dcache_tlb_entries_barrier_io_y_pr;
    assign dcache__tlb_entries_barrier_io_y_ppp = dcache_tlb_entries_barrier_io_y_ppp;
    assign dcache__tlb_entries_barrier_io_y_pal = dcache_tlb_entries_barrier_io_y_pal;
    assign dcache__tlb_entries_barrier_io_y_paa = dcache_tlb_entries_barrier_io_y_paa;
    assign dcache__tlb_entries_barrier_io_y_eff = dcache_tlb_entries_barrier_io_y_eff;
    assign dcache__tlb_entries_barrier_io_y_c = dcache_tlb_entries_barrier_io_y_c;
    assign dcache_tlb_entries_barrier_1_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_1_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_1_io_x_ppn = dcache_tlb__entries_WIRE_2_ppn;
    assign dcache_tlb_entries_barrier_1_io_x_u = dcache_tlb__entries_WIRE_2_u;
    assign dcache_tlb_entries_barrier_1_io_x_g = dcache_tlb__entries_WIRE_2_g;
    assign dcache_tlb_entries_barrier_1_io_x_ae_ptw = dcache_tlb__entries_WIRE_2_ae_ptw;
    assign dcache_tlb_entries_barrier_1_io_x_ae_final = dcache_tlb__entries_WIRE_2_ae_final;
    assign dcache_tlb_entries_barrier_1_io_x_ae_stage2 = dcache_tlb__entries_WIRE_2_ae_stage2;
    assign dcache_tlb_entries_barrier_1_io_x_pf = dcache_tlb__entries_WIRE_2_pf;
    assign dcache_tlb_entries_barrier_1_io_x_gf = dcache_tlb__entries_WIRE_2_gf;
    assign dcache_tlb_entries_barrier_1_io_x_sw = dcache_tlb__entries_WIRE_2_sw;
    assign dcache_tlb_entries_barrier_1_io_x_sx = dcache_tlb__entries_WIRE_2_sx;
    assign dcache_tlb_entries_barrier_1_io_x_sr = dcache_tlb__entries_WIRE_2_sr;
    assign dcache_tlb_entries_barrier_1_io_x_hw = dcache_tlb__entries_WIRE_2_hw;
    assign dcache_tlb_entries_barrier_1_io_x_hx = dcache_tlb__entries_WIRE_2_hx;
    assign dcache_tlb_entries_barrier_1_io_x_hr = dcache_tlb__entries_WIRE_2_hr;
    assign dcache_tlb_entries_barrier_1_io_x_pw = dcache_tlb__entries_WIRE_2_pw;
    assign dcache_tlb_entries_barrier_1_io_x_px = dcache_tlb__entries_WIRE_2_px;
    assign dcache_tlb_entries_barrier_1_io_x_pr = dcache_tlb__entries_WIRE_2_pr;
    assign dcache_tlb_entries_barrier_1_io_x_ppp = dcache_tlb__entries_WIRE_2_ppp;
    assign dcache_tlb_entries_barrier_1_io_x_pal = dcache_tlb__entries_WIRE_2_pal;
    assign dcache_tlb_entries_barrier_1_io_x_paa = dcache_tlb__entries_WIRE_2_paa;
    assign dcache_tlb_entries_barrier_1_io_x_eff = dcache_tlb__entries_WIRE_2_eff;
    assign dcache_tlb_entries_barrier_1_io_x_c = dcache_tlb__entries_WIRE_2_c;
    assign dcache_tlb_entries_barrier_1_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_2_fragmented_superpage;
    assign dcache__tlb_entries_barrier_1_io_y_ppn = dcache_tlb_entries_barrier_1_io_y_ppn;
    assign dcache__tlb_entries_barrier_1_io_y_u = dcache_tlb_entries_barrier_1_io_y_u;
    assign dcache__tlb_entries_barrier_1_io_y_ae_ptw = dcache_tlb_entries_barrier_1_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_1_io_y_ae_final = dcache_tlb_entries_barrier_1_io_y_ae_final;
    assign dcache__tlb_entries_barrier_1_io_y_ae_stage2 = dcache_tlb_entries_barrier_1_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_1_io_y_pf = dcache_tlb_entries_barrier_1_io_y_pf;
    assign dcache__tlb_entries_barrier_1_io_y_gf = dcache_tlb_entries_barrier_1_io_y_gf;
    assign dcache__tlb_entries_barrier_1_io_y_sw = dcache_tlb_entries_barrier_1_io_y_sw;
    assign dcache__tlb_entries_barrier_1_io_y_sx = dcache_tlb_entries_barrier_1_io_y_sx;
    assign dcache__tlb_entries_barrier_1_io_y_sr = dcache_tlb_entries_barrier_1_io_y_sr;
    assign dcache__tlb_entries_barrier_1_io_y_hw = dcache_tlb_entries_barrier_1_io_y_hw;
    assign dcache__tlb_entries_barrier_1_io_y_hx = dcache_tlb_entries_barrier_1_io_y_hx;
    assign dcache__tlb_entries_barrier_1_io_y_hr = dcache_tlb_entries_barrier_1_io_y_hr;
    assign dcache__tlb_entries_barrier_1_io_y_pw = dcache_tlb_entries_barrier_1_io_y_pw;
    assign dcache__tlb_entries_barrier_1_io_y_px = dcache_tlb_entries_barrier_1_io_y_px;
    assign dcache__tlb_entries_barrier_1_io_y_pr = dcache_tlb_entries_barrier_1_io_y_pr;
    assign dcache__tlb_entries_barrier_1_io_y_ppp = dcache_tlb_entries_barrier_1_io_y_ppp;
    assign dcache__tlb_entries_barrier_1_io_y_pal = dcache_tlb_entries_barrier_1_io_y_pal;
    assign dcache__tlb_entries_barrier_1_io_y_paa = dcache_tlb_entries_barrier_1_io_y_paa;
    assign dcache__tlb_entries_barrier_1_io_y_eff = dcache_tlb_entries_barrier_1_io_y_eff;
    assign dcache__tlb_entries_barrier_1_io_y_c = dcache_tlb_entries_barrier_1_io_y_c;
    assign dcache_tlb_entries_barrier_2_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_2_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_2_io_x_ppn = dcache_tlb__entries_WIRE_4_ppn;
    assign dcache_tlb_entries_barrier_2_io_x_u = dcache_tlb__entries_WIRE_4_u;
    assign dcache_tlb_entries_barrier_2_io_x_g = dcache_tlb__entries_WIRE_4_g;
    assign dcache_tlb_entries_barrier_2_io_x_ae_ptw = dcache_tlb__entries_WIRE_4_ae_ptw;
    assign dcache_tlb_entries_barrier_2_io_x_ae_final = dcache_tlb__entries_WIRE_4_ae_final;
    assign dcache_tlb_entries_barrier_2_io_x_ae_stage2 = dcache_tlb__entries_WIRE_4_ae_stage2;
    assign dcache_tlb_entries_barrier_2_io_x_pf = dcache_tlb__entries_WIRE_4_pf;
    assign dcache_tlb_entries_barrier_2_io_x_gf = dcache_tlb__entries_WIRE_4_gf;
    assign dcache_tlb_entries_barrier_2_io_x_sw = dcache_tlb__entries_WIRE_4_sw;
    assign dcache_tlb_entries_barrier_2_io_x_sx = dcache_tlb__entries_WIRE_4_sx;
    assign dcache_tlb_entries_barrier_2_io_x_sr = dcache_tlb__entries_WIRE_4_sr;
    assign dcache_tlb_entries_barrier_2_io_x_hw = dcache_tlb__entries_WIRE_4_hw;
    assign dcache_tlb_entries_barrier_2_io_x_hx = dcache_tlb__entries_WIRE_4_hx;
    assign dcache_tlb_entries_barrier_2_io_x_hr = dcache_tlb__entries_WIRE_4_hr;
    assign dcache_tlb_entries_barrier_2_io_x_pw = dcache_tlb__entries_WIRE_4_pw;
    assign dcache_tlb_entries_barrier_2_io_x_px = dcache_tlb__entries_WIRE_4_px;
    assign dcache_tlb_entries_barrier_2_io_x_pr = dcache_tlb__entries_WIRE_4_pr;
    assign dcache_tlb_entries_barrier_2_io_x_ppp = dcache_tlb__entries_WIRE_4_ppp;
    assign dcache_tlb_entries_barrier_2_io_x_pal = dcache_tlb__entries_WIRE_4_pal;
    assign dcache_tlb_entries_barrier_2_io_x_paa = dcache_tlb__entries_WIRE_4_paa;
    assign dcache_tlb_entries_barrier_2_io_x_eff = dcache_tlb__entries_WIRE_4_eff;
    assign dcache_tlb_entries_barrier_2_io_x_c = dcache_tlb__entries_WIRE_4_c;
    assign dcache_tlb_entries_barrier_2_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_4_fragmented_superpage;
    assign dcache__tlb_entries_barrier_2_io_y_ppn = dcache_tlb_entries_barrier_2_io_y_ppn;
    assign dcache__tlb_entries_barrier_2_io_y_u = dcache_tlb_entries_barrier_2_io_y_u;
    assign dcache__tlb_entries_barrier_2_io_y_ae_ptw = dcache_tlb_entries_barrier_2_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_2_io_y_ae_final = dcache_tlb_entries_barrier_2_io_y_ae_final;
    assign dcache__tlb_entries_barrier_2_io_y_ae_stage2 = dcache_tlb_entries_barrier_2_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_2_io_y_pf = dcache_tlb_entries_barrier_2_io_y_pf;
    assign dcache__tlb_entries_barrier_2_io_y_gf = dcache_tlb_entries_barrier_2_io_y_gf;
    assign dcache__tlb_entries_barrier_2_io_y_sw = dcache_tlb_entries_barrier_2_io_y_sw;
    assign dcache__tlb_entries_barrier_2_io_y_sx = dcache_tlb_entries_barrier_2_io_y_sx;
    assign dcache__tlb_entries_barrier_2_io_y_sr = dcache_tlb_entries_barrier_2_io_y_sr;
    assign dcache__tlb_entries_barrier_2_io_y_hw = dcache_tlb_entries_barrier_2_io_y_hw;
    assign dcache__tlb_entries_barrier_2_io_y_hx = dcache_tlb_entries_barrier_2_io_y_hx;
    assign dcache__tlb_entries_barrier_2_io_y_hr = dcache_tlb_entries_barrier_2_io_y_hr;
    assign dcache__tlb_entries_barrier_2_io_y_pw = dcache_tlb_entries_barrier_2_io_y_pw;
    assign dcache__tlb_entries_barrier_2_io_y_px = dcache_tlb_entries_barrier_2_io_y_px;
    assign dcache__tlb_entries_barrier_2_io_y_pr = dcache_tlb_entries_barrier_2_io_y_pr;
    assign dcache__tlb_entries_barrier_2_io_y_ppp = dcache_tlb_entries_barrier_2_io_y_ppp;
    assign dcache__tlb_entries_barrier_2_io_y_pal = dcache_tlb_entries_barrier_2_io_y_pal;
    assign dcache__tlb_entries_barrier_2_io_y_paa = dcache_tlb_entries_barrier_2_io_y_paa;
    assign dcache__tlb_entries_barrier_2_io_y_eff = dcache_tlb_entries_barrier_2_io_y_eff;
    assign dcache__tlb_entries_barrier_2_io_y_c = dcache_tlb_entries_barrier_2_io_y_c;
    assign dcache_tlb_entries_barrier_3_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_3_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_3_io_x_ppn = dcache_tlb__entries_WIRE_6_ppn;
    assign dcache_tlb_entries_barrier_3_io_x_u = dcache_tlb__entries_WIRE_6_u;
    assign dcache_tlb_entries_barrier_3_io_x_g = dcache_tlb__entries_WIRE_6_g;
    assign dcache_tlb_entries_barrier_3_io_x_ae_ptw = dcache_tlb__entries_WIRE_6_ae_ptw;
    assign dcache_tlb_entries_barrier_3_io_x_ae_final = dcache_tlb__entries_WIRE_6_ae_final;
    assign dcache_tlb_entries_barrier_3_io_x_ae_stage2 = dcache_tlb__entries_WIRE_6_ae_stage2;
    assign dcache_tlb_entries_barrier_3_io_x_pf = dcache_tlb__entries_WIRE_6_pf;
    assign dcache_tlb_entries_barrier_3_io_x_gf = dcache_tlb__entries_WIRE_6_gf;
    assign dcache_tlb_entries_barrier_3_io_x_sw = dcache_tlb__entries_WIRE_6_sw;
    assign dcache_tlb_entries_barrier_3_io_x_sx = dcache_tlb__entries_WIRE_6_sx;
    assign dcache_tlb_entries_barrier_3_io_x_sr = dcache_tlb__entries_WIRE_6_sr;
    assign dcache_tlb_entries_barrier_3_io_x_hw = dcache_tlb__entries_WIRE_6_hw;
    assign dcache_tlb_entries_barrier_3_io_x_hx = dcache_tlb__entries_WIRE_6_hx;
    assign dcache_tlb_entries_barrier_3_io_x_hr = dcache_tlb__entries_WIRE_6_hr;
    assign dcache_tlb_entries_barrier_3_io_x_pw = dcache_tlb__entries_WIRE_6_pw;
    assign dcache_tlb_entries_barrier_3_io_x_px = dcache_tlb__entries_WIRE_6_px;
    assign dcache_tlb_entries_barrier_3_io_x_pr = dcache_tlb__entries_WIRE_6_pr;
    assign dcache_tlb_entries_barrier_3_io_x_ppp = dcache_tlb__entries_WIRE_6_ppp;
    assign dcache_tlb_entries_barrier_3_io_x_pal = dcache_tlb__entries_WIRE_6_pal;
    assign dcache_tlb_entries_barrier_3_io_x_paa = dcache_tlb__entries_WIRE_6_paa;
    assign dcache_tlb_entries_barrier_3_io_x_eff = dcache_tlb__entries_WIRE_6_eff;
    assign dcache_tlb_entries_barrier_3_io_x_c = dcache_tlb__entries_WIRE_6_c;
    assign dcache_tlb_entries_barrier_3_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_6_fragmented_superpage;
    assign dcache__tlb_entries_barrier_3_io_y_ppn = dcache_tlb_entries_barrier_3_io_y_ppn;
    assign dcache__tlb_entries_barrier_3_io_y_u = dcache_tlb_entries_barrier_3_io_y_u;
    assign dcache__tlb_entries_barrier_3_io_y_ae_ptw = dcache_tlb_entries_barrier_3_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_3_io_y_ae_final = dcache_tlb_entries_barrier_3_io_y_ae_final;
    assign dcache__tlb_entries_barrier_3_io_y_ae_stage2 = dcache_tlb_entries_barrier_3_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_3_io_y_pf = dcache_tlb_entries_barrier_3_io_y_pf;
    assign dcache__tlb_entries_barrier_3_io_y_gf = dcache_tlb_entries_barrier_3_io_y_gf;
    assign dcache__tlb_entries_barrier_3_io_y_sw = dcache_tlb_entries_barrier_3_io_y_sw;
    assign dcache__tlb_entries_barrier_3_io_y_sx = dcache_tlb_entries_barrier_3_io_y_sx;
    assign dcache__tlb_entries_barrier_3_io_y_sr = dcache_tlb_entries_barrier_3_io_y_sr;
    assign dcache__tlb_entries_barrier_3_io_y_hw = dcache_tlb_entries_barrier_3_io_y_hw;
    assign dcache__tlb_entries_barrier_3_io_y_hx = dcache_tlb_entries_barrier_3_io_y_hx;
    assign dcache__tlb_entries_barrier_3_io_y_hr = dcache_tlb_entries_barrier_3_io_y_hr;
    assign dcache__tlb_entries_barrier_3_io_y_pw = dcache_tlb_entries_barrier_3_io_y_pw;
    assign dcache__tlb_entries_barrier_3_io_y_px = dcache_tlb_entries_barrier_3_io_y_px;
    assign dcache__tlb_entries_barrier_3_io_y_pr = dcache_tlb_entries_barrier_3_io_y_pr;
    assign dcache__tlb_entries_barrier_3_io_y_ppp = dcache_tlb_entries_barrier_3_io_y_ppp;
    assign dcache__tlb_entries_barrier_3_io_y_pal = dcache_tlb_entries_barrier_3_io_y_pal;
    assign dcache__tlb_entries_barrier_3_io_y_paa = dcache_tlb_entries_barrier_3_io_y_paa;
    assign dcache__tlb_entries_barrier_3_io_y_eff = dcache_tlb_entries_barrier_3_io_y_eff;
    assign dcache__tlb_entries_barrier_3_io_y_c = dcache_tlb_entries_barrier_3_io_y_c;
    assign dcache_tlb_entries_barrier_4_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_4_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_4_io_x_ppn = dcache_tlb__entries_WIRE_8_ppn;
    assign dcache_tlb_entries_barrier_4_io_x_u = dcache_tlb__entries_WIRE_8_u;
    assign dcache_tlb_entries_barrier_4_io_x_g = dcache_tlb__entries_WIRE_8_g;
    assign dcache_tlb_entries_barrier_4_io_x_ae_ptw = dcache_tlb__entries_WIRE_8_ae_ptw;
    assign dcache_tlb_entries_barrier_4_io_x_ae_final = dcache_tlb__entries_WIRE_8_ae_final;
    assign dcache_tlb_entries_barrier_4_io_x_ae_stage2 = dcache_tlb__entries_WIRE_8_ae_stage2;
    assign dcache_tlb_entries_barrier_4_io_x_pf = dcache_tlb__entries_WIRE_8_pf;
    assign dcache_tlb_entries_barrier_4_io_x_gf = dcache_tlb__entries_WIRE_8_gf;
    assign dcache_tlb_entries_barrier_4_io_x_sw = dcache_tlb__entries_WIRE_8_sw;
    assign dcache_tlb_entries_barrier_4_io_x_sx = dcache_tlb__entries_WIRE_8_sx;
    assign dcache_tlb_entries_barrier_4_io_x_sr = dcache_tlb__entries_WIRE_8_sr;
    assign dcache_tlb_entries_barrier_4_io_x_hw = dcache_tlb__entries_WIRE_8_hw;
    assign dcache_tlb_entries_barrier_4_io_x_hx = dcache_tlb__entries_WIRE_8_hx;
    assign dcache_tlb_entries_barrier_4_io_x_hr = dcache_tlb__entries_WIRE_8_hr;
    assign dcache_tlb_entries_barrier_4_io_x_pw = dcache_tlb__entries_WIRE_8_pw;
    assign dcache_tlb_entries_barrier_4_io_x_px = dcache_tlb__entries_WIRE_8_px;
    assign dcache_tlb_entries_barrier_4_io_x_pr = dcache_tlb__entries_WIRE_8_pr;
    assign dcache_tlb_entries_barrier_4_io_x_ppp = dcache_tlb__entries_WIRE_8_ppp;
    assign dcache_tlb_entries_barrier_4_io_x_pal = dcache_tlb__entries_WIRE_8_pal;
    assign dcache_tlb_entries_barrier_4_io_x_paa = dcache_tlb__entries_WIRE_8_paa;
    assign dcache_tlb_entries_barrier_4_io_x_eff = dcache_tlb__entries_WIRE_8_eff;
    assign dcache_tlb_entries_barrier_4_io_x_c = dcache_tlb__entries_WIRE_8_c;
    assign dcache_tlb_entries_barrier_4_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_8_fragmented_superpage;
    assign dcache__tlb_entries_barrier_4_io_y_ppn = dcache_tlb_entries_barrier_4_io_y_ppn;
    assign dcache__tlb_entries_barrier_4_io_y_u = dcache_tlb_entries_barrier_4_io_y_u;
    assign dcache__tlb_entries_barrier_4_io_y_ae_ptw = dcache_tlb_entries_barrier_4_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_4_io_y_ae_final = dcache_tlb_entries_barrier_4_io_y_ae_final;
    assign dcache__tlb_entries_barrier_4_io_y_ae_stage2 = dcache_tlb_entries_barrier_4_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_4_io_y_pf = dcache_tlb_entries_barrier_4_io_y_pf;
    assign dcache__tlb_entries_barrier_4_io_y_gf = dcache_tlb_entries_barrier_4_io_y_gf;
    assign dcache__tlb_entries_barrier_4_io_y_sw = dcache_tlb_entries_barrier_4_io_y_sw;
    assign dcache__tlb_entries_barrier_4_io_y_sx = dcache_tlb_entries_barrier_4_io_y_sx;
    assign dcache__tlb_entries_barrier_4_io_y_sr = dcache_tlb_entries_barrier_4_io_y_sr;
    assign dcache__tlb_entries_barrier_4_io_y_hw = dcache_tlb_entries_barrier_4_io_y_hw;
    assign dcache__tlb_entries_barrier_4_io_y_hx = dcache_tlb_entries_barrier_4_io_y_hx;
    assign dcache__tlb_entries_barrier_4_io_y_hr = dcache_tlb_entries_barrier_4_io_y_hr;
    assign dcache__tlb_entries_barrier_4_io_y_pw = dcache_tlb_entries_barrier_4_io_y_pw;
    assign dcache__tlb_entries_barrier_4_io_y_px = dcache_tlb_entries_barrier_4_io_y_px;
    assign dcache__tlb_entries_barrier_4_io_y_pr = dcache_tlb_entries_barrier_4_io_y_pr;
    assign dcache__tlb_entries_barrier_4_io_y_ppp = dcache_tlb_entries_barrier_4_io_y_ppp;
    assign dcache__tlb_entries_barrier_4_io_y_pal = dcache_tlb_entries_barrier_4_io_y_pal;
    assign dcache__tlb_entries_barrier_4_io_y_paa = dcache_tlb_entries_barrier_4_io_y_paa;
    assign dcache__tlb_entries_barrier_4_io_y_eff = dcache_tlb_entries_barrier_4_io_y_eff;
    assign dcache__tlb_entries_barrier_4_io_y_c = dcache_tlb_entries_barrier_4_io_y_c;
    assign dcache_tlb_entries_barrier_5_clock = dcache_tlb_clock;
    assign dcache_tlb_entries_barrier_5_reset = dcache_tlb_reset;
    assign dcache_tlb_entries_barrier_5_io_x_ppn = dcache_tlb__entries_WIRE_10_ppn;
    assign dcache_tlb_entries_barrier_5_io_x_u = dcache_tlb__entries_WIRE_10_u;
    assign dcache_tlb_entries_barrier_5_io_x_g = dcache_tlb__entries_WIRE_10_g;
    assign dcache_tlb_entries_barrier_5_io_x_ae_ptw = dcache_tlb__entries_WIRE_10_ae_ptw;
    assign dcache_tlb_entries_barrier_5_io_x_ae_final = dcache_tlb__entries_WIRE_10_ae_final;
    assign dcache_tlb_entries_barrier_5_io_x_ae_stage2 = dcache_tlb__entries_WIRE_10_ae_stage2;
    assign dcache_tlb_entries_barrier_5_io_x_pf = dcache_tlb__entries_WIRE_10_pf;
    assign dcache_tlb_entries_barrier_5_io_x_gf = dcache_tlb__entries_WIRE_10_gf;
    assign dcache_tlb_entries_barrier_5_io_x_sw = dcache_tlb__entries_WIRE_10_sw;
    assign dcache_tlb_entries_barrier_5_io_x_sx = dcache_tlb__entries_WIRE_10_sx;
    assign dcache_tlb_entries_barrier_5_io_x_sr = dcache_tlb__entries_WIRE_10_sr;
    assign dcache_tlb_entries_barrier_5_io_x_hw = dcache_tlb__entries_WIRE_10_hw;
    assign dcache_tlb_entries_barrier_5_io_x_hx = dcache_tlb__entries_WIRE_10_hx;
    assign dcache_tlb_entries_barrier_5_io_x_hr = dcache_tlb__entries_WIRE_10_hr;
    assign dcache_tlb_entries_barrier_5_io_x_pw = dcache_tlb__entries_WIRE_10_pw;
    assign dcache_tlb_entries_barrier_5_io_x_px = dcache_tlb__entries_WIRE_10_px;
    assign dcache_tlb_entries_barrier_5_io_x_pr = dcache_tlb__entries_WIRE_10_pr;
    assign dcache_tlb_entries_barrier_5_io_x_ppp = dcache_tlb__entries_WIRE_10_ppp;
    assign dcache_tlb_entries_barrier_5_io_x_pal = dcache_tlb__entries_WIRE_10_pal;
    assign dcache_tlb_entries_barrier_5_io_x_paa = dcache_tlb__entries_WIRE_10_paa;
    assign dcache_tlb_entries_barrier_5_io_x_eff = dcache_tlb__entries_WIRE_10_eff;
    assign dcache_tlb_entries_barrier_5_io_x_c = dcache_tlb__entries_WIRE_10_c;
    assign dcache_tlb_entries_barrier_5_io_x_fragmented_superpage = dcache_tlb__entries_WIRE_10_fragmented_superpage;
    assign dcache__tlb_entries_barrier_5_io_y_ppn = dcache_tlb_entries_barrier_5_io_y_ppn;
    assign dcache__tlb_entries_barrier_5_io_y_u = dcache_tlb_entries_barrier_5_io_y_u;
    assign dcache__tlb_entries_barrier_5_io_y_ae_ptw = dcache_tlb_entries_barrier_5_io_y_ae_ptw;
    assign dcache__tlb_entries_barrier_5_io_y_ae_final = dcache_tlb_entries_barrier_5_io_y_ae_final;
    assign dcache__tlb_entries_barrier_5_io_y_ae_stage2 = dcache_tlb_entries_barrier_5_io_y_ae_stage2;
    assign dcache__tlb_entries_barrier_5_io_y_pf = dcache_tlb_entries_barrier_5_io_y_pf;
    assign dcache__tlb_entries_barrier_5_io_y_gf = dcache_tlb_entries_barrier_5_io_y_gf;
    assign dcache__tlb_entries_barrier_5_io_y_sw = dcache_tlb_entries_barrier_5_io_y_sw;
    assign dcache__tlb_entries_barrier_5_io_y_sx = dcache_tlb_entries_barrier_5_io_y_sx;
    assign dcache__tlb_entries_barrier_5_io_y_sr = dcache_tlb_entries_barrier_5_io_y_sr;
    assign dcache__tlb_entries_barrier_5_io_y_hw = dcache_tlb_entries_barrier_5_io_y_hw;
    assign dcache__tlb_entries_barrier_5_io_y_hx = dcache_tlb_entries_barrier_5_io_y_hx;
    assign dcache__tlb_entries_barrier_5_io_y_hr = dcache_tlb_entries_barrier_5_io_y_hr;
    assign dcache_pma_checker_mpu_ppn_barrier_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_mpu_ppn_barrier_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_ppn = dcache_pma_checker__mpu_ppn_WIRE_ppn;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_u = dcache_pma_checker__mpu_ppn_WIRE_u;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_g = dcache_pma_checker__mpu_ppn_WIRE_g;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_ae_ptw = dcache_pma_checker__mpu_ppn_WIRE_ae_ptw;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_ae_final = dcache_pma_checker__mpu_ppn_WIRE_ae_final;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_ae_stage2 = dcache_pma_checker__mpu_ppn_WIRE_ae_stage2;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_pf = dcache_pma_checker__mpu_ppn_WIRE_pf;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_gf = dcache_pma_checker__mpu_ppn_WIRE_gf;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_sw = dcache_pma_checker__mpu_ppn_WIRE_sw;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_sx = dcache_pma_checker__mpu_ppn_WIRE_sx;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_sr = dcache_pma_checker__mpu_ppn_WIRE_sr;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_hw = dcache_pma_checker__mpu_ppn_WIRE_hw;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_hx = dcache_pma_checker__mpu_ppn_WIRE_hx;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_hr = dcache_pma_checker__mpu_ppn_WIRE_hr;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_pw = dcache_pma_checker__mpu_ppn_WIRE_pw;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_px = dcache_pma_checker__mpu_ppn_WIRE_px;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_pr = dcache_pma_checker__mpu_ppn_WIRE_pr;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_ppp = dcache_pma_checker__mpu_ppn_WIRE_ppp;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_pal = dcache_pma_checker__mpu_ppn_WIRE_pal;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_paa = dcache_pma_checker__mpu_ppn_WIRE_paa;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_eff = dcache_pma_checker__mpu_ppn_WIRE_eff;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_c = dcache_pma_checker__mpu_ppn_WIRE_c;
    assign dcache_pma_checker_mpu_ppn_barrier_io_x_fragmented_superpage = dcache_pma_checker__mpu_ppn_WIRE_fragmented_superpage;
    assign dcache__pma_checker_mpu_ppn_barrier_io_y_ppn = dcache_pma_checker_mpu_ppn_barrier_io_y_ppn;
    assign dcache_pma_checker_entries_barrier_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_io_x_ppn = dcache_pma_checker__entries_WIRE_ppn;
    assign dcache_pma_checker_entries_barrier_io_x_u = dcache_pma_checker__entries_WIRE_u;
    assign dcache_pma_checker_entries_barrier_io_x_g = dcache_pma_checker__entries_WIRE_g;
    assign dcache_pma_checker_entries_barrier_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_ae_ptw;
    assign dcache_pma_checker_entries_barrier_io_x_ae_final = dcache_pma_checker__entries_WIRE_ae_final;
    assign dcache_pma_checker_entries_barrier_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_ae_stage2;
    assign dcache_pma_checker_entries_barrier_io_x_pf = dcache_pma_checker__entries_WIRE_pf;
    assign dcache_pma_checker_entries_barrier_io_x_gf = dcache_pma_checker__entries_WIRE_gf;
    assign dcache_pma_checker_entries_barrier_io_x_sw = dcache_pma_checker__entries_WIRE_sw;
    assign dcache_pma_checker_entries_barrier_io_x_sx = dcache_pma_checker__entries_WIRE_sx;
    assign dcache_pma_checker_entries_barrier_io_x_sr = dcache_pma_checker__entries_WIRE_sr;
    assign dcache_pma_checker_entries_barrier_io_x_hw = dcache_pma_checker__entries_WIRE_hw;
    assign dcache_pma_checker_entries_barrier_io_x_hx = dcache_pma_checker__entries_WIRE_hx;
    assign dcache_pma_checker_entries_barrier_io_x_hr = dcache_pma_checker__entries_WIRE_hr;
    assign dcache_pma_checker_entries_barrier_io_x_pw = dcache_pma_checker__entries_WIRE_pw;
    assign dcache_pma_checker_entries_barrier_io_x_px = dcache_pma_checker__entries_WIRE_px;
    assign dcache_pma_checker_entries_barrier_io_x_pr = dcache_pma_checker__entries_WIRE_pr;
    assign dcache_pma_checker_entries_barrier_io_x_ppp = dcache_pma_checker__entries_WIRE_ppp;
    assign dcache_pma_checker_entries_barrier_io_x_pal = dcache_pma_checker__entries_WIRE_pal;
    assign dcache_pma_checker_entries_barrier_io_x_paa = dcache_pma_checker__entries_WIRE_paa;
    assign dcache_pma_checker_entries_barrier_io_x_eff = dcache_pma_checker__entries_WIRE_eff;
    assign dcache_pma_checker_entries_barrier_io_x_c = dcache_pma_checker__entries_WIRE_c;
    assign dcache_pma_checker_entries_barrier_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_io_y_ppn = dcache_pma_checker_entries_barrier_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_io_y_u = dcache_pma_checker_entries_barrier_io_y_u;
    assign dcache__pma_checker_entries_barrier_io_y_ae_ptw = dcache_pma_checker_entries_barrier_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_io_y_ae_final = dcache_pma_checker_entries_barrier_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_io_y_pf = dcache_pma_checker_entries_barrier_io_y_pf;
    assign dcache__pma_checker_entries_barrier_io_y_gf = dcache_pma_checker_entries_barrier_io_y_gf;
    assign dcache__pma_checker_entries_barrier_io_y_sw = dcache_pma_checker_entries_barrier_io_y_sw;
    assign dcache__pma_checker_entries_barrier_io_y_sx = dcache_pma_checker_entries_barrier_io_y_sx;
    assign dcache__pma_checker_entries_barrier_io_y_sr = dcache_pma_checker_entries_barrier_io_y_sr;
    assign dcache__pma_checker_entries_barrier_io_y_hw = dcache_pma_checker_entries_barrier_io_y_hw;
    assign dcache__pma_checker_entries_barrier_io_y_hx = dcache_pma_checker_entries_barrier_io_y_hx;
    assign dcache__pma_checker_entries_barrier_io_y_hr = dcache_pma_checker_entries_barrier_io_y_hr;
    assign dcache__pma_checker_entries_barrier_io_y_pw = dcache_pma_checker_entries_barrier_io_y_pw;
    assign dcache__pma_checker_entries_barrier_io_y_px = dcache_pma_checker_entries_barrier_io_y_px;
    assign dcache__pma_checker_entries_barrier_io_y_pr = dcache_pma_checker_entries_barrier_io_y_pr;
    assign dcache__pma_checker_entries_barrier_io_y_ppp = dcache_pma_checker_entries_barrier_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_io_y_pal = dcache_pma_checker_entries_barrier_io_y_pal;
    assign dcache__pma_checker_entries_barrier_io_y_paa = dcache_pma_checker_entries_barrier_io_y_paa;
    assign dcache__pma_checker_entries_barrier_io_y_eff = dcache_pma_checker_entries_barrier_io_y_eff;
    assign dcache__pma_checker_entries_barrier_io_y_c = dcache_pma_checker_entries_barrier_io_y_c;
    assign dcache_pma_checker_entries_barrier_1_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_1_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_1_io_x_ppn = dcache_pma_checker__entries_WIRE_2_ppn;
    assign dcache_pma_checker_entries_barrier_1_io_x_u = dcache_pma_checker__entries_WIRE_2_u;
    assign dcache_pma_checker_entries_barrier_1_io_x_g = dcache_pma_checker__entries_WIRE_2_g;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_2_ae_ptw;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_final = dcache_pma_checker__entries_WIRE_2_ae_final;
    assign dcache_pma_checker_entries_barrier_1_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_2_ae_stage2;
    assign dcache_pma_checker_entries_barrier_1_io_x_pf = dcache_pma_checker__entries_WIRE_2_pf;
    assign dcache_pma_checker_entries_barrier_1_io_x_gf = dcache_pma_checker__entries_WIRE_2_gf;
    assign dcache_pma_checker_entries_barrier_1_io_x_sw = dcache_pma_checker__entries_WIRE_2_sw;
    assign dcache_pma_checker_entries_barrier_1_io_x_sx = dcache_pma_checker__entries_WIRE_2_sx;
    assign dcache_pma_checker_entries_barrier_1_io_x_sr = dcache_pma_checker__entries_WIRE_2_sr;
    assign dcache_pma_checker_entries_barrier_1_io_x_hw = dcache_pma_checker__entries_WIRE_2_hw;
    assign dcache_pma_checker_entries_barrier_1_io_x_hx = dcache_pma_checker__entries_WIRE_2_hx;
    assign dcache_pma_checker_entries_barrier_1_io_x_hr = dcache_pma_checker__entries_WIRE_2_hr;
    assign dcache_pma_checker_entries_barrier_1_io_x_pw = dcache_pma_checker__entries_WIRE_2_pw;
    assign dcache_pma_checker_entries_barrier_1_io_x_px = dcache_pma_checker__entries_WIRE_2_px;
    assign dcache_pma_checker_entries_barrier_1_io_x_pr = dcache_pma_checker__entries_WIRE_2_pr;
    assign dcache_pma_checker_entries_barrier_1_io_x_ppp = dcache_pma_checker__entries_WIRE_2_ppp;
    assign dcache_pma_checker_entries_barrier_1_io_x_pal = dcache_pma_checker__entries_WIRE_2_pal;
    assign dcache_pma_checker_entries_barrier_1_io_x_paa = dcache_pma_checker__entries_WIRE_2_paa;
    assign dcache_pma_checker_entries_barrier_1_io_x_eff = dcache_pma_checker__entries_WIRE_2_eff;
    assign dcache_pma_checker_entries_barrier_1_io_x_c = dcache_pma_checker__entries_WIRE_2_c;
    assign dcache_pma_checker_entries_barrier_1_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_2_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_1_io_y_ppn = dcache_pma_checker_entries_barrier_1_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_1_io_y_u = dcache_pma_checker_entries_barrier_1_io_y_u;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_ptw = dcache_pma_checker_entries_barrier_1_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_final = dcache_pma_checker_entries_barrier_1_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_1_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_1_io_y_pf = dcache_pma_checker_entries_barrier_1_io_y_pf;
    assign dcache__pma_checker_entries_barrier_1_io_y_gf = dcache_pma_checker_entries_barrier_1_io_y_gf;
    assign dcache__pma_checker_entries_barrier_1_io_y_sw = dcache_pma_checker_entries_barrier_1_io_y_sw;
    assign dcache__pma_checker_entries_barrier_1_io_y_sx = dcache_pma_checker_entries_barrier_1_io_y_sx;
    assign dcache__pma_checker_entries_barrier_1_io_y_sr = dcache_pma_checker_entries_barrier_1_io_y_sr;
    assign dcache__pma_checker_entries_barrier_1_io_y_hw = dcache_pma_checker_entries_barrier_1_io_y_hw;
    assign dcache__pma_checker_entries_barrier_1_io_y_hx = dcache_pma_checker_entries_barrier_1_io_y_hx;
    assign dcache__pma_checker_entries_barrier_1_io_y_hr = dcache_pma_checker_entries_barrier_1_io_y_hr;
    assign dcache__pma_checker_entries_barrier_1_io_y_pw = dcache_pma_checker_entries_barrier_1_io_y_pw;
    assign dcache__pma_checker_entries_barrier_1_io_y_px = dcache_pma_checker_entries_barrier_1_io_y_px;
    assign dcache__pma_checker_entries_barrier_1_io_y_pr = dcache_pma_checker_entries_barrier_1_io_y_pr;
    assign dcache__pma_checker_entries_barrier_1_io_y_ppp = dcache_pma_checker_entries_barrier_1_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_1_io_y_pal = dcache_pma_checker_entries_barrier_1_io_y_pal;
    assign dcache__pma_checker_entries_barrier_1_io_y_paa = dcache_pma_checker_entries_barrier_1_io_y_paa;
    assign dcache__pma_checker_entries_barrier_1_io_y_eff = dcache_pma_checker_entries_barrier_1_io_y_eff;
    assign dcache__pma_checker_entries_barrier_1_io_y_c = dcache_pma_checker_entries_barrier_1_io_y_c;
    assign dcache_pma_checker_entries_barrier_2_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_2_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_2_io_x_ppn = dcache_pma_checker__entries_WIRE_4_ppn;
    assign dcache_pma_checker_entries_barrier_2_io_x_u = dcache_pma_checker__entries_WIRE_4_u;
    assign dcache_pma_checker_entries_barrier_2_io_x_g = dcache_pma_checker__entries_WIRE_4_g;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_4_ae_ptw;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_final = dcache_pma_checker__entries_WIRE_4_ae_final;
    assign dcache_pma_checker_entries_barrier_2_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_4_ae_stage2;
    assign dcache_pma_checker_entries_barrier_2_io_x_pf = dcache_pma_checker__entries_WIRE_4_pf;
    assign dcache_pma_checker_entries_barrier_2_io_x_gf = dcache_pma_checker__entries_WIRE_4_gf;
    assign dcache_pma_checker_entries_barrier_2_io_x_sw = dcache_pma_checker__entries_WIRE_4_sw;
    assign dcache_pma_checker_entries_barrier_2_io_x_sx = dcache_pma_checker__entries_WIRE_4_sx;
    assign dcache_pma_checker_entries_barrier_2_io_x_sr = dcache_pma_checker__entries_WIRE_4_sr;
    assign dcache_pma_checker_entries_barrier_2_io_x_hw = dcache_pma_checker__entries_WIRE_4_hw;
    assign dcache_pma_checker_entries_barrier_2_io_x_hx = dcache_pma_checker__entries_WIRE_4_hx;
    assign dcache_pma_checker_entries_barrier_2_io_x_hr = dcache_pma_checker__entries_WIRE_4_hr;
    assign dcache_pma_checker_entries_barrier_2_io_x_pw = dcache_pma_checker__entries_WIRE_4_pw;
    assign dcache_pma_checker_entries_barrier_2_io_x_px = dcache_pma_checker__entries_WIRE_4_px;
    assign dcache_pma_checker_entries_barrier_2_io_x_pr = dcache_pma_checker__entries_WIRE_4_pr;
    assign dcache_pma_checker_entries_barrier_2_io_x_ppp = dcache_pma_checker__entries_WIRE_4_ppp;
    assign dcache_pma_checker_entries_barrier_2_io_x_pal = dcache_pma_checker__entries_WIRE_4_pal;
    assign dcache_pma_checker_entries_barrier_2_io_x_paa = dcache_pma_checker__entries_WIRE_4_paa;
    assign dcache_pma_checker_entries_barrier_2_io_x_eff = dcache_pma_checker__entries_WIRE_4_eff;
    assign dcache_pma_checker_entries_barrier_2_io_x_c = dcache_pma_checker__entries_WIRE_4_c;
    assign dcache_pma_checker_entries_barrier_2_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_4_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_2_io_y_ppn = dcache_pma_checker_entries_barrier_2_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_2_io_y_u = dcache_pma_checker_entries_barrier_2_io_y_u;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_ptw = dcache_pma_checker_entries_barrier_2_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_final = dcache_pma_checker_entries_barrier_2_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_2_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_2_io_y_pf = dcache_pma_checker_entries_barrier_2_io_y_pf;
    assign dcache__pma_checker_entries_barrier_2_io_y_gf = dcache_pma_checker_entries_barrier_2_io_y_gf;
    assign dcache__pma_checker_entries_barrier_2_io_y_sw = dcache_pma_checker_entries_barrier_2_io_y_sw;
    assign dcache__pma_checker_entries_barrier_2_io_y_sx = dcache_pma_checker_entries_barrier_2_io_y_sx;
    assign dcache__pma_checker_entries_barrier_2_io_y_sr = dcache_pma_checker_entries_barrier_2_io_y_sr;
    assign dcache__pma_checker_entries_barrier_2_io_y_hw = dcache_pma_checker_entries_barrier_2_io_y_hw;
    assign dcache__pma_checker_entries_barrier_2_io_y_hx = dcache_pma_checker_entries_barrier_2_io_y_hx;
    assign dcache__pma_checker_entries_barrier_2_io_y_hr = dcache_pma_checker_entries_barrier_2_io_y_hr;
    assign dcache__pma_checker_entries_barrier_2_io_y_pw = dcache_pma_checker_entries_barrier_2_io_y_pw;
    assign dcache__pma_checker_entries_barrier_2_io_y_px = dcache_pma_checker_entries_barrier_2_io_y_px;
    assign dcache__pma_checker_entries_barrier_2_io_y_pr = dcache_pma_checker_entries_barrier_2_io_y_pr;
    assign dcache__pma_checker_entries_barrier_2_io_y_ppp = dcache_pma_checker_entries_barrier_2_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_2_io_y_pal = dcache_pma_checker_entries_barrier_2_io_y_pal;
    assign dcache__pma_checker_entries_barrier_2_io_y_paa = dcache_pma_checker_entries_barrier_2_io_y_paa;
    assign dcache__pma_checker_entries_barrier_2_io_y_eff = dcache_pma_checker_entries_barrier_2_io_y_eff;
    assign dcache__pma_checker_entries_barrier_2_io_y_c = dcache_pma_checker_entries_barrier_2_io_y_c;
    assign dcache_pma_checker_entries_barrier_3_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_3_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_3_io_x_ppn = dcache_pma_checker__entries_WIRE_6_ppn;
    assign dcache_pma_checker_entries_barrier_3_io_x_u = dcache_pma_checker__entries_WIRE_6_u;
    assign dcache_pma_checker_entries_barrier_3_io_x_g = dcache_pma_checker__entries_WIRE_6_g;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_6_ae_ptw;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_final = dcache_pma_checker__entries_WIRE_6_ae_final;
    assign dcache_pma_checker_entries_barrier_3_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_6_ae_stage2;
    assign dcache_pma_checker_entries_barrier_3_io_x_pf = dcache_pma_checker__entries_WIRE_6_pf;
    assign dcache_pma_checker_entries_barrier_3_io_x_gf = dcache_pma_checker__entries_WIRE_6_gf;
    assign dcache_pma_checker_entries_barrier_3_io_x_sw = dcache_pma_checker__entries_WIRE_6_sw;
    assign dcache_pma_checker_entries_barrier_3_io_x_sx = dcache_pma_checker__entries_WIRE_6_sx;
    assign dcache_pma_checker_entries_barrier_3_io_x_sr = dcache_pma_checker__entries_WIRE_6_sr;
    assign dcache_pma_checker_entries_barrier_3_io_x_hw = dcache_pma_checker__entries_WIRE_6_hw;
    assign dcache_pma_checker_entries_barrier_3_io_x_hx = dcache_pma_checker__entries_WIRE_6_hx;
    assign dcache_pma_checker_entries_barrier_3_io_x_hr = dcache_pma_checker__entries_WIRE_6_hr;
    assign dcache_pma_checker_entries_barrier_3_io_x_pw = dcache_pma_checker__entries_WIRE_6_pw;
    assign dcache_pma_checker_entries_barrier_3_io_x_px = dcache_pma_checker__entries_WIRE_6_px;
    assign dcache_pma_checker_entries_barrier_3_io_x_pr = dcache_pma_checker__entries_WIRE_6_pr;
    assign dcache_pma_checker_entries_barrier_3_io_x_ppp = dcache_pma_checker__entries_WIRE_6_ppp;
    assign dcache_pma_checker_entries_barrier_3_io_x_pal = dcache_pma_checker__entries_WIRE_6_pal;
    assign dcache_pma_checker_entries_barrier_3_io_x_paa = dcache_pma_checker__entries_WIRE_6_paa;
    assign dcache_pma_checker_entries_barrier_3_io_x_eff = dcache_pma_checker__entries_WIRE_6_eff;
    assign dcache_pma_checker_entries_barrier_3_io_x_c = dcache_pma_checker__entries_WIRE_6_c;
    assign dcache_pma_checker_entries_barrier_3_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_6_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_3_io_y_ppn = dcache_pma_checker_entries_barrier_3_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_3_io_y_u = dcache_pma_checker_entries_barrier_3_io_y_u;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_ptw = dcache_pma_checker_entries_barrier_3_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_final = dcache_pma_checker_entries_barrier_3_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_3_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_3_io_y_pf = dcache_pma_checker_entries_barrier_3_io_y_pf;
    assign dcache__pma_checker_entries_barrier_3_io_y_gf = dcache_pma_checker_entries_barrier_3_io_y_gf;
    assign dcache__pma_checker_entries_barrier_3_io_y_sw = dcache_pma_checker_entries_barrier_3_io_y_sw;
    assign dcache__pma_checker_entries_barrier_3_io_y_sx = dcache_pma_checker_entries_barrier_3_io_y_sx;
    assign dcache__pma_checker_entries_barrier_3_io_y_sr = dcache_pma_checker_entries_barrier_3_io_y_sr;
    assign dcache__pma_checker_entries_barrier_3_io_y_hw = dcache_pma_checker_entries_barrier_3_io_y_hw;
    assign dcache__pma_checker_entries_barrier_3_io_y_hx = dcache_pma_checker_entries_barrier_3_io_y_hx;
    assign dcache__pma_checker_entries_barrier_3_io_y_hr = dcache_pma_checker_entries_barrier_3_io_y_hr;
    assign dcache__pma_checker_entries_barrier_3_io_y_pw = dcache_pma_checker_entries_barrier_3_io_y_pw;
    assign dcache__pma_checker_entries_barrier_3_io_y_px = dcache_pma_checker_entries_barrier_3_io_y_px;
    assign dcache__pma_checker_entries_barrier_3_io_y_pr = dcache_pma_checker_entries_barrier_3_io_y_pr;
    assign dcache__pma_checker_entries_barrier_3_io_y_ppp = dcache_pma_checker_entries_barrier_3_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_3_io_y_pal = dcache_pma_checker_entries_barrier_3_io_y_pal;
    assign dcache__pma_checker_entries_barrier_3_io_y_paa = dcache_pma_checker_entries_barrier_3_io_y_paa;
    assign dcache__pma_checker_entries_barrier_3_io_y_eff = dcache_pma_checker_entries_barrier_3_io_y_eff;
    assign dcache__pma_checker_entries_barrier_3_io_y_c = dcache_pma_checker_entries_barrier_3_io_y_c;
    assign dcache_pma_checker_entries_barrier_4_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_4_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_4_io_x_ppn = dcache_pma_checker__entries_WIRE_8_ppn;
    assign dcache_pma_checker_entries_barrier_4_io_x_u = dcache_pma_checker__entries_WIRE_8_u;
    assign dcache_pma_checker_entries_barrier_4_io_x_g = dcache_pma_checker__entries_WIRE_8_g;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_8_ae_ptw;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_final = dcache_pma_checker__entries_WIRE_8_ae_final;
    assign dcache_pma_checker_entries_barrier_4_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_8_ae_stage2;
    assign dcache_pma_checker_entries_barrier_4_io_x_pf = dcache_pma_checker__entries_WIRE_8_pf;
    assign dcache_pma_checker_entries_barrier_4_io_x_gf = dcache_pma_checker__entries_WIRE_8_gf;
    assign dcache_pma_checker_entries_barrier_4_io_x_sw = dcache_pma_checker__entries_WIRE_8_sw;
    assign dcache_pma_checker_entries_barrier_4_io_x_sx = dcache_pma_checker__entries_WIRE_8_sx;
    assign dcache_pma_checker_entries_barrier_4_io_x_sr = dcache_pma_checker__entries_WIRE_8_sr;
    assign dcache_pma_checker_entries_barrier_4_io_x_hw = dcache_pma_checker__entries_WIRE_8_hw;
    assign dcache_pma_checker_entries_barrier_4_io_x_hx = dcache_pma_checker__entries_WIRE_8_hx;
    assign dcache_pma_checker_entries_barrier_4_io_x_hr = dcache_pma_checker__entries_WIRE_8_hr;
    assign dcache_pma_checker_entries_barrier_4_io_x_pw = dcache_pma_checker__entries_WIRE_8_pw;
    assign dcache_pma_checker_entries_barrier_4_io_x_px = dcache_pma_checker__entries_WIRE_8_px;
    assign dcache_pma_checker_entries_barrier_4_io_x_pr = dcache_pma_checker__entries_WIRE_8_pr;
    assign dcache_pma_checker_entries_barrier_4_io_x_ppp = dcache_pma_checker__entries_WIRE_8_ppp;
    assign dcache_pma_checker_entries_barrier_4_io_x_pal = dcache_pma_checker__entries_WIRE_8_pal;
    assign dcache_pma_checker_entries_barrier_4_io_x_paa = dcache_pma_checker__entries_WIRE_8_paa;
    assign dcache_pma_checker_entries_barrier_4_io_x_eff = dcache_pma_checker__entries_WIRE_8_eff;
    assign dcache_pma_checker_entries_barrier_4_io_x_c = dcache_pma_checker__entries_WIRE_8_c;
    assign dcache_pma_checker_entries_barrier_4_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_8_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_4_io_y_ppn = dcache_pma_checker_entries_barrier_4_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_4_io_y_u = dcache_pma_checker_entries_barrier_4_io_y_u;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_ptw = dcache_pma_checker_entries_barrier_4_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_final = dcache_pma_checker_entries_barrier_4_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_4_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_4_io_y_pf = dcache_pma_checker_entries_barrier_4_io_y_pf;
    assign dcache__pma_checker_entries_barrier_4_io_y_gf = dcache_pma_checker_entries_barrier_4_io_y_gf;
    assign dcache__pma_checker_entries_barrier_4_io_y_sw = dcache_pma_checker_entries_barrier_4_io_y_sw;
    assign dcache__pma_checker_entries_barrier_4_io_y_sx = dcache_pma_checker_entries_barrier_4_io_y_sx;
    assign dcache__pma_checker_entries_barrier_4_io_y_sr = dcache_pma_checker_entries_barrier_4_io_y_sr;
    assign dcache__pma_checker_entries_barrier_4_io_y_hw = dcache_pma_checker_entries_barrier_4_io_y_hw;
    assign dcache__pma_checker_entries_barrier_4_io_y_hx = dcache_pma_checker_entries_barrier_4_io_y_hx;
    assign dcache__pma_checker_entries_barrier_4_io_y_hr = dcache_pma_checker_entries_barrier_4_io_y_hr;
    assign dcache__pma_checker_entries_barrier_4_io_y_pw = dcache_pma_checker_entries_barrier_4_io_y_pw;
    assign dcache__pma_checker_entries_barrier_4_io_y_px = dcache_pma_checker_entries_barrier_4_io_y_px;
    assign dcache__pma_checker_entries_barrier_4_io_y_pr = dcache_pma_checker_entries_barrier_4_io_y_pr;
    assign dcache__pma_checker_entries_barrier_4_io_y_ppp = dcache_pma_checker_entries_barrier_4_io_y_ppp;
    assign dcache__pma_checker_entries_barrier_4_io_y_pal = dcache_pma_checker_entries_barrier_4_io_y_pal;
    assign dcache__pma_checker_entries_barrier_4_io_y_paa = dcache_pma_checker_entries_barrier_4_io_y_paa;
    assign dcache__pma_checker_entries_barrier_4_io_y_eff = dcache_pma_checker_entries_barrier_4_io_y_eff;
    assign dcache__pma_checker_entries_barrier_4_io_y_c = dcache_pma_checker_entries_barrier_4_io_y_c;
    assign dcache_pma_checker_entries_barrier_5_clock = dcache_pma_checker_clock;
    assign dcache_pma_checker_entries_barrier_5_reset = dcache_pma_checker_reset;
    assign dcache_pma_checker_entries_barrier_5_io_x_ppn = dcache_pma_checker__entries_WIRE_10_ppn;
    assign dcache_pma_checker_entries_barrier_5_io_x_u = dcache_pma_checker__entries_WIRE_10_u;
    assign dcache_pma_checker_entries_barrier_5_io_x_g = dcache_pma_checker__entries_WIRE_10_g;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_ptw = dcache_pma_checker__entries_WIRE_10_ae_ptw;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_final = dcache_pma_checker__entries_WIRE_10_ae_final;
    assign dcache_pma_checker_entries_barrier_5_io_x_ae_stage2 = dcache_pma_checker__entries_WIRE_10_ae_stage2;
    assign dcache_pma_checker_entries_barrier_5_io_x_pf = dcache_pma_checker__entries_WIRE_10_pf;
    assign dcache_pma_checker_entries_barrier_5_io_x_gf = dcache_pma_checker__entries_WIRE_10_gf;
    assign dcache_pma_checker_entries_barrier_5_io_x_sw = dcache_pma_checker__entries_WIRE_10_sw;
    assign dcache_pma_checker_entries_barrier_5_io_x_sx = dcache_pma_checker__entries_WIRE_10_sx;
    assign dcache_pma_checker_entries_barrier_5_io_x_sr = dcache_pma_checker__entries_WIRE_10_sr;
    assign dcache_pma_checker_entries_barrier_5_io_x_hw = dcache_pma_checker__entries_WIRE_10_hw;
    assign dcache_pma_checker_entries_barrier_5_io_x_hx = dcache_pma_checker__entries_WIRE_10_hx;
    assign dcache_pma_checker_entries_barrier_5_io_x_hr = dcache_pma_checker__entries_WIRE_10_hr;
    assign dcache_pma_checker_entries_barrier_5_io_x_pw = dcache_pma_checker__entries_WIRE_10_pw;
    assign dcache_pma_checker_entries_barrier_5_io_x_px = dcache_pma_checker__entries_WIRE_10_px;
    assign dcache_pma_checker_entries_barrier_5_io_x_pr = dcache_pma_checker__entries_WIRE_10_pr;
    assign dcache_pma_checker_entries_barrier_5_io_x_ppp = dcache_pma_checker__entries_WIRE_10_ppp;
    assign dcache_pma_checker_entries_barrier_5_io_x_pal = dcache_pma_checker__entries_WIRE_10_pal;
    assign dcache_pma_checker_entries_barrier_5_io_x_paa = dcache_pma_checker__entries_WIRE_10_paa;
    assign dcache_pma_checker_entries_barrier_5_io_x_eff = dcache_pma_checker__entries_WIRE_10_eff;
    assign dcache_pma_checker_entries_barrier_5_io_x_c = dcache_pma_checker__entries_WIRE_10_c;
    assign dcache_pma_checker_entries_barrier_5_io_x_fragmented_superpage = dcache_pma_checker__entries_WIRE_10_fragmented_superpage;
    assign dcache__pma_checker_entries_barrier_5_io_y_ppn = dcache_pma_checker_entries_barrier_5_io_y_ppn;
    assign dcache__pma_checker_entries_barrier_5_io_y_u = dcache_pma_checker_entries_barrier_5_io_y_u;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_ptw = dcache_pma_checker_entries_barrier_5_io_y_ae_ptw;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_final = dcache_pma_checker_entries_barrier_5_io_y_ae_final;
    assign dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 = dcache_pma_checker_entries_barrier_5_io_y_ae_stage2;
    assign dcache__pma_checker_entries_barrier_5_io_y_pf = dcache_pma_checker_entries_barrier_5_io_y_pf;
    assign dcache__pma_checker_entries_barrier_5_io_y_gf = dcache_pma_checker_entries_barrier_5_io_y_gf;
    assign dcache__pma_checker_entries_barrier_5_io_y_sw = dcache_pma_checker_entries_barrier_5_io_y_sw;
    assign dcache__pma_checker_entries_barrier_5_io_y_sx = dcache_pma_checker_entries_barrier_5_io_y_sx;
    assign dcache__pma_checker_entries_barrier_5_io_y_sr = dcache_pma_checker_entries_barrier_5_io_y_sr;
    assign dcache__pma_checker_entries_barrier_5_io_y_hw = dcache_pma_checker_entries_barrier_5_io_y_hw;
    assign dcache__pma_checker_entries_barrier_5_io_y_hx = dcache_pma_checker_entries_barrier_5_io_y_hx;
    assign dcache__pma_checker_entries_barrier_5_io_y_hr = dcache_pma_checker_entries_barrier_5_io_y_hr;
     
    wire[19:0] dcache_pma_checker_ppn =( dcache_pma_checker_hitsVec_0  ?  dcache__pma_checker_entries_barrier_io_y_ppn :20'h0)|( dcache_pma_checker_hitsVec_1  ?  dcache__pma_checker_entries_barrier_1_io_y_ppn :20'h0)|( dcache_pma_checker_hitsVec_2  ?  dcache__pma_checker_entries_barrier_2_io_y_ppn :20'h0)|( dcache_pma_checker_hitsVec_3  ?  dcache__pma_checker_entries_barrier_3_io_y_ppn :20'h0)|( dcache_pma_checker_hitsVec_4  ?  dcache__pma_checker_entries_barrier_4_io_y_ppn :20'h0)|( dcache_pma_checker_hitsVec_5  ?  dcache__pma_checker_entries_barrier_5_io_y_ppn :20'h0)|( dcache_pma_checker_vm_enabled ==1'h0 ?  dcache_pma_checker_vpn [19:0]:20'h0); 
    wire[1:0] dcache_pma_checker_ptw_ae_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_ptw , dcache__pma_checker_entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] dcache_pma_checker_ptw_ae_array_lo ={ dcache_pma_checker_ptw_ae_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_ptw }; 
    wire[1:0] dcache_pma_checker_ptw_ae_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_ptw , dcache__pma_checker_entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] dcache_pma_checker_ptw_ae_array_hi ={ dcache_pma_checker_ptw_ae_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] dcache_pma_checker_ptw_ae_array ={1'h0,{ dcache_pma_checker_ptw_ae_array_hi , dcache_pma_checker_ptw_ae_array_lo }}; 
    wire[1:0] dcache_pma_checker_final_ae_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_final , dcache__pma_checker_entries_barrier_1_io_y_ae_final }; 
    wire[2:0] dcache_pma_checker_final_ae_array_lo ={ dcache_pma_checker_final_ae_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_final }; 
    wire[1:0] dcache_pma_checker_final_ae_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_final , dcache__pma_checker_entries_barrier_4_io_y_ae_final }; 
    wire[2:0] dcache_pma_checker_final_ae_array_hi ={ dcache_pma_checker_final_ae_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_final }; 
    wire[6:0] dcache_pma_checker_final_ae_array ={1'h0,{ dcache_pma_checker_final_ae_array_hi , dcache_pma_checker_final_ae_array_lo }}; 
    wire[1:0] dcache_pma_checker_ptw_pf_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_pf , dcache__pma_checker_entries_barrier_1_io_y_pf }; 
    wire[2:0] dcache_pma_checker_ptw_pf_array_lo ={ dcache_pma_checker_ptw_pf_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_pf }; 
    wire[1:0] dcache_pma_checker_ptw_pf_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_pf , dcache__pma_checker_entries_barrier_4_io_y_pf }; 
    wire[2:0] dcache_pma_checker_ptw_pf_array_hi ={ dcache_pma_checker_ptw_pf_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_pf }; 
    wire[6:0] dcache_pma_checker_ptw_pf_array ={1'h0,{ dcache_pma_checker_ptw_pf_array_hi , dcache_pma_checker_ptw_pf_array_lo }}; 
    wire[1:0] dcache_pma_checker_ptw_gf_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_gf , dcache__pma_checker_entries_barrier_1_io_y_gf }; 
    wire[2:0] dcache_pma_checker_ptw_gf_array_lo ={ dcache_pma_checker_ptw_gf_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_gf }; 
    wire[1:0] dcache_pma_checker_ptw_gf_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_gf , dcache__pma_checker_entries_barrier_4_io_y_gf }; 
    wire[2:0] dcache_pma_checker_ptw_gf_array_hi ={ dcache_pma_checker_ptw_gf_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_gf }; 
    wire[6:0] dcache_pma_checker_ptw_gf_array ={1'h0,{ dcache_pma_checker_ptw_gf_array_hi , dcache_pma_checker_ptw_gf_array_lo }}; 
    wire dcache_pma_checker_sum = dcache_pma_checker_priv_v  ?  dcache_pma_checker_io_ptw_gstatus_sum : dcache_pma_checker_io_ptw_status_sum ; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_u , dcache__pma_checker_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_lo ={ dcache_pma_checker_priv_rw_ok_lo_hi , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_u , dcache__pma_checker_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_hi ={ dcache_pma_checker_priv_rw_ok_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_lo_hi_1 ={ dcache__pma_checker_entries_barrier_2_io_y_u , dcache__pma_checker_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_lo_1 ={ dcache_pma_checker_priv_rw_ok_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_rw_ok_hi_hi_1 ={ dcache__pma_checker_entries_barrier_5_io_y_u , dcache__pma_checker_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_rw_ok_hi_1 ={ dcache_pma_checker_priv_rw_ok_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_pma_checker_priv_rw_ok =( dcache_pma_checker_priv_s ==1'h0| dcache_pma_checker_sum  ? { dcache_pma_checker_priv_rw_ok_hi , dcache_pma_checker_priv_rw_ok_lo }:6'h0)|( dcache_pma_checker_priv_s  ? ~{ dcache_pma_checker_priv_rw_ok_hi_1 , dcache_pma_checker_priv_rw_ok_lo_1 }:6'h0); 
    wire[1:0] dcache_pma_checker_priv_x_ok_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_u , dcache__pma_checker_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_lo ={ dcache_pma_checker_priv_x_ok_lo_hi , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_x_ok_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_u , dcache__pma_checker_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_hi ={ dcache_pma_checker_priv_x_ok_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_x_ok_lo_hi_1 ={ dcache__pma_checker_entries_barrier_2_io_y_u , dcache__pma_checker_entries_barrier_1_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_lo_1 ={ dcache_pma_checker_priv_x_ok_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_u }; 
    wire[1:0] dcache_pma_checker_priv_x_ok_hi_hi_1 ={ dcache__pma_checker_entries_barrier_5_io_y_u , dcache__pma_checker_entries_barrier_4_io_y_u }; 
    wire[2:0] dcache_pma_checker_priv_x_ok_hi_1 ={ dcache_pma_checker_priv_x_ok_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_u }; 
    wire[5:0] dcache_pma_checker_priv_x_ok = dcache_pma_checker_priv_s  ? ~{ dcache_pma_checker_priv_x_ok_hi , dcache_pma_checker_priv_x_ok_lo }:{ dcache_pma_checker_priv_x_ok_hi_1 , dcache_pma_checker_priv_x_ok_lo_1 }; 
    wire[1:0] dcache_pma_checker_stage1_bypass_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_ae_stage2 , dcache__pma_checker_entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] dcache_pma_checker_stage1_bypass_lo ={ dcache_pma_checker_stage1_bypass_lo_hi , dcache__pma_checker_entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] dcache_pma_checker_stage1_bypass_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_ae_stage2 , dcache__pma_checker_entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] dcache_pma_checker_stage1_bypass_hi ={ dcache_pma_checker_stage1_bypass_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_ae_stage2 }; 
    wire dcache_pma_checker_mxr = dcache_pma_checker_io_ptw_status_mxr |( dcache_pma_checker_priv_v  ?  dcache_pma_checker_io_ptw_gstatus_mxr :1'h0); 
    wire[1:0] dcache_pma_checker_r_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_sr , dcache__pma_checker_entries_barrier_1_io_y_sr }; 
    wire[2:0] dcache_pma_checker_r_array_lo ={ dcache_pma_checker_r_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sr }; 
    wire[1:0] dcache_pma_checker_r_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_sr , dcache__pma_checker_entries_barrier_4_io_y_sr }; 
    wire[2:0] dcache_pma_checker_r_array_hi ={ dcache_pma_checker_r_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sr }; 
    wire[1:0] dcache_pma_checker_r_array_lo_hi_1 ={ dcache__pma_checker_entries_barrier_2_io_y_sx , dcache__pma_checker_entries_barrier_1_io_y_sx }; 
    wire[2:0] dcache_pma_checker_r_array_lo_1 ={ dcache_pma_checker_r_array_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_sx }; 
    wire[1:0] dcache_pma_checker_r_array_hi_hi_1 ={ dcache__pma_checker_entries_barrier_5_io_y_sx , dcache__pma_checker_entries_barrier_4_io_y_sx }; 
    wire[2:0] dcache_pma_checker_r_array_hi_1 ={ dcache_pma_checker_r_array_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_pma_checker_r_array ={1'h1, dcache_pma_checker_priv_rw_ok &({ dcache_pma_checker_r_array_hi , dcache_pma_checker_r_array_lo }|( dcache_pma_checker_mxr  ? { dcache_pma_checker_r_array_hi_1 , dcache_pma_checker_r_array_lo_1 }:6'h0))| dcache_pma_checker_stage1_bypass }; 
    wire[1:0] dcache_pma_checker_w_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_sw , dcache__pma_checker_entries_barrier_1_io_y_sw }; 
    wire[2:0] dcache_pma_checker_w_array_lo ={ dcache_pma_checker_w_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sw }; 
    wire[1:0] dcache_pma_checker_w_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_sw , dcache__pma_checker_entries_barrier_4_io_y_sw }; 
    wire[2:0] dcache_pma_checker_w_array_hi ={ dcache_pma_checker_w_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sw }; 
    wire[6:0] dcache_pma_checker_w_array ={1'h1, dcache_pma_checker_priv_rw_ok &{ dcache_pma_checker_w_array_hi , dcache_pma_checker_w_array_lo }| dcache_pma_checker_stage1_bypass }; 
    wire[1:0] dcache_pma_checker_x_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_sx , dcache__pma_checker_entries_barrier_1_io_y_sx }; 
    wire[2:0] dcache_pma_checker_x_array_lo ={ dcache_pma_checker_x_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_sx }; 
    wire[1:0] dcache_pma_checker_x_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_sx , dcache__pma_checker_entries_barrier_4_io_y_sx }; 
    wire[2:0] dcache_pma_checker_x_array_hi ={ dcache_pma_checker_x_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_sx }; 
    wire[6:0] dcache_pma_checker_x_array ={1'h1, dcache_pma_checker_priv_x_ok &{ dcache_pma_checker_x_array_hi , dcache_pma_checker_x_array_lo }| dcache_pma_checker_stage1_bypass }; 
    wire[5:0] dcache_pma_checker_stage2_bypass = dcache_pma_checker_stage2_en ==1'h0 ? 6'h3F:6'h0; 
    wire[1:0] dcache_pma_checker_hr_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_hr , dcache__pma_checker_entries_barrier_1_io_y_hr }; 
    wire[2:0] dcache_pma_checker_hr_array_lo ={ dcache_pma_checker_hr_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hr }; 
    wire[1:0] dcache_pma_checker_hr_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_hr , dcache__pma_checker_entries_barrier_4_io_y_hr }; 
    wire[2:0] dcache_pma_checker_hr_array_hi ={ dcache_pma_checker_hr_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hr }; 
    wire[1:0] dcache_pma_checker_hr_array_lo_hi_1 ={ dcache__pma_checker_entries_barrier_2_io_y_hx , dcache__pma_checker_entries_barrier_1_io_y_hx }; 
    wire[2:0] dcache_pma_checker_hr_array_lo_1 ={ dcache_pma_checker_hr_array_lo_hi_1 , dcache__pma_checker_entries_barrier_io_y_hx }; 
    wire[1:0] dcache_pma_checker_hr_array_hi_hi_1 ={ dcache__pma_checker_entries_barrier_5_io_y_hx , dcache__pma_checker_entries_barrier_4_io_y_hx }; 
    wire[2:0] dcache_pma_checker_hr_array_hi_1 ={ dcache_pma_checker_hr_array_hi_hi_1 , dcache__pma_checker_entries_barrier_3_io_y_hx }; 
    wire[6:0] dcache_pma_checker_hr_array ={1'h1,{ dcache_pma_checker_hr_array_hi , dcache_pma_checker_hr_array_lo }|( dcache_pma_checker_io_ptw_status_mxr  ? { dcache_pma_checker_hr_array_hi_1 , dcache_pma_checker_hr_array_lo_1 }:6'h0)| dcache_pma_checker_stage2_bypass }; 
    wire[1:0] dcache_pma_checker_hw_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_hw , dcache__pma_checker_entries_barrier_1_io_y_hw }; 
    wire[2:0] dcache_pma_checker_hw_array_lo ={ dcache_pma_checker_hw_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hw }; 
    wire[1:0] dcache_pma_checker_hw_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_hw , dcache__pma_checker_entries_barrier_4_io_y_hw }; 
    wire[2:0] dcache_pma_checker_hw_array_hi ={ dcache_pma_checker_hw_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hw }; 
    wire[6:0] dcache_pma_checker_hw_array ={1'h1,{ dcache_pma_checker_hw_array_hi , dcache_pma_checker_hw_array_lo }| dcache_pma_checker_stage2_bypass }; 
    wire[1:0] dcache_pma_checker_hx_array_lo_hi ={ dcache__pma_checker_entries_barrier_2_io_y_hx , dcache__pma_checker_entries_barrier_1_io_y_hx }; 
    wire[2:0] dcache_pma_checker_hx_array_lo ={ dcache_pma_checker_hx_array_lo_hi , dcache__pma_checker_entries_barrier_io_y_hx }; 
    wire[1:0] dcache_pma_checker_hx_array_hi_hi ={ dcache__pma_checker_entries_barrier_5_io_y_hx , dcache__pma_checker_entries_barrier_4_io_y_hx }; 
    wire[2:0] dcache_pma_checker_hx_array_hi ={ dcache_pma_checker_hx_array_hi_hi , dcache__pma_checker_entries_barrier_3_io_y_hx }; 
    wire[6:0] dcache_pma_checker_hx_array ={1'h1,{ dcache_pma_checker_hx_array_hi , dcache_pma_checker_hx_array_lo }| dcache_pma_checker_stage2_bypass }; 
    wire[1:0] dcache_pma_checker_pr_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pr , dcache__pma_checker_entries_barrier_io_y_pr }; 
    wire[1:0] dcache_pma_checker_pr_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pr , dcache__pma_checker_entries_barrier_3_io_y_pr }; 
    wire[2:0] dcache_pma_checker_pr_array_hi ={ dcache_pma_checker_pr_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pr }; 
    wire[6:0] dcache_pma_checker_pr_array ={ dcache_pma_checker_prot_r  ? 2'h3:2'h0,{ dcache_pma_checker_pr_array_hi , dcache_pma_checker_pr_array_lo }}&~( dcache_pma_checker_ptw_ae_array | dcache_pma_checker_final_ae_array ); 
    wire[1:0] dcache_pma_checker_pw_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pw , dcache__pma_checker_entries_barrier_io_y_pw }; 
    wire[1:0] dcache_pma_checker_pw_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pw , dcache__pma_checker_entries_barrier_3_io_y_pw }; 
    wire[2:0] dcache_pma_checker_pw_array_hi ={ dcache_pma_checker_pw_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pw }; 
    wire[6:0] dcache_pma_checker_pw_array ={ dcache_pma_checker_prot_w  ? 2'h3:2'h0,{ dcache_pma_checker_pw_array_hi , dcache_pma_checker_pw_array_lo }}&~( dcache_pma_checker_ptw_ae_array | dcache_pma_checker_final_ae_array ); 
    wire[1:0] dcache_pma_checker_px_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_px , dcache__pma_checker_entries_barrier_io_y_px }; 
    wire[1:0] dcache_pma_checker_px_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_px , dcache__pma_checker_entries_barrier_3_io_y_px }; 
    wire[2:0] dcache_pma_checker_px_array_hi ={ dcache_pma_checker_px_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_px }; 
    wire[6:0] dcache_pma_checker_px_array ={ dcache_pma_checker_prot_x  ? 2'h3:2'h0,{ dcache_pma_checker_px_array_hi , dcache_pma_checker_px_array_lo }}&~( dcache_pma_checker_ptw_ae_array | dcache_pma_checker_final_ae_array ); 
    wire[1:0] dcache_pma_checker_eff_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_eff , dcache__pma_checker_entries_barrier_io_y_eff }; 
    wire[1:0] dcache_pma_checker_eff_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_eff , dcache__pma_checker_entries_barrier_3_io_y_eff }; 
    wire[2:0] dcache_pma_checker_eff_array_hi ={ dcache_pma_checker_eff_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_eff }; 
    wire[6:0] dcache_pma_checker_eff_array ={ dcache_pma_checker_prot_eff  ? 2'h3:2'h0,{ dcache_pma_checker_eff_array_hi , dcache_pma_checker_eff_array_lo }}; 
    wire[1:0] dcache_pma_checker_c_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_c , dcache__pma_checker_entries_barrier_io_y_c }; 
    wire[1:0] dcache_pma_checker_c_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_c , dcache__pma_checker_entries_barrier_3_io_y_c }; 
    wire[2:0] dcache_pma_checker_c_array_hi ={ dcache_pma_checker_c_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_pma_checker_c_array ={ dcache_pma_checker_cacheable  ? 2'h3:2'h0,{ dcache_pma_checker_c_array_hi , dcache_pma_checker_c_array_lo }}; 
    wire[6:0] dcache_pma_checker_lrscAllowed = dcache_pma_checker_c_array ; 
    wire[1:0] dcache_pma_checker_ppp_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_ppp , dcache__pma_checker_entries_barrier_io_y_ppp }; 
    wire[1:0] dcache_pma_checker_ppp_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_ppp , dcache__pma_checker_entries_barrier_3_io_y_ppp }; 
    wire[2:0] dcache_pma_checker_ppp_array_hi ={ dcache_pma_checker_ppp_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_ppp }; 
    wire[6:0] dcache_pma_checker_ppp_array ={ dcache_pma_checker_prot_pp  ? 2'h3:2'h0,{ dcache_pma_checker_ppp_array_hi , dcache_pma_checker_ppp_array_lo }}; 
    wire[1:0] dcache_pma_checker_paa_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_paa , dcache__pma_checker_entries_barrier_io_y_paa }; 
    wire[1:0] dcache_pma_checker_paa_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_paa , dcache__pma_checker_entries_barrier_3_io_y_paa }; 
    wire[2:0] dcache_pma_checker_paa_array_hi ={ dcache_pma_checker_paa_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_paa }; 
    wire[6:0] dcache_pma_checker_paa_array ={ dcache_pma_checker_prot_aa  ? 2'h3:2'h0,{ dcache_pma_checker_paa_array_hi , dcache_pma_checker_paa_array_lo }}; 
    wire[1:0] dcache_pma_checker_pal_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_pal , dcache__pma_checker_entries_barrier_io_y_pal }; 
    wire[1:0] dcache_pma_checker_pal_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_pal , dcache__pma_checker_entries_barrier_3_io_y_pal }; 
    wire[2:0] dcache_pma_checker_pal_array_hi ={ dcache_pma_checker_pal_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_pal }; 
    wire[6:0] dcache_pma_checker_pal_array ={ dcache_pma_checker_prot_al  ? 2'h3:2'h0,{ dcache_pma_checker_pal_array_hi , dcache_pma_checker_pal_array_lo }}; 
    wire[6:0] dcache_pma_checker_ppp_array_if_cached = dcache_pma_checker_ppp_array | dcache_pma_checker_c_array ; 
    wire[6:0] dcache_pma_checker_paa_array_if_cached = dcache_pma_checker_paa_array | dcache_pma_checker_c_array ; 
    wire[6:0] dcache_pma_checker_pal_array_if_cached = dcache_pma_checker_pal_array | dcache_pma_checker_c_array ; 
    wire[1:0] dcache_pma_checker_prefetchable_array_lo ={ dcache__pma_checker_entries_barrier_1_io_y_c , dcache__pma_checker_entries_barrier_io_y_c }; 
    wire[1:0] dcache_pma_checker_prefetchable_array_hi_hi ={ dcache__pma_checker_entries_barrier_4_io_y_c , dcache__pma_checker_entries_barrier_3_io_y_c }; 
    wire[2:0] dcache_pma_checker_prefetchable_array_hi ={ dcache_pma_checker_prefetchable_array_hi_hi , dcache__pma_checker_entries_barrier_2_io_y_c }; 
    wire[6:0] dcache_pma_checker_prefetchable_array ={{ dcache_pma_checker_cacheable & dcache_pma_checker_homogeneous ,1'h0},{ dcache_pma_checker_prefetchable_array_hi , dcache_pma_checker_prefetchable_array_lo }}; 
    wire[4:0] dcache__GEN_74 ={1'h0,4'h1<< dcache_pma_checker_io_req_bits_size }-5'h1; 
    wire dcache_pma_checker_misaligned =|( dcache_pma_checker_io_req_bits_vaddr &{30'h0, dcache__GEN_74 [3:0]}); 
    wire[4:0] dcache_pma_checker_io_req_bits_cmd ; 
    wire dcache_pma_checker_cmd_lrsc =( dcache_pma_checker_io_req_bits_cmd ==5'h6| dcache_pma_checker_io_req_bits_cmd ==5'h7)&1'h1; 
    wire dcache_pma_checker_cmd_amo_logical =( dcache_pma_checker_io_req_bits_cmd ==5'h4| dcache_pma_checker_io_req_bits_cmd ==5'h9| dcache_pma_checker_io_req_bits_cmd ==5'hA| dcache_pma_checker_io_req_bits_cmd ==5'hB)&1'h1; 
    wire dcache_pma_checker_cmd_amo_arithmetic =( dcache_pma_checker_io_req_bits_cmd ==5'h8| dcache_pma_checker_io_req_bits_cmd ==5'hC| dcache_pma_checker_io_req_bits_cmd ==5'hD| dcache_pma_checker_io_req_bits_cmd ==5'hE| dcache_pma_checker_io_req_bits_cmd ==5'hF)&1'h1; 
    wire dcache_pma_checker_cmd_put_partial = dcache_pma_checker_io_req_bits_cmd ==5'h11; 
    wire dcache_pma_checker_cmd_read = dcache_pma_checker_io_req_bits_cmd ==5'h0| dcache_pma_checker_io_req_bits_cmd ==5'h10| dcache_pma_checker_io_req_bits_cmd ==5'h6| dcache_pma_checker_io_req_bits_cmd ==5'h7| dcache_pma_checker_io_req_bits_cmd ==5'h4| dcache_pma_checker_io_req_bits_cmd ==5'h9| dcache_pma_checker_io_req_bits_cmd ==5'hA| dcache_pma_checker_io_req_bits_cmd ==5'hB| dcache_pma_checker_io_req_bits_cmd ==5'h8| dcache_pma_checker_io_req_bits_cmd ==5'hC| dcache_pma_checker_io_req_bits_cmd ==5'hD| dcache_pma_checker_io_req_bits_cmd ==5'hE| dcache_pma_checker_io_req_bits_cmd ==5'hF; 
    wire dcache_pma_checker_cmd_write = dcache_pma_checker_io_req_bits_cmd ==5'h1| dcache_pma_checker_io_req_bits_cmd ==5'h11| dcache_pma_checker_io_req_bits_cmd ==5'h7| dcache_pma_checker_io_req_bits_cmd ==5'h4| dcache_pma_checker_io_req_bits_cmd ==5'h9| dcache_pma_checker_io_req_bits_cmd ==5'hA| dcache_pma_checker_io_req_bits_cmd ==5'hB| dcache_pma_checker_io_req_bits_cmd ==5'h8| dcache_pma_checker_io_req_bits_cmd ==5'hC| dcache_pma_checker_io_req_bits_cmd ==5'hD| dcache_pma_checker_io_req_bits_cmd ==5'hE| dcache_pma_checker_io_req_bits_cmd ==5'hF; 
    wire dcache_pma_checker_cmd_write_perms = dcache_pma_checker_cmd_write | dcache_pma_checker_io_req_bits_cmd ==5'h5| dcache_pma_checker_io_req_bits_cmd ==5'h17; 
    wire[6:0] dcache_pma_checker_ae_array =( dcache_pma_checker_misaligned  ?  dcache_pma_checker_eff_array :7'h0)|( dcache_pma_checker_cmd_lrsc  ? ~ dcache_pma_checker_lrscAllowed :7'h0); 
    wire[6:0] dcache_pma_checker_ae_ld_array = dcache_pma_checker_cmd_read  ?  dcache_pma_checker_ae_array |~ dcache_pma_checker_pr_array :7'h0; 
    wire[6:0] dcache_pma_checker_ae_st_array =( dcache_pma_checker_cmd_write_perms  ?  dcache_pma_checker_ae_array |~ dcache_pma_checker_pw_array :7'h0)|( dcache_pma_checker_cmd_put_partial  ? ~ dcache_pma_checker_ppp_array_if_cached :7'h0)|( dcache_pma_checker_cmd_amo_logical  ? ~ dcache_pma_checker_pal_array_if_cached :7'h0)|( dcache_pma_checker_cmd_amo_arithmetic  ? ~ dcache_pma_checker_paa_array_if_cached :7'h0); 
    wire[6:0] dcache_pma_checker_must_alloc_array =( dcache_pma_checker_cmd_put_partial  ? ~ dcache_pma_checker_ppp_array :7'h0)|( dcache_pma_checker_cmd_amo_logical  ? ~ dcache_pma_checker_pal_array :7'h0)|( dcache_pma_checker_cmd_amo_arithmetic  ? ~ dcache_pma_checker_paa_array :7'h0)|( dcache_pma_checker_cmd_lrsc  ? 7'h7F:7'h0); 
    wire[6:0] dcache_pma_checker_pf_ld_array = dcache_pma_checker_cmd_read  ? (~( dcache_pma_checker_cmd_readx  ?  dcache_pma_checker_x_array : dcache_pma_checker_r_array )&~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array :7'h0; 
    wire[6:0] dcache_pma_checker_pf_st_array = dcache_pma_checker_cmd_write_perms  ? (~ dcache_pma_checker_w_array &~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array :7'h0; 
    wire[6:0] dcache_pma_checker_pf_inst_array =(~ dcache_pma_checker_x_array &~ dcache_pma_checker_ptw_ae_array | dcache_pma_checker_ptw_pf_array )&~ dcache_pma_checker_ptw_gf_array ; 
    wire[6:0] dcache_pma_checker_gf_ld_array = dcache_pma_checker_priv_v & dcache_pma_checker_cmd_read  ? (~( dcache_pma_checker_cmd_readx  ?  dcache_pma_checker_hx_array : dcache_pma_checker_hr_array )| dcache_pma_checker_ptw_gf_array )&~ dcache_pma_checker_ptw_ae_array :7'h0; 
    wire[6:0] dcache_pma_checker_gf_st_array = dcache_pma_checker_priv_v & dcache_pma_checker_cmd_write_perms  ? (~ dcache_pma_checker_hw_array | dcache_pma_checker_ptw_gf_array )&~ dcache_pma_checker_ptw_ae_array :7'h0; 
    wire[6:0] dcache_pma_checker_gf_inst_array = dcache_pma_checker_priv_v  ? (~ dcache_pma_checker_hx_array | dcache_pma_checker_ptw_gf_array )&~ dcache_pma_checker_ptw_ae_array :7'h0; 
    wire[6:0] dcache_pma_checker_gpa_hits_need_gpa_mask = dcache_pma_checker_gf_ld_array | dcache_pma_checker_gf_st_array ; 
    wire[5:0] dcache_pma_checker_gpa_hits_hit_mask ={1'h0, dcache_pma_checker_r_gpa_valid & dcache_pma_checker_r_gpa_vpn == dcache_pma_checker_vpn  ? 5'h1F:5'h0}|( dcache_pma_checker_vstage1_en ==1'h0 ? 6'h3F:6'h0); 
    wire[5:0] dcache_pma_checker_gpa_hits = dcache_pma_checker_gpa_hits_hit_mask |~( dcache_pma_checker_gpa_hits_need_gpa_mask [5:0]); 
    wire dcache_pma_checker_tlb_hit_if_not_gpa_miss =| dcache_pma_checker_real_hits ; 
    wire dcache_pma_checker_tlb_hit =|( dcache_pma_checker_real_hits & dcache_pma_checker_gpa_hits ); 
    wire dcache_pma_checker_tlb_miss = dcache_pma_checker_vm_enabled & dcache_pma_checker_vsatp_mode_mismatch ==1'h0& dcache_pma_checker_tlb_hit ==1'h0; reg[2:0] dcache_pma_checker_state_reg_1 ; 
    wire dcache__GEN_75 = dcache_pma_checker_io_req_valid & dcache_pma_checker_vm_enabled ; 
    wire dcache__GEN_76 = dcache_pma_checker_superpage_hits_0 | dcache_pma_checker_superpage_hits_1 | dcache_pma_checker_superpage_hits_2 | dcache_pma_checker_superpage_hits_3 ; 
    wire[1:0] dcache_pma_checker_lo ={ dcache_pma_checker_superpage_hits_1 , dcache_pma_checker_superpage_hits_0 }; 
    wire[1:0] dcache_pma_checker_hi ={ dcache_pma_checker_superpage_hits_3 , dcache_pma_checker_superpage_hits_2 }; 
    wire[3:0] dcache__GEN_77 ={ dcache_pma_checker_hi , dcache_pma_checker_lo }; 
    wire[1:0] dcache_pma_checker_hi_1 = dcache__GEN_77 [3:2]; 
    wire[1:0] dcache_pma_checker_lo_1 = dcache__GEN_77 [1:0]; 
    wire[1:0] dcache__GEN_78 = dcache_pma_checker_hi_1 | dcache_pma_checker_lo_1 ; 
    wire[1:0] dcache_pma_checker_state_reg_touch_way_sized ={| dcache_pma_checker_hi_1 , dcache__GEN_78 [1]}; 
    wire dcache_pma_checker_state_reg_set_left_older = dcache_pma_checker_state_reg_touch_way_sized [1]==1'h0; 
    wire dcache_pma_checker_state_reg_left_subtree_state = dcache_pma_checker_state_reg_1 [1]; 
    wire dcache_pma_checker_state_reg_right_subtree_state = dcache_pma_checker_state_reg_1 [0]; 
    wire[1:0] dcache_pma_checker_state_reg_hi ={ dcache_pma_checker_state_reg_set_left_older , dcache_pma_checker_state_reg_set_left_older  ?  dcache_pma_checker_state_reg_left_subtree_state : dcache_pma_checker_state_reg_touch_way_sized [0]==1'h0}; 
    wire[2:0] dcache__GEN_79 ={ dcache_pma_checker_state_reg_hi , dcache_pma_checker_state_reg_set_left_older  ?  dcache_pma_checker_state_reg_touch_way_sized [0]==1'h0: dcache_pma_checker_state_reg_right_subtree_state }; 
    wire[2:0] dcache__pma_checker_real_hits_2to0 = dcache_pma_checker_real_hits [2:0]; 
    wire dcache_pma_checker_multipleHits_leftOne = dcache__pma_checker_real_hits_2to0 [0]; 
    wire[1:0] dcache__pma_checker_real_hits_2to0_2to1 = dcache__pma_checker_real_hits_2to0 [2:1]; 
    wire dcache_pma_checker_multipleHits_leftOne_1 = dcache__pma_checker_real_hits_2to0_2to1 [0]; 
    wire dcache_pma_checker_multipleHits_rightOne = dcache__pma_checker_real_hits_2to0_2to1 [1]; 
    wire dcache_pma_checker_multipleHits_rightOne_1 = dcache_pma_checker_multipleHits_leftOne_1 | dcache_pma_checker_multipleHits_rightOne ; 
    wire dcache_pma_checker_multipleHits_rightTwo = dcache_pma_checker_multipleHits_leftOne_1 & dcache_pma_checker_multipleHits_rightOne |1'h0; 
    wire dcache_pma_checker_multipleHits_leftOne_2 = dcache_pma_checker_multipleHits_leftOne | dcache_pma_checker_multipleHits_rightOne_1 ; 
    wire dcache_pma_checker_multipleHits_leftTwo = dcache_pma_checker_multipleHits_rightTwo |1'h0| dcache_pma_checker_multipleHits_leftOne & dcache_pma_checker_multipleHits_rightOne_1 ; 
    wire[2:0] dcache__pma_checker_real_hits_5to3 = dcache_pma_checker_real_hits [5:3]; 
    wire dcache_pma_checker_multipleHits_leftOne_3 = dcache__pma_checker_real_hits_5to3 [0]; 
    wire[1:0] dcache__pma_checker_real_hits_5to3_2to1 = dcache__pma_checker_real_hits_5to3 [2:1]; 
    wire dcache_pma_checker_multipleHits_leftOne_4 = dcache__pma_checker_real_hits_5to3_2to1 [0]; 
    wire dcache_pma_checker_multipleHits_rightOne_2 = dcache__pma_checker_real_hits_5to3_2to1 [1]; 
    wire dcache_pma_checker_multipleHits_rightOne_3 = dcache_pma_checker_multipleHits_leftOne_4 | dcache_pma_checker_multipleHits_rightOne_2 ; 
    wire dcache_pma_checker_multipleHits_rightTwo_1 = dcache_pma_checker_multipleHits_leftOne_4 & dcache_pma_checker_multipleHits_rightOne_2 |1'h0; 
    wire dcache_pma_checker_multipleHits_rightOne_4 = dcache_pma_checker_multipleHits_leftOne_3 | dcache_pma_checker_multipleHits_rightOne_3 ; 
    wire dcache_pma_checker_multipleHits_rightTwo_2 = dcache_pma_checker_multipleHits_rightTwo_1 |1'h0| dcache_pma_checker_multipleHits_leftOne_3 & dcache_pma_checker_multipleHits_rightOne_3 ; 
    wire dcache_pma_checker_multipleHits = dcache_pma_checker_multipleHits_leftTwo | dcache_pma_checker_multipleHits_rightTwo_2 | dcache_pma_checker_multipleHits_leftOne_2 & dcache_pma_checker_multipleHits_rightOne_4 ; 
    wire dcache_pma_checker_io_req_ready = dcache_pma_checker_state ==2'h0; 
    wire dcache_pma_checker_io_resp_pf_ld =(|( dcache_pma_checker_pf_ld_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_pf_st =(|( dcache_pma_checker_pf_st_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_pf_inst =(|( dcache_pma_checker_pf_inst_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_gf_ld =(|( dcache_pma_checker_gf_ld_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_gf_st =(|( dcache_pma_checker_gf_st_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_gf_inst =(|( dcache_pma_checker_gf_inst_array & dcache_pma_checker_hits ))|1'h0; 
    wire dcache_pma_checker_io_resp_ae_ld =|( dcache_pma_checker_ae_ld_array & dcache_pma_checker_hits ); 
    wire dcache_pma_checker_io_resp_ae_st =|( dcache_pma_checker_ae_st_array & dcache_pma_checker_hits ); 
    wire dcache_pma_checker_io_resp_ae_inst =|(~ dcache_pma_checker_px_array & dcache_pma_checker_hits ); 
    wire dcache_pma_checker_io_resp_ma_ld = dcache_pma_checker_misaligned & dcache_pma_checker_cmd_read ; 
    wire dcache_pma_checker_io_resp_ma_st = dcache_pma_checker_misaligned & dcache_pma_checker_cmd_write ; 
    wire dcache_pma_checker_io_resp_cacheable =|( dcache_pma_checker_c_array & dcache_pma_checker_hits ); 
    wire dcache_pma_checker_io_resp_must_alloc =|( dcache_pma_checker_must_alloc_array & dcache_pma_checker_hits ); 
    wire dcache_pma_checker_io_resp_miss = dcache_pma_checker_do_refill | dcache_pma_checker_vsatp_mode_mismatch | dcache_pma_checker_tlb_miss | dcache_pma_checker_multipleHits ; 
    wire[31:0] dcache_pma_checker_io_resp_paddr ={ dcache_pma_checker_ppn , dcache_pma_checker_io_req_bits_vaddr [11:0]}; 
    wire dcache_pma_checker_io_resp_gpa_is_pte = dcache_pma_checker_vstage1_en & dcache_pma_checker_r_gpa_is_pte ; 
    wire[21:0] dcache_pma_checker_io_resp_gpa_page = dcache_pma_checker_vstage1_en ==1'h0 ? {1'h0, dcache_pma_checker_vpn }:{1'h0, dcache_pma_checker_r_gpa [32:12]}; 
    wire[11:0] dcache_pma_checker_io_resp_gpa_offset = dcache_pma_checker_io_resp_gpa_is_pte  ?  dcache_pma_checker_r_gpa [11:0]: dcache_pma_checker_io_req_bits_vaddr [11:0]; 
    wire[33:0] dcache_pma_checker_io_resp_gpa ={ dcache_pma_checker_io_resp_gpa_page , dcache_pma_checker_io_resp_gpa_offset }; 
    wire dcache_pma_checker_io_ptw_req_valid = dcache_pma_checker_state ==2'h1; 
    wire dcache_pma_checker_io_ptw_req_bits_valid = dcache_pma_checker_io_kill ==1'h0; 
    wire dcache_replace ;  
    wire dcache_lfsr_prng_clock;
    wire dcache_lfsr_prng_reset;
    wire dcache_lfsr_prng_io_seed_valid;
    wire dcache_lfsr_prng_io_seed_bits_0;
    wire dcache_lfsr_prng_io_seed_bits_1;
    wire dcache_lfsr_prng_io_seed_bits_2;
    wire dcache_lfsr_prng_io_seed_bits_3;
    wire dcache_lfsr_prng_io_seed_bits_4;
    wire dcache_lfsr_prng_io_seed_bits_5;
    wire dcache_lfsr_prng_io_seed_bits_6;
    wire dcache_lfsr_prng_io_seed_bits_7;
    wire dcache_lfsr_prng_io_seed_bits_8;
    wire dcache_lfsr_prng_io_seed_bits_9;
    wire dcache_lfsr_prng_io_seed_bits_10;
    wire dcache_lfsr_prng_io_seed_bits_11;
    wire dcache_lfsr_prng_io_seed_bits_12;
    wire dcache_lfsr_prng_io_seed_bits_13;
    wire dcache_lfsr_prng_io_seed_bits_14;
    wire dcache_lfsr_prng_io_seed_bits_15;
    wire dcache_lfsr_prng_io_increment;
    wire dcache_lfsr_prng_io_out_0;
    wire dcache_lfsr_prng_io_out_1;
    wire dcache_lfsr_prng_io_out_2;
    wire dcache_lfsr_prng_io_out_3;
    wire dcache_lfsr_prng_io_out_4;
    wire dcache_lfsr_prng_io_out_5;
    wire dcache_lfsr_prng_io_out_6;
    wire dcache_lfsr_prng_io_out_7;
    wire dcache_lfsr_prng_io_out_8;
    wire dcache_lfsr_prng_io_out_9;
    wire dcache_lfsr_prng_io_out_10;
    wire dcache_lfsr_prng_io_out_11;
    wire dcache_lfsr_prng_io_out_12;
    wire dcache_lfsr_prng_io_out_13;
    wire dcache_lfsr_prng_io_out_14;
    wire dcache_lfsr_prng_io_out_15;

    wire dcache_lfsr_prng__state_WIRE_1 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_2 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_3 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_4 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_5 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_6 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_7 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_8 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_9 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_10 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_11 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_12 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_13 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_14 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_15 =1'h0; 
    wire dcache_lfsr_prng__state_WIRE_0 =1'h1; 
    reg dcache_lfsr_prng_state_0 ; 
    reg dcache_lfsr_prng_state_1 ; 
    reg dcache_lfsr_prng_state_2 ; 
    reg dcache_lfsr_prng_state_3 ; 
    reg dcache_lfsr_prng_state_4 ; 
    reg dcache_lfsr_prng_state_5 ; 
    reg dcache_lfsr_prng_state_6 ; 
    reg dcache_lfsr_prng_state_7 ; 
    reg dcache_lfsr_prng_state_8 ; 
    reg dcache_lfsr_prng_state_9 ; 
    reg dcache_lfsr_prng_state_10 ; 
    reg dcache_lfsr_prng_state_11 ; 
    reg dcache_lfsr_prng_state_12 ; 
    reg dcache_lfsr_prng_state_13 ; 
    reg dcache_lfsr_prng_state_14 ; 
    reg dcache_lfsr_prng_state_15 ; 
    wire dcache_lfsr_prng__GEN = dcache_lfsr_prng_state_15 ^ dcache_lfsr_prng_state_13 ^ dcache_lfsr_prng_state_12 ^ dcache_lfsr_prng_state_10 ; 
  always @( posedge  dcache_lfsr_prng_clock )
         begin 
             if ( dcache_lfsr_prng_reset )
                 begin  
                     dcache_lfsr_prng_state_0  <= dcache_lfsr_prng__state_WIRE_0 ; 
                     dcache_lfsr_prng_state_1  <= dcache_lfsr_prng__state_WIRE_1 ; 
                     dcache_lfsr_prng_state_2  <= dcache_lfsr_prng__state_WIRE_2 ; 
                     dcache_lfsr_prng_state_3  <= dcache_lfsr_prng__state_WIRE_3 ; 
                     dcache_lfsr_prng_state_4  <= dcache_lfsr_prng__state_WIRE_4 ; 
                     dcache_lfsr_prng_state_5  <= dcache_lfsr_prng__state_WIRE_5 ; 
                     dcache_lfsr_prng_state_6  <= dcache_lfsr_prng__state_WIRE_6 ; 
                     dcache_lfsr_prng_state_7  <= dcache_lfsr_prng__state_WIRE_7 ; 
                     dcache_lfsr_prng_state_8  <= dcache_lfsr_prng__state_WIRE_8 ; 
                     dcache_lfsr_prng_state_9  <= dcache_lfsr_prng__state_WIRE_9 ; 
                     dcache_lfsr_prng_state_10  <= dcache_lfsr_prng__state_WIRE_10 ; 
                     dcache_lfsr_prng_state_11  <= dcache_lfsr_prng__state_WIRE_11 ; 
                     dcache_lfsr_prng_state_12  <= dcache_lfsr_prng__state_WIRE_12 ; 
                     dcache_lfsr_prng_state_13  <= dcache_lfsr_prng__state_WIRE_13 ; 
                     dcache_lfsr_prng_state_14  <= dcache_lfsr_prng__state_WIRE_14 ; 
                     dcache_lfsr_prng_state_15  <= dcache_lfsr_prng__state_WIRE_15 ;
                 end 
              else 
                 if ( dcache_lfsr_prng_io_seed_valid )
                     begin  
                         dcache_lfsr_prng_state_0  <= dcache_lfsr_prng_io_seed_bits_0 ; 
                         dcache_lfsr_prng_state_1  <= dcache_lfsr_prng_io_seed_bits_1 ; 
                         dcache_lfsr_prng_state_2  <= dcache_lfsr_prng_io_seed_bits_2 ; 
                         dcache_lfsr_prng_state_3  <= dcache_lfsr_prng_io_seed_bits_3 ; 
                         dcache_lfsr_prng_state_4  <= dcache_lfsr_prng_io_seed_bits_4 ; 
                         dcache_lfsr_prng_state_5  <= dcache_lfsr_prng_io_seed_bits_5 ; 
                         dcache_lfsr_prng_state_6  <= dcache_lfsr_prng_io_seed_bits_6 ; 
                         dcache_lfsr_prng_state_7  <= dcache_lfsr_prng_io_seed_bits_7 ; 
                         dcache_lfsr_prng_state_8  <= dcache_lfsr_prng_io_seed_bits_8 ; 
                         dcache_lfsr_prng_state_9  <= dcache_lfsr_prng_io_seed_bits_9 ; 
                         dcache_lfsr_prng_state_10  <= dcache_lfsr_prng_io_seed_bits_10 ; 
                         dcache_lfsr_prng_state_11  <= dcache_lfsr_prng_io_seed_bits_11 ; 
                         dcache_lfsr_prng_state_12  <= dcache_lfsr_prng_io_seed_bits_12 ; 
                         dcache_lfsr_prng_state_13  <= dcache_lfsr_prng_io_seed_bits_13 ; 
                         dcache_lfsr_prng_state_14  <= dcache_lfsr_prng_io_seed_bits_14 ; 
                         dcache_lfsr_prng_state_15  <= dcache_lfsr_prng_io_seed_bits_15 ;
                     end 
                  else 
                     if ( dcache_lfsr_prng_io_increment )
                         begin  
                             dcache_lfsr_prng_state_0  <= dcache_lfsr_prng__GEN ; 
                             dcache_lfsr_prng_state_1  <= dcache_lfsr_prng_state_0 ; 
                             dcache_lfsr_prng_state_2  <= dcache_lfsr_prng_state_1 ; 
                             dcache_lfsr_prng_state_3  <= dcache_lfsr_prng_state_2 ; 
                             dcache_lfsr_prng_state_4  <= dcache_lfsr_prng_state_3 ; 
                             dcache_lfsr_prng_state_5  <= dcache_lfsr_prng_state_4 ; 
                             dcache_lfsr_prng_state_6  <= dcache_lfsr_prng_state_5 ; 
                             dcache_lfsr_prng_state_7  <= dcache_lfsr_prng_state_6 ; 
                             dcache_lfsr_prng_state_8  <= dcache_lfsr_prng_state_7 ; 
                             dcache_lfsr_prng_state_9  <= dcache_lfsr_prng_state_8 ; 
                             dcache_lfsr_prng_state_10  <= dcache_lfsr_prng_state_9 ; 
                             dcache_lfsr_prng_state_11  <= dcache_lfsr_prng_state_10 ; 
                             dcache_lfsr_prng_state_12  <= dcache_lfsr_prng_state_11 ; 
                             dcache_lfsr_prng_state_13  <= dcache_lfsr_prng_state_12 ; 
                             dcache_lfsr_prng_state_14  <= dcache_lfsr_prng_state_13 ; 
                             dcache_lfsr_prng_state_15  <= dcache_lfsr_prng_state_14 ;
                         end 
                      else 
                         begin 
                         end 
         end
  assign  dcache_lfsr_prng_io_out_0 = dcache_lfsr_prng_state_0 ; 
  assign  dcache_lfsr_prng_io_out_1 = dcache_lfsr_prng_state_1 ; 
  assign  dcache_lfsr_prng_io_out_2 = dcache_lfsr_prng_state_2 ; 
  assign  dcache_lfsr_prng_io_out_3 = dcache_lfsr_prng_state_3 ; 
  assign  dcache_lfsr_prng_io_out_4 = dcache_lfsr_prng_state_4 ; 
  assign  dcache_lfsr_prng_io_out_5 = dcache_lfsr_prng_state_5 ; 
  assign  dcache_lfsr_prng_io_out_6 = dcache_lfsr_prng_state_6 ; 
  assign  dcache_lfsr_prng_io_out_7 = dcache_lfsr_prng_state_7 ; 
  assign  dcache_lfsr_prng_io_out_8 = dcache_lfsr_prng_state_8 ; 
  assign  dcache_lfsr_prng_io_out_9 = dcache_lfsr_prng_state_9 ; 
  assign  dcache_lfsr_prng_io_out_10 = dcache_lfsr_prng_state_10 ; 
  assign  dcache_lfsr_prng_io_out_11 = dcache_lfsr_prng_state_11 ; 
  assign  dcache_lfsr_prng_io_out_12 = dcache_lfsr_prng_state_12 ; 
  assign  dcache_lfsr_prng_io_out_13 = dcache_lfsr_prng_state_13 ; 
  assign  dcache_lfsr_prng_io_out_14 = dcache_lfsr_prng_state_14 ; 
  assign  dcache_lfsr_prng_io_out_15 = dcache_lfsr_prng_state_15 ;
    assign dcache_lfsr_prng_clock = dcache_clock;
    assign dcache_lfsr_prng_reset = dcache_reset;
    assign dcache_lfsr_prng_io_seed_valid = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_0 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_1 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_2 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_3 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_4 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_5 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_6 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_7 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_8 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_9 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_10 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_11 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_12 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_13 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_14 = 1'h0;
    assign dcache_lfsr_prng_io_seed_bits_15 = 1'h0;
    assign dcache_lfsr_prng_io_increment = dcache_replace;
    assign dcache__lfsr_prng_io_out_0 = dcache_lfsr_prng_io_out_0;
    assign dcache__lfsr_prng_io_out_1 = dcache_lfsr_prng_io_out_1;
    assign dcache__lfsr_prng_io_out_2 = dcache_lfsr_prng_io_out_2;
    assign dcache__lfsr_prng_io_out_3 = dcache_lfsr_prng_io_out_3;
    assign dcache__lfsr_prng_io_out_4 = dcache_lfsr_prng_io_out_4;
    assign dcache__lfsr_prng_io_out_5 = dcache_lfsr_prng_io_out_5;
    assign dcache__lfsr_prng_io_out_6 = dcache_lfsr_prng_io_out_6;
    assign dcache__lfsr_prng_io_out_7 = dcache_lfsr_prng_io_out_7;
    assign dcache__lfsr_prng_io_out_8 = dcache_lfsr_prng_io_out_8;
    assign dcache__lfsr_prng_io_out_9 = dcache_lfsr_prng_io_out_9;
    assign dcache__lfsr_prng_io_out_10 = dcache_lfsr_prng_io_out_10;
    assign dcache__lfsr_prng_io_out_11 = dcache_lfsr_prng_io_out_11;
    assign dcache__lfsr_prng_io_out_12 = dcache_lfsr_prng_io_out_12;
    assign dcache__lfsr_prng_io_out_13 = dcache_lfsr_prng_io_out_13;
    assign dcache__lfsr_prng_io_out_14 = dcache_lfsr_prng_io_out_14;
    assign dcache__lfsr_prng_io_out_15 = dcache_lfsr_prng_io_out_15;
     
    wire[1:0] dcache_lfsr_lo_lo_lo ={ dcache__lfsr_prng_io_out_1 , dcache__lfsr_prng_io_out_0 }; 
    wire[1:0] dcache_lfsr_lo_lo_hi ={ dcache__lfsr_prng_io_out_3 , dcache__lfsr_prng_io_out_2 }; 
    wire[3:0] dcache_lfsr_lo_lo ={ dcache_lfsr_lo_lo_hi , dcache_lfsr_lo_lo_lo }; 
    wire[1:0] dcache_lfsr_lo_hi_lo ={ dcache__lfsr_prng_io_out_5 , dcache__lfsr_prng_io_out_4 }; 
    wire[1:0] dcache_lfsr_lo_hi_hi ={ dcache__lfsr_prng_io_out_7 , dcache__lfsr_prng_io_out_6 }; 
    wire[3:0] dcache_lfsr_lo_hi ={ dcache_lfsr_lo_hi_hi , dcache_lfsr_lo_hi_lo }; 
    wire[7:0] dcache_lfsr_lo ={ dcache_lfsr_lo_hi , dcache_lfsr_lo_lo }; 
    wire[1:0] dcache_lfsr_hi_lo_lo ={ dcache__lfsr_prng_io_out_9 , dcache__lfsr_prng_io_out_8 }; 
    wire[1:0] dcache_lfsr_hi_lo_hi ={ dcache__lfsr_prng_io_out_11 , dcache__lfsr_prng_io_out_10 }; 
    wire[3:0] dcache_lfsr_hi_lo ={ dcache_lfsr_hi_lo_hi , dcache_lfsr_hi_lo_lo }; 
    wire[1:0] dcache_lfsr_hi_hi_lo ={ dcache__lfsr_prng_io_out_13 , dcache__lfsr_prng_io_out_12 }; 
    wire[1:0] dcache_lfsr_hi_hi_hi ={ dcache__lfsr_prng_io_out_15 , dcache__lfsr_prng_io_out_14 }; 
    wire[3:0] dcache_lfsr_hi_hi ={ dcache_lfsr_hi_hi_hi , dcache_lfsr_hi_hi_lo }; 
    wire[7:0] dcache_lfsr_hi ={ dcache_lfsr_hi_hi , dcache_lfsr_hi_lo }; 
    wire[15:0] dcache_lfsr ={ dcache_lfsr_hi , dcache_lfsr_lo }; 
    wire[33:0] dcache_metaArb_io_in_5_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_5_bits_idx ; 
    wire dcache_metaArb_io_in_5_bits_way_en = dcache_metaArb_io_in_4_bits_way_en ; 
    wire dcache_metaArb_io_in_6_bits_way_en = dcache_metaArb_io_in_4_bits_way_en ; 
    wire dcache_metaArb_io_in_7_bits_way_en = dcache_metaArb_io_in_4_bits_way_en ; 
    wire[21:0] dcache_metaArb_io_in_5_bits_data = dcache_metaArb_io_in_4_bits_data ; 
    wire[21:0] dcache_metaArb_io_in_6_bits_data = dcache_metaArb_io_in_4_bits_data ; 
    wire[21:0] dcache_metaArb_io_in_7_bits_data = dcache_metaArb_io_in_4_bits_data ; 
    wire[33:0] dcache_metaArb_io_in_0_bits_addr = dcache_metaArb_io_in_5_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_0_bits_idx = dcache_metaArb_io_in_5_bits_idx ; 
    wire[5:0] dcache_tag_array_MPORT_addr = dcache_metaArb_io_out_bits_idx ; 
    wire[5:0] dcache__s1_meta_WIRE = dcache_metaArb_io_out_bits_idx ; 
    wire[21:0] dcache__GEN_80 = dcache_metaArb_io_out_bits_data ; 
    wire dcache_metaArb_io_in_6_valid ; 
    wire[33:0] dcache_metaArb_io_in_6_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_6_bits_idx ; 
    wire[5:0] dcache_metaArb_io_in_7_bits_idx ; 
    wire dcache_metaArb_io_in_5_valid ; 
    wire dcache_metaArb_io_in_4_valid ; 
    wire[33:0] dcache_metaArb_io_in_4_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_4_bits_idx ; 
    wire dcache_metaArb_io_in_3_valid ; 
    wire[33:0] dcache_metaArb_io_in_3_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_3_bits_idx ; 
    wire dcache_metaArb_io_in_3_bits_way_en ; 
    wire[21:0] dcache_metaArb_io_in_3_bits_data ; 
    wire dcache_metaArb_io_in_2_valid ; 
    wire dcache_metaArb_io_in_2_bits_write ; 
    wire[33:0] dcache_metaArb_io_in_2_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_2_bits_idx ; 
    wire dcache_metaArb_io_in_2_bits_way_en ; 
    wire[21:0] dcache_metaArb_io_in_2_bits_data ; 
    wire dcache_metaArb_io_in_1_valid ; 
    wire[33:0] dcache_metaArb_io_in_1_bits_addr ; 
    wire[5:0] dcache_metaArb_io_in_1_bits_idx ; 
    wire dcache_metaArb_io_in_1_bits_way_en ; 
    wire[21:0] dcache_metaArb_io_in_1_bits_data ; 
    wire dcache_metaArb_io_in_0_valid ; 
    wire[2:0] dcache_metaArb_io_chosen = dcache_metaArb_io_in_0_valid  ? 3'h0: dcache_metaArb_io_in_1_valid  ? 3'h1: dcache_metaArb_io_in_2_valid  ? 3'h2: dcache_metaArb_io_in_3_valid  ? 3'h3: dcache_metaArb_io_in_4_valid  ? 3'h4: dcache_metaArb_io_in_5_valid  ? 3'h5: dcache_metaArb_io_in_6_valid  ? 3'h6:3'h7; 
    wire dcache_metaArb_io_out_bits_write = dcache_metaArb_io_in_0_valid  ?  dcache_metaArb_io_in_0_bits_write : dcache_metaArb_io_in_1_valid  ?  dcache_metaArb_io_in_1_bits_write : dcache_metaArb_io_in_2_valid  ?  dcache_metaArb_io_in_2_bits_write : dcache_metaArb_io_in_3_valid  ?  dcache_metaArb_io_in_3_bits_write : dcache_metaArb_io_in_4_valid  ?  dcache_metaArb_io_in_4_bits_write : dcache_metaArb_io_in_5_valid  ?  dcache_metaArb_io_in_5_bits_write : dcache_metaArb_io_in_6_valid  ?  dcache_metaArb_io_in_6_bits_write : dcache_metaArb_io_in_7_bits_write ; 
    wire[33:0] dcache_metaArb_io_out_bits_addr = dcache_metaArb_io_in_0_valid  ?  dcache_metaArb_io_in_0_bits_addr : dcache_metaArb_io_in_1_valid  ?  dcache_metaArb_io_in_1_bits_addr : dcache_metaArb_io_in_2_valid  ?  dcache_metaArb_io_in_2_bits_addr : dcache_metaArb_io_in_3_valid  ?  dcache_metaArb_io_in_3_bits_addr : dcache_metaArb_io_in_4_valid  ?  dcache_metaArb_io_in_4_bits_addr : dcache_metaArb_io_in_5_valid  ?  dcache_metaArb_io_in_5_bits_addr : dcache_metaArb_io_in_6_valid  ?  dcache_metaArb_io_in_6_bits_addr : dcache_metaArb_io_in_7_bits_addr ; 
  assign  dcache_metaArb_io_out_bits_idx = dcache_metaArb_io_in_0_valid  ?  dcache_metaArb_io_in_0_bits_idx : dcache_metaArb_io_in_1_valid  ?  dcache_metaArb_io_in_1_bits_idx : dcache_metaArb_io_in_2_valid  ?  dcache_metaArb_io_in_2_bits_idx : dcache_metaArb_io_in_3_valid  ?  dcache_metaArb_io_in_3_bits_idx : dcache_metaArb_io_in_4_valid  ?  dcache_metaArb_io_in_4_bits_idx : dcache_metaArb_io_in_5_valid  ?  dcache_metaArb_io_in_5_bits_idx : dcache_metaArb_io_in_6_valid  ?  dcache_metaArb_io_in_6_bits_idx : dcache_metaArb_io_in_7_bits_idx ; 
    wire[21:0] dcache_metaArb_io_in_0_bits_data ; 
    wire dcache_metaArb_io_out_bits_way_en = dcache_metaArb_io_in_0_valid  ?  dcache_metaArb_io_in_0_bits_way_en : dcache_metaArb_io_in_1_valid  ?  dcache_metaArb_io_in_1_bits_way_en : dcache_metaArb_io_in_2_valid  ?  dcache_metaArb_io_in_2_bits_way_en : dcache_metaArb_io_in_3_valid  ?  dcache_metaArb_io_in_3_bits_way_en : dcache_metaArb_io_in_4_valid  ?  dcache_metaArb_io_in_4_bits_way_en : dcache_metaArb_io_in_5_valid  ?  dcache_metaArb_io_in_5_bits_way_en : dcache_metaArb_io_in_6_valid  ?  dcache_metaArb_io_in_6_bits_way_en : dcache_metaArb_io_in_7_bits_way_en ; 
  assign  dcache_metaArb_io_out_bits_data = dcache_metaArb_io_in_0_valid  ?  dcache_metaArb_io_in_0_bits_data : dcache_metaArb_io_in_1_valid  ?  dcache_metaArb_io_in_1_bits_data : dcache_metaArb_io_in_2_valid  ?  dcache_metaArb_io_in_2_bits_data : dcache_metaArb_io_in_3_valid  ?  dcache_metaArb_io_in_3_bits_data : dcache_metaArb_io_in_4_valid  ?  dcache_metaArb_io_in_4_bits_data : dcache_metaArb_io_in_5_valid  ?  dcache_metaArb_io_in_5_bits_data : dcache_metaArb_io_in_6_valid  ?  dcache_metaArb_io_in_6_bits_data : dcache_metaArb_io_in_7_bits_data ; 
    wire dcache__GEN_81 = dcache_metaArb_io_in_0_valid | dcache_metaArb_io_in_1_valid ; 
    wire dcache__GEN_82 = dcache__GEN_81 | dcache_metaArb_io_in_2_valid ; 
    wire dcache__GEN_83 = dcache__GEN_82 | dcache_metaArb_io_in_3_valid ; 
    wire dcache__GEN_84 = dcache__GEN_83 | dcache_metaArb_io_in_4_valid ; 
    wire dcache__GEN_85 = dcache__GEN_84 | dcache_metaArb_io_in_5_valid ; 
    wire dcache_metaArb_grant_1 = dcache_metaArb_io_in_0_valid ==1'h0; 
    wire dcache_metaArb_grant_2 = dcache__GEN_81 ==1'h0; 
    wire dcache_metaArb_grant_3 = dcache__GEN_82 ==1'h0; 
    wire dcache_metaArb_grant_4 = dcache__GEN_83 ==1'h0; 
    wire dcache_metaArb_grant_5 = dcache__GEN_84 ==1'h0; 
    wire dcache_metaArb_grant_6 = dcache__GEN_85 ==1'h0; 
    wire dcache_metaArb_grant_7 =( dcache__GEN_85 | dcache_metaArb_io_in_6_valid )==1'h0; 
    wire dcache_metaArb_io_in_0_ready = dcache_metaArb_io_out_ready &1'h1; 
    wire dcache_metaArb_io_in_1_ready = dcache_metaArb_grant_1 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_2_ready = dcache_metaArb_grant_2 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_3_ready = dcache_metaArb_grant_3 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_4_ready = dcache_metaArb_grant_4 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_5_ready = dcache_metaArb_grant_5 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_6_ready = dcache_metaArb_grant_6 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_in_7_ready = dcache_metaArb_grant_7 & dcache_metaArb_io_out_ready ; 
    wire dcache_metaArb_io_out_valid = dcache_metaArb_grant_7 ==1'h0| dcache_metaArb_io_in_7_valid ; 
    wire[21:0] dcache_tag_array_MPORT_data_0 ; 
    wire[5:0] dcache_tag_array_s1_meta_addr ; 
    wire dcache_tag_array_s1_meta_en ; 
    wire[21:0] dcache__s1_meta_uncorrected_WIRE = dcache_tag_array_s1_meta_data_0 ;  
    wire[5:0] dcache_tag_array_0_ext_R0_addr;
    wire dcache_tag_array_0_ext_R0_en;
    wire dcache_tag_array_0_ext_R0_clk;
    wire[21:0] dcache_tag_array_0_ext_R0_data;
    wire[5:0] dcache_tag_array_0_ext_W0_addr;
    wire dcache_tag_array_0_ext_W0_en;
    wire dcache_tag_array_0_ext_W0_clk;
    wire[21:0] dcache_tag_array_0_ext_W0_data;

    reg[21:0] dcache_tag_array_0_ext_Memory [0:63]; 
    reg dcache_tag_array_0_ext__R0_en_d0 ; reg[5:0] dcache_tag_array_0_ext__R0_addr_d0 ; 
  always @( posedge  dcache_tag_array_0_ext_R0_clk )
         begin  
             dcache_tag_array_0_ext__R0_en_d0  <= dcache_tag_array_0_ext_R0_en ; 
             dcache_tag_array_0_ext__R0_addr_d0  <= dcache_tag_array_0_ext_R0_addr ;
         end
  always @( posedge  dcache_tag_array_0_ext_W0_clk )
         begin 
             if ( dcache_tag_array_0_ext_W0_en &1'h1) 
                 dcache_tag_array_0_ext_Memory  [ dcache_tag_array_0_ext_W0_addr ]<= dcache_tag_array_0_ext_W0_data ;
         end
  assign  dcache_tag_array_0_ext_R0_data = dcache_tag_array_0_ext__R0_en_d0  ?  dcache_tag_array_0_ext_Memory [ dcache_tag_array_0_ext__R0_addr_d0 ]:22'bx;
    assign dcache_tag_array_0_ext_R0_addr = dcache_tag_array_s1_meta_addr;
    assign dcache_tag_array_0_ext_R0_en = dcache_tag_array_s1_meta_en;
    assign dcache_tag_array_0_ext_R0_clk = dcache_tag_array_s1_meta_clk;
    assign dcache_tag_array_s1_meta_data_0 = dcache_tag_array_0_ext_R0_data;
    assign dcache_tag_array_0_ext_W0_addr = dcache_tag_array_MPORT_addr;
    assign dcache_tag_array_0_ext_W0_en = dcache__GEN;
    assign dcache_tag_array_0_ext_W0_clk = dcache_tag_array_MPORT_clk;
    assign dcache_tag_array_0_ext_W0_data = dcache_tag_array_MPORT_data_0;
     
    wire dcache_tag_array_MPORT_en ; 
  assign  dcache__GEN = dcache_tag_array_MPORT_en & dcache_tag_array_MPORT_mask_0 ; 
    wire dcache_dataArb_io_out_valid ; 
    wire[11:0] dcache_dataArb_io_out_bits_addr ; 
    wire dcache_dataArb_io_out_bits_write ; 
    wire[63:0] dcache_dataArb_io_out_bits_wdata ; 
    wire dcache_dataArb_io_out_bits_wordMask ; 
    wire[7:0] dcache_dataArb_io_out_bits_eccMask ; 
    wire dcache_dataArb_io_out_bits_way_en ;  
    wire dcache_data_clock;
    wire dcache_data_reset;
    wire dcache_data_io_req_valid;
    wire[11:0] dcache_data_io_req_bits_addr;
    wire dcache_data_io_req_bits_write;
    wire[63:0] dcache_data_io_req_bits_wdata;
    wire dcache_data_io_req_bits_wordMask;
    wire[7:0] dcache_data_io_req_bits_eccMask;
    wire dcache_data_io_req_bits_way_en;
    wire[63:0] dcache_data_io_resp_0;

    wire[7:0] dcache_data__GEN ; 
    wire[63:0] dcache_data__GEN_0 ; 
    wire[63:0] dcache_data__data_arrays_0_ext_R0_data ; 
    wire[63:0] dcache_data_wWords_0 = dcache_data_io_req_bits_wdata ; 
    wire dcache_data_data_arrays_0_rdata_MPORT_clk = dcache_data_clock ; 
    wire dcache_data_data_arrays_0_rdata_data_clk = dcache_data_clock ; 
    wire dcache_data_rdata_valid = dcache_data_io_req_valid ; 
    wire dcache_data_eccMask_0 = dcache_data_io_req_bits_eccMask [0]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_0 = dcache_data_eccMask_0 ; 
    wire dcache_data_eccMask_1 = dcache_data_io_req_bits_eccMask [1]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_1 = dcache_data_eccMask_1 ; 
    wire dcache_data_eccMask_2 = dcache_data_io_req_bits_eccMask [2]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_2 = dcache_data_eccMask_2 ; 
    wire dcache_data_eccMask_3 = dcache_data_io_req_bits_eccMask [3]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_3 = dcache_data_eccMask_3 ; 
    wire dcache_data_eccMask_4 = dcache_data_io_req_bits_eccMask [4]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_4 = dcache_data_eccMask_4 ; 
    wire dcache_data_eccMask_5 = dcache_data_io_req_bits_eccMask [5]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_5 = dcache_data_eccMask_5 ; 
    wire dcache_data_eccMask_6 = dcache_data_io_req_bits_eccMask [6]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_6 = dcache_data_eccMask_6 ; 
    wire dcache_data_eccMask_7 = dcache_data_io_req_bits_eccMask [7]; 
    wire dcache_data_data_arrays_0_rdata_MPORT_mask_7 = dcache_data_eccMask_7 ; 
    wire[8:0] dcache_data_addr = dcache_data_io_req_bits_addr [11:3]; 
    wire[8:0] dcache_data_data_arrays_0_rdata_MPORT_addr = dcache_data_addr ; 
    wire dcache_data_data_arrays_0_rdata_MPORT_en ; 
    wire[8:0] dcache_data_data_arrays_0_rdata_data_addr ; 
    wire dcache_data_data_arrays_0_rdata_data_en ; 
    wire[8:0] dcache_data__rdata_data_WIRE = dcache_data_addr ;  
    wire[8:0] dcache_data_data_arrays_0_ext_R0_addr;
    wire dcache_data_data_arrays_0_ext_R0_en;
    wire dcache_data_data_arrays_0_ext_R0_clk;
    wire[63:0] dcache_data_data_arrays_0_ext_R0_data;
    wire[8:0] dcache_data_data_arrays_0_ext_W0_addr;
    wire dcache_data_data_arrays_0_ext_W0_en;
    wire dcache_data_data_arrays_0_ext_W0_clk;
    wire[63:0] dcache_data_data_arrays_0_ext_W0_data;
    wire[7:0] dcache_data_data_arrays_0_ext_W0_mask;

    reg[63:0] dcache_data_data_arrays_0_ext_Memory [0:511]; 
    reg dcache_data_data_arrays_0_ext__R0_en_d0 ; reg[8:0] dcache_data_data_arrays_0_ext__R0_addr_d0 ; 
  always @( posedge  dcache_data_data_arrays_0_ext_R0_clk )
         begin  
             dcache_data_data_arrays_0_ext__R0_en_d0  <= dcache_data_data_arrays_0_ext_R0_en ; 
             dcache_data_data_arrays_0_ext__R0_addr_d0  <= dcache_data_data_arrays_0_ext_R0_addr ;
         end
  always @( posedge  dcache_data_data_arrays_0_ext_W0_clk )
         begin 
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [0]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h0+:8]<= dcache_data_data_arrays_0_ext_W0_data [7:0];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [1]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h8+:8]<= dcache_data_data_arrays_0_ext_W0_data [15:8];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [2]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h10+:8]<= dcache_data_data_arrays_0_ext_W0_data [23:16];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [3]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h18+:8]<= dcache_data_data_arrays_0_ext_W0_data [31:24];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [4]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h20+:8]<= dcache_data_data_arrays_0_ext_W0_data [39:32];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [5]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h28+:8]<= dcache_data_data_arrays_0_ext_W0_data [47:40];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [6]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h30+:8]<= dcache_data_data_arrays_0_ext_W0_data [55:48];
             if ( dcache_data_data_arrays_0_ext_W0_en & dcache_data_data_arrays_0_ext_W0_mask [7]) 
                 dcache_data_data_arrays_0_ext_Memory  [ dcache_data_data_arrays_0_ext_W0_addr ][32'h38+:8]<= dcache_data_data_arrays_0_ext_W0_data [63:56];
         end
  assign  dcache_data_data_arrays_0_ext_R0_data = dcache_data_data_arrays_0_ext__R0_en_d0  ?  dcache_data_data_arrays_0_ext_Memory [ dcache_data_data_arrays_0_ext__R0_addr_d0 ]:64'bx;
    assign dcache_data_data_arrays_0_ext_R0_addr = dcache_data_data_arrays_0_rdata_data_addr;
    assign dcache_data_data_arrays_0_ext_R0_en = dcache_data_data_arrays_0_rdata_data_en;
    assign dcache_data_data_arrays_0_ext_R0_clk = dcache_data_data_arrays_0_rdata_data_clk;
    assign dcache_data__data_arrays_0_ext_R0_data = dcache_data_data_arrays_0_ext_R0_data;
    assign dcache_data_data_arrays_0_ext_W0_addr = dcache_data_data_arrays_0_rdata_MPORT_addr;
    assign dcache_data_data_arrays_0_ext_W0_en = dcache_data_data_arrays_0_rdata_MPORT_en;
    assign dcache_data_data_arrays_0_ext_W0_clk = dcache_data_data_arrays_0_rdata_MPORT_clk;
    assign dcache_data_data_arrays_0_ext_W0_data = dcache_data__GEN_0;
    assign dcache_data_data_arrays_0_ext_W0_mask = dcache_data__GEN;
     
    wire[7:0] dcache_data__rdata_WIRE_0 ; 
    wire[7:0] dcache_data__rdata_WIRE_1 ; 
    wire[7:0] dcache_data__rdata_WIRE_2 ; 
    wire[7:0] dcache_data__rdata_WIRE_3 ; 
    wire[7:0] dcache_data__rdata_WIRE_4 ; 
    wire[7:0] dcache_data__rdata_WIRE_5 ; 
    wire[7:0] dcache_data__rdata_WIRE_6 ; 
    wire[7:0] dcache_data__rdata_WIRE_7 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_0 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_1 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_2 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_3 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_4 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_5 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_6 ; 
    wire[7:0] dcache_data_data_arrays_0_rdata_MPORT_data_7 ; 
  assign  dcache_data__GEN_0 ={ dcache_data_data_arrays_0_rdata_MPORT_data_7 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_6 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_5 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_4 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_3 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_2 ,{ dcache_data_data_arrays_0_rdata_MPORT_data_1 , dcache_data_data_arrays_0_rdata_MPORT_data_0 }}}}}}}; 
  assign  dcache_data__GEN ={ dcache_data_data_arrays_0_rdata_MPORT_mask_7 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_6 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_5 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_4 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_3 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_2 ,{ dcache_data_data_arrays_0_rdata_MPORT_mask_1 , dcache_data_data_arrays_0_rdata_MPORT_mask_0 }}}}}}}; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_0 = dcache_data__data_arrays_0_ext_R0_data [7:0]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_1 = dcache_data__data_arrays_0_ext_R0_data [15:8]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_2 = dcache_data__data_arrays_0_ext_R0_data [23:16]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_3 = dcache_data__data_arrays_0_ext_R0_data [31:24]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_4 = dcache_data__data_arrays_0_ext_R0_data [39:32]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_5 = dcache_data__data_arrays_0_ext_R0_data [47:40]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_6 = dcache_data__data_arrays_0_ext_R0_data [55:48]; 
    wire[7:0] dcache_data_data_arrays_0_rdata_data_data_7 = dcache_data__data_arrays_0_ext_R0_data [63:56]; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_en = dcache_data_rdata_valid & dcache_data_io_req_bits_write ; 
    wire[7:0] dcache_data_rdata_wData_0 = dcache_data_wWords_0 [7:0]; 
  assign  dcache_data__rdata_WIRE_0 = dcache_data_rdata_wData_0 ; 
    wire[7:0] dcache_data_rdata_wData_1 = dcache_data_wWords_0 [15:8]; 
  assign  dcache_data__rdata_WIRE_1 = dcache_data_rdata_wData_1 ; 
    wire[7:0] dcache_data_rdata_wData_2 = dcache_data_wWords_0 [23:16]; 
  assign  dcache_data__rdata_WIRE_2 = dcache_data_rdata_wData_2 ; 
    wire[7:0] dcache_data_rdata_wData_3 = dcache_data_wWords_0 [31:24]; 
  assign  dcache_data__rdata_WIRE_3 = dcache_data_rdata_wData_3 ; 
    wire[7:0] dcache_data_rdata_wData_4 = dcache_data_wWords_0 [39:32]; 
  assign  dcache_data__rdata_WIRE_4 = dcache_data_rdata_wData_4 ; 
    wire[7:0] dcache_data_rdata_wData_5 = dcache_data_wWords_0 [47:40]; 
  assign  dcache_data__rdata_WIRE_5 = dcache_data_rdata_wData_5 ; 
    wire[7:0] dcache_data_rdata_wData_6 = dcache_data_wWords_0 [55:48]; 
  assign  dcache_data__rdata_WIRE_6 = dcache_data_rdata_wData_6 ; 
    wire[7:0] dcache_data_rdata_wData_7 = dcache_data_wWords_0 [63:56]; 
  assign  dcache_data__rdata_WIRE_7 = dcache_data_rdata_wData_7 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_0 = dcache_data__rdata_WIRE_0 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_1 = dcache_data__rdata_WIRE_1 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_2 = dcache_data__rdata_WIRE_2 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_3 = dcache_data__rdata_WIRE_3 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_4 = dcache_data__rdata_WIRE_4 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_5 = dcache_data__rdata_WIRE_5 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_6 = dcache_data__rdata_WIRE_6 ; 
  assign  dcache_data_data_arrays_0_rdata_MPORT_data_7 = dcache_data__rdata_WIRE_7 ; 
  assign  dcache_data_data_arrays_0_rdata_data_en = dcache_data_rdata_valid & dcache_data_io_req_bits_write ==1'h0; 
  assign  dcache_data_data_arrays_0_rdata_data_addr = dcache_data__rdata_data_WIRE ; 
    wire[15:0] dcache_data_rdata_lo_lo ={ dcache_data_data_arrays_0_rdata_data_data_1 , dcache_data_data_arrays_0_rdata_data_data_0 }; 
    wire[15:0] dcache_data_rdata_lo_hi ={ dcache_data_data_arrays_0_rdata_data_data_3 , dcache_data_data_arrays_0_rdata_data_data_2 }; 
    wire[31:0] dcache_data_rdata_lo ={ dcache_data_rdata_lo_hi , dcache_data_rdata_lo_lo }; 
    wire[15:0] dcache_data_rdata_hi_lo ={ dcache_data_data_arrays_0_rdata_data_data_5 , dcache_data_data_arrays_0_rdata_data_data_4 }; 
    wire[15:0] dcache_data_rdata_hi_hi ={ dcache_data_data_arrays_0_rdata_data_data_7 , dcache_data_data_arrays_0_rdata_data_data_6 }; 
    wire[31:0] dcache_data_rdata_hi ={ dcache_data_rdata_hi_hi , dcache_data_rdata_hi_lo }; 
    wire[63:0] dcache_data_rdata_0_0 ={ dcache_data_rdata_hi , dcache_data_rdata_lo }; 
  assign  dcache_data_io_resp_0 = dcache_data_rdata_0_0 ;
    assign dcache_data_clock = dcache_clock;
    assign dcache_data_reset = dcache_reset;
    assign dcache_data_io_req_valid = dcache_dataArb_io_out_valid;
    assign dcache_data_io_req_bits_addr = dcache_dataArb_io_out_bits_addr;
    assign dcache_data_io_req_bits_write = dcache_dataArb_io_out_bits_write;
    assign dcache_data_io_req_bits_wdata = dcache_dataArb_io_out_bits_wdata;
    assign dcache_data_io_req_bits_wordMask = dcache_dataArb_io_out_bits_wordMask;
    assign dcache_data_io_req_bits_eccMask = dcache_dataArb_io_out_bits_eccMask;
    assign dcache_data_io_req_bits_way_en = dcache_dataArb_io_out_bits_way_en;
    assign dcache_s1_all_data_ways_0 = dcache_data_io_resp_0;
     
    wire dcache_pstore_drain ; 
    wire[63:0] dcache_tl_d_data_encoded ; 
    wire[63:0] dcache_dataArb_io_in_2_bits_wdata = dcache_dataArb_io_in_1_bits_wdata ; 
    wire[63:0] dcache_dataArb_io_in_3_bits_wdata = dcache_dataArb_io_in_1_bits_wdata ; 
    wire dcache_dataArb_io_in_2_valid ; 
    wire[11:0] dcache_dataArb_io_in_2_bits_addr ; 
    wire[11:0] dcache_dataArb_io_in_3_bits_addr ; 
    wire dcache_dataArb_io_in_1_valid ; 
    wire[11:0] dcache_dataArb_io_in_1_bits_addr ; 
    wire dcache_dataArb_io_in_1_bits_write ; 
    wire dcache_dataArb_io_in_1_bits_way_en ; 
    wire dcache_dataArb_io_in_0_valid ; 
    wire[11:0] dcache_dataArb_io_in_0_bits_addr ; 
    wire[1:0] dcache_dataArb_io_chosen = dcache_dataArb_io_in_0_valid  ? 2'h0: dcache_dataArb_io_in_1_valid  ? 2'h1: dcache_dataArb_io_in_2_valid  ? 2'h2:2'h3; 
    wire dcache_dataArb_io_in_0_bits_write ; 
  assign  dcache_dataArb_io_out_bits_addr = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_addr : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_addr : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_addr : dcache_dataArb_io_in_3_bits_addr ; 
    wire[63:0] dcache_dataArb_io_in_0_bits_wdata ; 
  assign  dcache_dataArb_io_out_bits_write = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_write : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_write : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_write : dcache_dataArb_io_in_3_bits_write ; 
    wire dcache_dataArb_io_in_0_bits_wordMask ; 
  assign  dcache_dataArb_io_out_bits_wdata = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_wdata : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_wdata : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_wdata : dcache_dataArb_io_in_3_bits_wdata ; 
    wire[7:0] dcache_dataArb_io_in_0_bits_eccMask ; 
  assign  dcache_dataArb_io_out_bits_wordMask = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_wordMask : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_wordMask : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_wordMask : dcache_dataArb_io_in_3_bits_wordMask ; 
    wire dcache_dataArb_io_in_0_bits_way_en ; 
  assign  dcache_dataArb_io_out_bits_eccMask = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_eccMask : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_eccMask : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_eccMask : dcache_dataArb_io_in_3_bits_eccMask ; 
  assign  dcache_dataArb_io_out_bits_way_en = dcache_dataArb_io_in_0_valid  ?  dcache_dataArb_io_in_0_bits_way_en : dcache_dataArb_io_in_1_valid  ?  dcache_dataArb_io_in_1_bits_way_en : dcache_dataArb_io_in_2_valid  ?  dcache_dataArb_io_in_2_bits_way_en : dcache_dataArb_io_in_3_bits_way_en ; 
    wire dcache__GEN_86 = dcache_dataArb_io_in_0_valid | dcache_dataArb_io_in_1_valid ; 
    wire dcache_dataArb_grant_1 = dcache_dataArb_io_in_0_valid ==1'h0; 
    wire dcache_dataArb_grant_2 = dcache__GEN_86 ==1'h0; 
    wire dcache_dataArb_grant_3 =( dcache__GEN_86 | dcache_dataArb_io_in_2_valid )==1'h0; 
    wire dcache_dataArb_io_in_0_ready = dcache_dataArb_io_out_ready &1'h1; 
    wire dcache_dataArb_io_in_1_ready = dcache_dataArb_grant_1 & dcache_dataArb_io_out_ready ; 
    wire dcache_dataArb_io_in_2_ready = dcache_dataArb_grant_2 & dcache_dataArb_io_out_ready ; 
    wire dcache_dataArb_io_in_3_ready = dcache_dataArb_grant_3 & dcache_dataArb_io_out_ready ; 
    wire dcache_dataArb_io_in_3_valid ; 
  assign  dcache_dataArb_io_out_valid = dcache_dataArb_grant_3 ==1'h0| dcache_dataArb_io_in_3_valid ; 
  assign  dcache_nodeOut_a_deq_valid = dcache_tl_out_a_valid ; 
  assign  dcache_nodeOut_a_deq_bits_opcode = dcache_tl_out_a_bits_opcode ; 
  assign  dcache_nodeOut_a_deq_bits_param = dcache_tl_out_a_bits_param ; 
  assign  dcache_nodeOut_a_deq_bits_size = dcache_tl_out_a_bits_size ; 
  assign  dcache_nodeOut_a_deq_bits_source = dcache_tl_out_a_bits_source ; 
  assign  dcache_nodeOut_a_deq_bits_address = dcache_tl_out_a_bits_address ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable = dcache_tl_out_a_bits_user_amba_prot_bufferable ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable = dcache_tl_out_a_bits_user_amba_prot_modifiable ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc = dcache_tl_out_a_bits_user_amba_prot_readalloc ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc = dcache_tl_out_a_bits_user_amba_prot_writealloc ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_privileged = dcache_tl_out_a_bits_user_amba_prot_privileged ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_secure = dcache_tl_out_a_bits_user_amba_prot_secure ; 
  assign  dcache_nodeOut_a_deq_bits_user_amba_prot_fetch = dcache_tl_out_a_bits_user_amba_prot_fetch ; 
  assign  dcache_nodeOut_a_deq_bits_mask = dcache_tl_out_a_bits_mask ; 
  assign  dcache_nodeOut_a_deq_bits_data = dcache_tl_out_a_bits_data ; 
  assign  dcache_nodeOut_a_deq_bits_corrupt = dcache_tl_out_a_bits_corrupt ; 
    wire dcache_tl_out_a_ready = dcache_nodeOut_a_deq_ready ; 
    wire dcache_nodeOut_a_valid = dcache_nodeOut_a_deq_valid ; 
    wire[2:0] dcache_nodeOut_a_bits_opcode = dcache_nodeOut_a_deq_bits_opcode ; 
    wire[2:0] dcache_nodeOut_a_bits_param = dcache_nodeOut_a_deq_bits_param ; 
    wire[3:0] dcache_nodeOut_a_bits_size = dcache_nodeOut_a_deq_bits_size ; 
    wire dcache_nodeOut_a_bits_source = dcache_nodeOut_a_deq_bits_source ; 
    wire[31:0] dcache_nodeOut_a_bits_address = dcache_nodeOut_a_deq_bits_address ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_bufferable = dcache_nodeOut_a_deq_bits_user_amba_prot_bufferable ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_modifiable = dcache_nodeOut_a_deq_bits_user_amba_prot_modifiable ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_readalloc = dcache_nodeOut_a_deq_bits_user_amba_prot_readalloc ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_writealloc = dcache_nodeOut_a_deq_bits_user_amba_prot_writealloc ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_privileged = dcache_nodeOut_a_deq_bits_user_amba_prot_privileged ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_secure = dcache_nodeOut_a_deq_bits_user_amba_prot_secure ; 
    wire dcache_nodeOut_a_bits_user_amba_prot_fetch = dcache_nodeOut_a_deq_bits_user_amba_prot_fetch ; 
    wire[7:0] dcache_nodeOut_a_bits_mask = dcache_nodeOut_a_deq_bits_mask ; 
    wire[63:0] dcache_nodeOut_a_bits_data = dcache_nodeOut_a_deq_bits_data ; 
    wire dcache__io_cpu_req_ready_output ; 
    wire dcache_nodeOut_a_bits_corrupt = dcache_nodeOut_a_deq_bits_corrupt ; 
    reg dcache_s1_valid ; 
    wire dcache_nodeOut_b_ready ; 
    wire dcache__GEN_87 = dcache_nodeOut_b_ready & dcache_nodeOut_b_valid ; 
    reg dcache_s1_probe ; 
    wire dcache__GEN_88 = dcache_nodeOut_b_ready & dcache_nodeOut_b_valid ; reg[2:0] dcache_probe_bits_opcode ; reg[1:0] dcache_probe_bits_param ; reg[3:0] dcache_probe_bits_size ; 
    wire[3:0] dcache_nackResponseMessage_size = dcache_probe_bits_size ; 
    wire[3:0] dcache_cleanReleaseMessage_size = dcache_probe_bits_size ; 
    wire[3:0] dcache_dirtyReleaseMessage_size = dcache_probe_bits_size ; 
    reg dcache_probe_bits_source ; 
    wire dcache_nodeOut_c_bits_source = dcache_probe_bits_source ; 
    wire dcache_nackResponseMessage_source = dcache_probe_bits_source ; 
    wire dcache_cleanReleaseMessage_source = dcache_probe_bits_source ; 
    wire dcache_dirtyReleaseMessage_source = dcache_probe_bits_source ; reg[31:0] dcache_probe_bits_address ; 
    wire[31:0] dcache_nodeOut_c_bits_address = dcache_probe_bits_address ; 
    wire[31:0] dcache_nackResponseMessage_address = dcache_probe_bits_address ; 
    wire[31:0] dcache_cleanReleaseMessage_address = dcache_probe_bits_address ; 
    wire[31:0] dcache_dirtyReleaseMessage_address = dcache_probe_bits_address ; reg[7:0] dcache_probe_bits_mask ; reg[63:0] dcache_probe_bits_data ; 
    reg dcache_probe_bits_corrupt ; 
    wire dcache_s1_valid_masked = dcache_s1_valid & dcache_io_cpu_s1_kill ==1'h0; 
    wire dcache_s1_nack ; 
    wire dcache_s1_valid_not_nacked = dcache_s1_valid & dcache_s1_nack ==1'h0; 
    reg dcache_s1_tlb_req_valid ; 
    reg dcache_s2_tlb_req_valid ; 
    wire dcache_s0_clk_en = dcache_metaArb_io_out_valid & dcache_metaArb_io_out_bits_write ==1'h0; 
    wire[33:0] dcache_s0_req_addr ={ dcache_metaArb_io_out_bits_addr [33:6], dcache_io_cpu_req_bits_addr [5:0]}; 
    wire dcache_s0_req_phys = dcache_metaArb_io_in_7_ready ==1'h0 ? 1'h1: dcache_io_cpu_req_bits_phys ; reg[33:0] dcache_s1_req_addr ; 
  assign  dcache_pma_checker_io_req_bits_vaddr = dcache_s1_req_addr ; reg[5:0] dcache_s1_req_tag ; reg[4:0] dcache_s1_req_cmd ; 
  assign  dcache_pma_checker_io_req_bits_cmd = dcache_s1_req_cmd ; reg[1:0] dcache_s1_req_size ; 
  assign  dcache_pma_checker_io_req_bits_size = dcache_s1_req_size ; 
    wire[1:0] dcache_s1_mask_xwr_size = dcache_s1_req_size ; 
    reg dcache_s1_req_signed ; reg[1:0] dcache_s1_req_dprv ; 
  assign  dcache_pma_checker_io_req_bits_prv = dcache_s1_req_dprv ; 
    reg dcache_s1_req_dv ; 
    wire dcache_pma_checker_io_req_bits_v = dcache_s1_req_dv ; 
    reg dcache_s1_req_phys ; 
    reg dcache_s1_req_no_alloc ; 
    reg dcache_s1_req_no_xcpt ; reg[63:0] dcache_s1_req_data ; reg[7:0] dcache_s1_req_mask ; 
    wire[33:0] dcache_s1_vaddr ={ dcache_s1_req_addr [33:12], dcache_s1_req_addr [11:0]}; 
    wire dcache__GEN_89 =( dcache__tlb_port_req_ready_output & dcache_tlb_port_req_valid )==1'h0; 
    wire dcache_s0_tlb_req_passthrough = dcache__GEN_89  ?  dcache_s0_req_phys : dcache_tlb_port_req_bits_passthrough ; 
    wire[33:0] dcache_s0_tlb_req_vaddr = dcache__GEN_89  ?  dcache_s0_req_addr : dcache_tlb_port_req_bits_vaddr ; 
    wire[1:0] dcache_s0_tlb_req_size = dcache__GEN_89  ?  dcache_s0_req_size : dcache_tlb_port_req_bits_size ; 
    wire[4:0] dcache_s0_tlb_req_cmd = dcache__GEN_89  ?  dcache_s0_req_cmd : dcache_tlb_port_req_bits_cmd ; 
    wire[1:0] dcache_s0_tlb_req_prv = dcache__GEN_89  ?  dcache_s0_req_dprv : dcache_tlb_port_req_bits_prv ; 
    wire dcache_s0_tlb_req_v = dcache__GEN_89  ?  dcache_s0_req_dv : dcache_tlb_port_req_bits_v ; 
    wire dcache__GEN_90 = dcache_s0_clk_en | dcache_tlb_port_req_valid ; reg[33:0] dcache_s1_tlb_req_vaddr ; 
  assign  dcache_tlb_io_req_bits_vaddr = dcache_s1_tlb_req_vaddr ; 
    reg dcache_s1_tlb_req_passthrough ; 
  assign  dcache_tlb_io_req_bits_passthrough = dcache_s1_tlb_req_passthrough ; reg[1:0] dcache_s1_tlb_req_size ; 
  assign  dcache_tlb_io_req_bits_size = dcache_s1_tlb_req_size ; reg[4:0] dcache_s1_tlb_req_cmd ; 
  assign  dcache_tlb_io_req_bits_cmd = dcache_s1_tlb_req_cmd ; reg[1:0] dcache_s1_tlb_req_prv ; 
  assign  dcache_tlb_io_req_bits_prv = dcache_s1_tlb_req_prv ; 
    reg dcache_s1_tlb_req_v ; 
    wire dcache_tlb_io_req_bits_v = dcache_s1_tlb_req_v ; 
    wire dcache_s1_read = dcache_s1_req_cmd ==5'h0| dcache_s1_req_cmd ==5'h10| dcache_s1_req_cmd ==5'h6| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF; 
    wire dcache_s1_write = dcache_s1_req_cmd ==5'h1| dcache_s1_req_cmd ==5'h11| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF; 
    wire dcache_s1_readwrite = dcache_s1_read | dcache_s1_write ; 
    wire dcache_s1_sfence = dcache_s1_req_cmd ==5'h14| dcache_s1_req_cmd ==5'h15| dcache_s1_req_cmd ==5'h16; 
    wire dcache_s1_flush_line = dcache_s1_req_cmd ==5'h5& dcache_s1_req_size [0]; 
    reg dcache_s1_flush_valid ; 
    reg dcache_flushed ; 
    reg dcache_flushing ; reg[33:0] dcache_flushing_req_addr ; reg[5:0] dcache_flushing_req_tag ; reg[4:0] dcache_flushing_req_cmd ; reg[1:0] dcache_flushing_req_size ; 
    reg dcache_flushing_req_signed ; reg[1:0] dcache_flushing_req_dprv ; 
    reg dcache_flushing_req_dv ; 
    reg dcache_flushing_req_phys ; 
    reg dcache_flushing_req_no_alloc ; 
    reg dcache_flushing_req_no_xcpt ; reg[63:0] dcache_flushing_req_data ; reg[7:0] dcache_flushing_req_mask ; 
    reg dcache_cached_grant_wait ; 
    reg dcache_resetting ; 
  assign  dcache_metaArb_io_in_0_valid = dcache_resetting ; reg[5:0] dcache_flushCounter ; 
  assign  dcache_metaArb_io_in_5_bits_idx = dcache_flushCounter ; 
    reg dcache_release_ack_wait ; reg[31:0] dcache_release_ack_addr ; reg[3:0] dcache_release_state ; reg[1:0] dcache_refill_way ; 
    wire dcache_inWriteback = dcache_release_state ==4'h1| dcache_release_state ==4'h2; 
    reg dcache_uncachedInFlight_0 ; reg[33:0] dcache_uncachedReqs_0_addr ; 
    wire[33:0] dcache_uncachedResp_addr = dcache_uncachedReqs_0_addr ; reg[5:0] dcache_uncachedReqs_0_tag ; 
    wire[5:0] dcache_uncachedResp_tag = dcache_uncachedReqs_0_tag ; reg[4:0] dcache_uncachedReqs_0_cmd ; 
    wire[4:0] dcache_uncachedResp_cmd = dcache_uncachedReqs_0_cmd ; reg[1:0] dcache_uncachedReqs_0_size ; 
    wire[1:0] dcache_uncachedResp_size = dcache_uncachedReqs_0_size ; 
    reg dcache_uncachedReqs_0_signed ; 
    wire dcache_uncachedResp_signed = dcache_uncachedReqs_0_signed ; reg[1:0] dcache_uncachedReqs_0_dprv ; 
    wire[1:0] dcache_uncachedResp_dprv = dcache_uncachedReqs_0_dprv ; 
    reg dcache_uncachedReqs_0_dv ; 
    wire dcache_uncachedResp_dv = dcache_uncachedReqs_0_dv ; 
    reg dcache_uncachedReqs_0_phys ; 
    wire dcache_uncachedResp_phys = dcache_uncachedReqs_0_phys ; 
    reg dcache_uncachedReqs_0_no_alloc ; 
    wire dcache_uncachedResp_no_alloc = dcache_uncachedReqs_0_no_alloc ; 
    reg dcache_uncachedReqs_0_no_xcpt ; 
    wire dcache_uncachedResp_no_xcpt = dcache_uncachedReqs_0_no_xcpt ; reg[63:0] dcache_uncachedReqs_0_data ; 
    wire[63:0] dcache_uncachedResp_data = dcache_uncachedReqs_0_data ; reg[7:0] dcache_uncachedReqs_0_mask ; 
    wire[7:0] dcache_uncachedResp_mask = dcache_uncachedReqs_0_mask ; 
    wire dcache_s0_read = dcache_io_cpu_req_bits_cmd ==5'h0| dcache_io_cpu_req_bits_cmd ==5'h10| dcache_io_cpu_req_bits_cmd ==5'h6| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF; 
    wire dcache_dataArb_io_in_3_valid_res =( dcache_io_cpu_req_bits_cmd ==5'h1| dcache_io_cpu_req_bits_cmd ==5'h3)==1'h0| dcache_io_cpu_req_bits_size <2'h0; 
    wire dcache__GEN_91 =(( dcache_io_cpu_req_bits_cmd ==5'h0| dcache_io_cpu_req_bits_cmd ==5'h10| dcache_io_cpu_req_bits_cmd ==5'h6| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF|( dcache_io_cpu_req_bits_cmd ==5'h1| dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF)&( dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_size <2'h0))==1'h0| dcache_dataArb_io_in_3_valid_res )==1'h0; 
  assign  dcache_dataArb_io_in_3_valid = dcache_io_cpu_req_valid & dcache_dataArb_io_in_3_valid_res ; 
    wire[33:0] dcache__GEN_92 ={ dcache_io_cpu_req_bits_addr [33:12], dcache_io_cpu_req_bits_addr [11:0]}; 
  assign  dcache_dataArb_io_in_3_bits_addr = dcache__GEN_92 [11:0]; 
    wire dcache__GEN_93 = dcache_dataArb_io_in_3_ready & dcache_io_cpu_req_valid &( dcache_io_cpu_req_bits_cmd ==5'h0| dcache_io_cpu_req_bits_cmd ==5'h10| dcache_io_cpu_req_bits_cmd ==5'h6| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF|( dcache_io_cpu_req_bits_cmd ==5'h1| dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF)&( dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_size <2'h0)); 
    reg dcache_s1_did_read ; 
    reg dcache_s1_read_mask ; 
  assign  dcache_metaArb_io_in_7_bits_idx = dcache_dataArb_io_in_3_bits_addr [11:6]; 
    wire dcache_s1_cmd_uses_tlb = dcache_s1_readwrite | dcache_s1_flush_line | dcache_s1_req_cmd ==5'h17; 
  assign  dcache_tlb_io_kill = dcache_io_cpu_s2_kill | dcache_s2_tlb_req_valid & dcache_tlb_port_s2_kill ; 
  assign  dcache_tlb_io_req_valid = dcache_s1_tlb_req_valid | dcache_s1_valid & dcache_io_cpu_s1_kill ==1'h0& dcache_s1_cmd_uses_tlb ; 
    wire dcache__GEN_94 = dcache_tlb_io_req_ready ==1'h0& dcache_tlb_io_ptw_resp_valid ==1'h0& dcache_io_cpu_req_bits_phys ==1'h0 ? 1'h0: dcache_metaArb_io_in_7_ready ==1'h0 ? 1'h0: dcache_dataArb_io_in_3_ready ==1'h0& dcache_s0_read  ? 1'h0: dcache_release_state ==4'h0& dcache_cached_grant_wait ==1'h0& dcache_s1_nack ==1'h0; 
  assign  dcache_tlb_io_sfence_valid = dcache_s1_valid & dcache_io_cpu_s1_kill ==1'h0& dcache_s1_sfence ; 
    wire dcache_tlb_io_sfence_bits_rs1 = dcache_s1_req_size [0]; 
    wire dcache_tlb_io_sfence_bits_rs2 = dcache_s1_req_size [1]; 
    wire dcache_tlb_io_sfence_bits_asid = dcache_io_cpu_s1_data_data [0]; 
    wire[32:0] dcache_tlb_io_sfence_bits_addr = dcache_s1_req_addr [32:0]; 
    wire dcache_tlb_io_sfence_bits_hv = dcache_s1_req_cmd ==5'h15; 
    wire dcache_tlb_io_sfence_bits_hg = dcache_s1_req_cmd ==5'h16; 
    wire[31:0] dcache_s1_paddr ={ dcache_s1_tlb_req_valid  ?  dcache_s1_req_addr [31:12]: dcache_tlb_io_resp_paddr [31:12], dcache_s1_req_addr [11:0]}; 
  assign  dcache_tag_array_MPORT_en = dcache_metaArb_io_out_valid & dcache_metaArb_io_out_bits_write ; 
  assign  dcache_tag_array_MPORT_data_0 = dcache__GEN_80 ; 
  assign  dcache_tag_array_s1_meta_en = dcache_metaArb_io_out_valid & dcache_metaArb_io_out_bits_write ==1'h0; 
  assign  dcache_tag_array_s1_meta_addr = dcache__s1_meta_WIRE ; 
    wire[19:0] dcache_s1_meta_uncorrected_0_tag = dcache__s1_meta_uncorrected_WIRE [19:0]; 
    wire[1:0] dcache_s1_meta_uncorrected_0_coh_state = dcache__s1_meta_uncorrected_WIRE [21:20]; 
    wire[19:0] dcache_s1_tag = dcache_s1_paddr [31:12]; 
    wire dcache_s1_hit_way = dcache_s1_meta_uncorrected_0_coh_state >2'h0& dcache_s1_meta_uncorrected_0_tag == dcache_s1_tag ; 
    wire[1:0] dcache__s1_meta_hit_state_WIRE = dcache_s1_meta_uncorrected_0_tag == dcache_s1_tag & dcache_s1_flush_valid ==1'h0 ?  dcache_s1_meta_uncorrected_0_coh_state :2'h0; 
    wire[1:0] dcache_s1_hit_state_state = dcache__s1_meta_hit_state_WIRE ; 
    wire[15:0] dcache_tl_d_data_encoded_lo_lo ={ dcache_nodeOut_d_bits_data [15:8], dcache_nodeOut_d_bits_data [7:0]}; 
    wire[15:0] dcache_tl_d_data_encoded_lo_hi ={ dcache_nodeOut_d_bits_data [31:24], dcache_nodeOut_d_bits_data [23:16]}; 
    wire[31:0] dcache_tl_d_data_encoded_lo ={ dcache_tl_d_data_encoded_lo_hi , dcache_tl_d_data_encoded_lo_lo }; 
    wire[15:0] dcache_tl_d_data_encoded_hi_lo ={ dcache_nodeOut_d_bits_data [47:40], dcache_nodeOut_d_bits_data [39:32]}; 
    wire[15:0] dcache_tl_d_data_encoded_hi_hi ={ dcache_nodeOut_d_bits_data [63:56], dcache_nodeOut_d_bits_data [55:48]}; 
    wire[31:0] dcache_tl_d_data_encoded_hi ={ dcache_tl_d_data_encoded_hi_hi , dcache_tl_d_data_encoded_hi_lo }; 
  assign  dcache_dataArb_io_in_1_bits_wdata = dcache_tl_d_data_encoded ; 
    wire[63:0] dcache_s1_all_data_ways_1 = dcache_tl_d_data_encoded ; 
    wire[63:0] dcache_s2_data_s1_way_words_0_0 = dcache_s1_all_data_ways_0 ; 
    wire[63:0] dcache_s2_data_s1_way_words_1_0 = dcache_s1_all_data_ways_1 ; 
    wire dcache_s1_mask_xwr_upper = dcache_s1_req_addr [0]| dcache_s1_mask_xwr_size >=2'h1; 
    wire dcache_s1_mask_xwr_lower = dcache_s1_req_addr [0] ? 1'h0:1'h1; 
    wire[1:0] dcache__GEN_95 ={ dcache_s1_mask_xwr_upper , dcache_s1_mask_xwr_lower }; 
    wire[1:0] dcache_s1_mask_xwr_upper_1 =( dcache_s1_req_addr [1] ?  dcache__GEN_95 :2'h0)|( dcache_s1_mask_xwr_size >=2'h2 ? 2'h3:2'h0); 
    wire[1:0] dcache_s1_mask_xwr_lower_1 = dcache_s1_req_addr [1] ? 2'h0: dcache__GEN_95 ; 
    wire[3:0] dcache__GEN_96 ={ dcache_s1_mask_xwr_upper_1 , dcache_s1_mask_xwr_lower_1 }; 
    wire[3:0] dcache_s1_mask_xwr_upper_2 =( dcache_s1_req_addr [2] ?  dcache__GEN_96 :4'h0)|( dcache_s1_mask_xwr_size >=2'h3 ? 4'hF:4'h0); 
    wire[3:0] dcache_s1_mask_xwr_lower_2 = dcache_s1_req_addr [2] ? 4'h0: dcache__GEN_96 ; 
    wire[7:0] dcache_s1_mask_xwr ={ dcache_s1_mask_xwr_upper_2 , dcache_s1_mask_xwr_lower_2 }; 
    wire[7:0] dcache_s1_mask = dcache_s1_req_cmd ==5'h11 ?  dcache_io_cpu_s1_data_mask : dcache_s1_mask_xwr ; 
    wire dcache__GEN_97 =(( dcache_s1_valid_masked & dcache_s1_req_cmd ==5'h11)==1'h0|(&( dcache_s1_mask_xwr |~ dcache_io_cpu_s1_data_mask )))==1'h0; 
    reg dcache_s2_valid ; 
    wire dcache__io_cpu_s2_xcpt_ae_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_ae_st_output ; 
    wire[1:0] dcache_s2_valid_no_xcpt_lo_lo ={ dcache__io_cpu_s2_xcpt_ae_ld_output , dcache__io_cpu_s2_xcpt_ae_st_output }; 
    wire dcache__io_cpu_s2_xcpt_gf_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_gf_st_output ; 
    wire[1:0] dcache_s2_valid_no_xcpt_lo_hi ={ dcache__io_cpu_s2_xcpt_gf_ld_output , dcache__io_cpu_s2_xcpt_gf_st_output }; 
    wire[3:0] dcache_s2_valid_no_xcpt_lo ={ dcache_s2_valid_no_xcpt_lo_hi , dcache_s2_valid_no_xcpt_lo_lo }; 
    wire dcache__io_cpu_s2_xcpt_pf_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_pf_st_output ; 
    wire[1:0] dcache_s2_valid_no_xcpt_hi_lo ={ dcache__io_cpu_s2_xcpt_pf_ld_output , dcache__io_cpu_s2_xcpt_pf_st_output }; 
    wire dcache__io_cpu_s2_xcpt_ma_ld_output ; 
    wire dcache__io_cpu_s2_xcpt_ma_st_output ; 
    wire[1:0] dcache_s2_valid_no_xcpt_hi_hi ={ dcache__io_cpu_s2_xcpt_ma_ld_output , dcache__io_cpu_s2_xcpt_ma_st_output }; 
    wire[3:0] dcache_s2_valid_no_xcpt_hi ={ dcache_s2_valid_no_xcpt_hi_hi , dcache_s2_valid_no_xcpt_hi_lo }; 
    wire dcache_s2_valid_no_xcpt = dcache_s2_valid &(|{ dcache_s2_valid_no_xcpt_hi , dcache_s2_valid_no_xcpt_lo })==1'h0; 
    reg dcache_s2_probe ; 
    wire dcache_releaseInFlight = dcache_s1_probe | dcache_s2_probe |(| dcache_release_state ); 
    reg dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_not_nacked_in_s1 = dcache_s2_valid & dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_masked = dcache_s2_valid_no_xcpt & dcache_s2_not_nacked_in_s1 ; 
    wire dcache_s2_valid_not_killed = dcache_s2_valid_masked & dcache_io_cpu_s2_kill ==1'h0; reg[33:0] dcache_s2_req_addr ; reg[5:0] dcache_s2_req_tag ; reg[4:0] dcache_s2_req_cmd ; reg[1:0] dcache_s2_req_size ; 
    wire[1:0] dcache_size = dcache_s2_req_size ; 
    reg dcache_s2_req_signed ; reg[1:0] dcache_s2_req_dprv ; 
    reg dcache_s2_req_dv ; 
    reg dcache_s2_req_phys ; 
    reg dcache_s2_req_no_alloc ; 
    reg dcache_s2_req_no_xcpt ; reg[63:0] dcache_s2_req_data ; reg[7:0] dcache_s2_req_mask ; 
    wire dcache_s2_cmd_flush_all = dcache_s2_req_cmd ==5'h5& dcache_s2_req_size [0]==1'h0; 
    wire dcache_s2_cmd_flush_line = dcache_s2_req_cmd ==5'h5& dcache_s2_req_size [0]; 
    reg dcache_s2_tlb_xcpt_miss ; reg[31:0] dcache_s2_tlb_xcpt_paddr ; reg[33:0] dcache_s2_tlb_xcpt_gpa ; 
    reg dcache_s2_tlb_xcpt_gpa_is_pte ; 
    reg dcache_s2_tlb_xcpt_pf_ld ; 
    reg dcache_s2_tlb_xcpt_pf_st ; 
    reg dcache_s2_tlb_xcpt_pf_inst ; 
    reg dcache_s2_tlb_xcpt_gf_ld ; 
    reg dcache_s2_tlb_xcpt_gf_st ; 
    reg dcache_s2_tlb_xcpt_gf_inst ; 
    reg dcache_s2_tlb_xcpt_ae_ld ; 
    reg dcache_s2_tlb_xcpt_ae_st ; 
    reg dcache_s2_tlb_xcpt_ae_inst ; 
    reg dcache_s2_tlb_xcpt_ma_ld ; 
    reg dcache_s2_tlb_xcpt_ma_st ; 
    reg dcache_s2_tlb_xcpt_ma_inst ; 
    reg dcache_s2_tlb_xcpt_cacheable ; 
    reg dcache_s2_tlb_xcpt_must_alloc ; 
    reg dcache_s2_tlb_xcpt_prefetchable ; 
    reg dcache_s2_pma_miss ; reg[31:0] dcache_s2_pma_paddr ; reg[33:0] dcache_s2_pma_gpa ; 
    reg dcache_s2_pma_gpa_is_pte ; 
    reg dcache_s2_pma_pf_ld ; 
    reg dcache_s2_pma_pf_st ; 
    reg dcache_s2_pma_pf_inst ; 
    reg dcache_s2_pma_gf_ld ; 
    reg dcache_s2_pma_gf_st ; 
    reg dcache_s2_pma_gf_inst ; 
    reg dcache_s2_pma_ae_ld ; 
    reg dcache_s2_pma_ae_st ; 
    reg dcache_s2_pma_ae_inst ; 
    reg dcache_s2_pma_ma_ld ; 
    reg dcache_s2_pma_ma_st ; 
    reg dcache_s2_pma_ma_inst ; 
    reg dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_bufferable = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_modifiable = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_readalloc = dcache_s2_pma_cacheable ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_writealloc = dcache_s2_pma_cacheable ; 
    reg dcache_s2_pma_must_alloc ; 
    reg dcache_s2_pma_prefetchable ; reg[33:0] dcache_s2_uncached_resp_addr ; 
    wire dcache__GEN_98 = dcache_s1_valid_not_nacked | dcache_s1_flush_valid ; 
    wire[5:0] dcache__GEN_99 = dcache__GEN_98  ?  dcache_s1_req_tag : dcache_s2_req_tag ; 
    wire[4:0] dcache__GEN_100 = dcache__GEN_98  ?  dcache_s1_req_cmd : dcache_s2_req_cmd ; 
    wire[1:0] dcache__GEN_101 = dcache__GEN_98  ?  dcache_s1_req_size : dcache_s2_req_size ; 
    wire dcache__GEN_102 = dcache__GEN_98  ?  dcache_s1_req_signed : dcache_s2_req_signed ; 
    wire[33:0] dcache__GEN_103 ={2'h0, dcache_s1_paddr }; 
    wire[33:0] dcache__GEN_104 = dcache__GEN_98  ?  dcache__GEN_103 : dcache_s2_req_addr ; 
    wire dcache__GEN_105 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_miss : dcache_tlb_io_resp_miss ; 
    wire[31:0] dcache__GEN_106 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_paddr : dcache_tlb_io_resp_paddr ; 
    wire[33:0] dcache__GEN_107 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_gpa : dcache_tlb_io_resp_gpa ; 
    wire dcache__GEN_108 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_gpa_is_pte : dcache_tlb_io_resp_gpa_is_pte ; 
    wire dcache__GEN_109 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_pf_ld : dcache_tlb_io_resp_pf_ld ; 
    wire dcache__GEN_110 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_pf_st : dcache_tlb_io_resp_pf_st ; 
    wire dcache__GEN_111 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_pf_inst : dcache_tlb_io_resp_pf_inst ; 
    wire dcache__GEN_112 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_gf_ld : dcache_tlb_io_resp_gf_ld ; 
    wire dcache__GEN_113 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_gf_st : dcache_tlb_io_resp_gf_st ; 
    wire dcache__GEN_114 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_gf_inst : dcache_tlb_io_resp_gf_inst ; 
    wire dcache__GEN_115 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ae_ld : dcache_tlb_io_resp_ae_ld ; 
    wire dcache__GEN_116 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ae_st : dcache_tlb_io_resp_ae_st ; 
    wire dcache__GEN_117 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ae_inst : dcache_tlb_io_resp_ae_inst ; 
    wire dcache__GEN_118 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ma_ld : dcache_tlb_io_resp_ma_ld ; 
    wire dcache__GEN_119 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ma_st : dcache_tlb_io_resp_ma_st ; 
    wire dcache__GEN_120 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_ma_inst : dcache_tlb_io_resp_ma_inst ; 
    wire dcache__GEN_121 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_cacheable : dcache_tlb_io_resp_cacheable ; 
    wire dcache__GEN_122 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_must_alloc : dcache_tlb_io_resp_must_alloc ; 
    wire dcache__GEN_123 = dcache_s1_tlb_req_valid  ?  dcache_pma_checker_io_resp_prefetchable : dcache_tlb_io_resp_prefetchable ; 
    wire dcache__GEN_124 = dcache_s1_valid_not_nacked | dcache_s1_flush_valid ; reg[33:0] dcache_s2_vaddr_r ; 
    wire[33:0] dcache_s2_vaddr ={ dcache_s2_vaddr_r [33:12], dcache_s2_req_addr [11:0]}; 
    wire dcache_s2_read = dcache_s2_req_cmd ==5'h0| dcache_s2_req_cmd ==5'h10| dcache_s2_req_cmd ==5'h6| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF; 
    wire dcache_s2_write = dcache_s2_req_cmd ==5'h1| dcache_s2_req_cmd ==5'h11| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF; 
    wire dcache_s2_readwrite = dcache_s2_read | dcache_s2_write ; 
    reg dcache_s2_flush_valid_pre_tag_ecc ; 
    wire dcache_s1_meta_clk_en = dcache_s1_valid_not_nacked | dcache_s1_flush_valid | dcache_s1_probe ; 
    reg dcache_s2_meta_correctable_errors ; 
    reg dcache_s2_meta_uncorrectable_errors ; 
    wire dcache_s2_meta_error_uncorrectable =| dcache_s2_meta_uncorrectable_errors ; reg[21:0] dcache_s2_meta_corrected_r ; 
    wire[21:0] dcache__s2_meta_corrected_WIRE = dcache_s2_meta_corrected_r ; 
    wire[19:0] dcache_metaArb_io_in_1_bits_data_new_meta_tag = dcache_s2_meta_corrected_0_tag ; 
  assign  dcache_s2_meta_corrected_0_tag = dcache__s2_meta_corrected_WIRE [19:0]; 
    wire[1:0] dcache_s2_meta_corrected_0_coh_state = dcache__s2_meta_corrected_WIRE [21:20]; 
    wire dcache_s2_meta_error =|( dcache_s2_meta_uncorrectable_errors | dcache_s2_meta_correctable_errors ); 
    wire dcache_s2_flush_valid = dcache_s2_flush_valid_pre_tag_ecc & dcache_s2_meta_error ==1'h0; 
    wire dcache__io_cpu_replay_next_output ; 
    wire dcache_s2_data_en = dcache_s1_valid | dcache_inWriteback | dcache__io_cpu_replay_next_output ; 
    wire dcache_s2_data_word_en = dcache_inWriteback  ? 1'h1: dcache_s1_did_read  ?  dcache_s1_read_mask :1'h0; 
    wire dcache_s2_data_s1_word_en = dcache__io_cpu_replay_next_output ==1'h0 ?  dcache_s2_data_word_en :1'h1; 
    wire[1:0] dcache_s1_data_way ; 
    wire[1:0] dcache__GEN_125 = dcache_s2_data_s1_word_en  ?  dcache_s1_data_way :2'h0; 
    wire[63:0] dcache__s2_data_WIRE =( dcache__GEN_125 [0] ?  dcache_s2_data_s1_way_words_0_0 :64'h0)|( dcache__GEN_125 [1] ?  dcache_s2_data_s1_way_words_1_0 :64'h0); reg[63:0] dcache_s2_data ; 
    reg dcache_s2_probe_way ; reg[1:0] dcache_s2_probe_state_state ; 
    reg dcache_s2_hit_way ; 
    wire dcache__GEN_126 = dcache_s1_valid_not_nacked | dcache_s1_flush_valid ; reg[1:0] dcache_s2_hit_state_state ; 
    reg dcache_s2_waw_hazard ; 
    wire dcache_s2_hit_valid = dcache_s2_hit_state_state >2'h0; 
    wire[1:0] dcache_c ={ dcache_s2_req_cmd ==5'h1| dcache_s2_req_cmd ==5'h11| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF, dcache_s2_req_cmd ==5'h1| dcache_s2_req_cmd ==5'h11| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF| dcache_s2_req_cmd ==5'h3| dcache_s2_req_cmd ==5'h6}; 
    wire[3:0] dcache__GEN_127 ={ dcache_c , dcache_s2_hit_state_state }; 
    wire dcache__GEN_128 =4'hE== dcache__GEN_127 ; 
    wire dcache__GEN_129 =4'hF== dcache__GEN_127 ; 
    wire dcache__GEN_130 =4'h6== dcache__GEN_127 ; 
    wire dcache__GEN_131 =4'h7== dcache__GEN_127 ; 
    wire dcache__GEN_132 =4'h1== dcache__GEN_127 ; 
    wire dcache__GEN_133 =4'h2== dcache__GEN_127 ; 
    wire dcache__GEN_134 =4'h3== dcache__GEN_127 ; 
    wire dcache_s2_hit = dcache__GEN_134  ? 1'h1: dcache__GEN_133  ? 1'h1: dcache__GEN_132  ? 1'h1: dcache__GEN_131  ? 1'h1: dcache__GEN_130  ? 1'h1: dcache__GEN_129  ? 1'h1: dcache__GEN_128 ; 
    wire[1:0] dcache_s2_grow_param = dcache__GEN_134  ? 2'h3: dcache__GEN_133  ? 2'h2: dcache__GEN_132  ? 2'h1: dcache__GEN_131  ? 2'h3: dcache__GEN_130  ? 2'h2: dcache__GEN_129  ? 2'h3: dcache__GEN_128  ? 2'h3:4'h0== dcache__GEN_127  ? 2'h0:4'h5== dcache__GEN_127  ? 2'h2:4'h4== dcache__GEN_127  ? 2'h1:4'hD== dcache__GEN_127  ? 2'h2:4'hC== dcache__GEN_127  ? 2'h1:2'h0; 
    wire[1:0] dcache_s2_new_hit_state_state = dcache_s2_grow_param ; 
    wire[1:0] dcache_metaArb_io_in_2_bits_data_meta_coh_state = dcache_s2_new_hit_state_state ; 
    wire[15:0] dcache_s2_data_corrected_lo_lo ={ dcache_s2_data [15:8], dcache_s2_data [7:0]}; 
    wire[15:0] dcache_s2_data_corrected_lo_hi ={ dcache_s2_data [31:24], dcache_s2_data [23:16]}; 
    wire[31:0] dcache_s2_data_corrected_lo ={ dcache_s2_data_corrected_lo_hi , dcache_s2_data_corrected_lo_lo }; 
    wire[15:0] dcache_s2_data_corrected_hi_lo ={ dcache_s2_data [47:40], dcache_s2_data [39:32]}; 
    wire[15:0] dcache_s2_data_corrected_hi_hi ={ dcache_s2_data [63:56], dcache_s2_data [55:48]}; 
    wire[31:0] dcache_s2_data_corrected_hi ={ dcache_s2_data_corrected_hi_hi , dcache_s2_data_corrected_hi_lo }; 
  assign  dcache_s2_data_corrected ={ dcache_s2_data_corrected_hi , dcache_s2_data_corrected_lo }; 
    wire[63:0] dcache_nodeOut_c_bits_data = dcache_s2_data_corrected ; 
    wire[63:0] dcache_s2_data_word_corrected = dcache_s2_data_corrected ; 
    wire[15:0] dcache_s2_data_uncorrected_lo_lo ={ dcache_s2_data [15:8], dcache_s2_data [7:0]}; 
    wire[15:0] dcache_s2_data_uncorrected_lo_hi ={ dcache_s2_data [31:24], dcache_s2_data [23:16]}; 
    wire[31:0] dcache_s2_data_uncorrected_lo ={ dcache_s2_data_uncorrected_lo_hi , dcache_s2_data_uncorrected_lo_lo }; 
    wire[15:0] dcache_s2_data_uncorrected_hi_lo ={ dcache_s2_data [47:40], dcache_s2_data [39:32]}; 
    wire[15:0] dcache_s2_data_uncorrected_hi_hi ={ dcache_s2_data [63:56], dcache_s2_data [55:48]}; 
    wire[31:0] dcache_s2_data_uncorrected_hi ={ dcache_s2_data_uncorrected_hi_hi , dcache_s2_data_uncorrected_hi_lo }; 
    wire[63:0] dcache_s2_data_uncorrected ={ dcache_s2_data_uncorrected_hi , dcache_s2_data_uncorrected_lo }; 
    wire[63:0] dcache_s2_data_word = dcache_s2_data_uncorrected ; 
    wire dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw = dcache_s2_valid_masked & dcache_s2_meta_error ==1'h0& dcache_s2_hit ; 
    wire dcache_s2_valid_hit_pre_data_ecc_and_waw = dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & dcache_s2_readwrite ; 
    wire dcache_s2_valid_flush_line = dcache_s2_valid_hit_maybe_flush_pre_data_ecc_and_waw & dcache_s2_cmd_flush_line ; 
    wire dcache_s2_valid_hit_pre_data_ecc = dcache_s2_valid_hit_pre_data_ecc_and_waw &( dcache_s2_waw_hazard ==1'h0| dcache_s2_store_merge ); 
    wire dcache_s2_valid_data_error = dcache_s2_valid_hit_pre_data_ecc_and_waw & dcache_s2_data_error ; 
    wire dcache_s2_valid_hit = dcache_s2_valid_hit_pre_data_ecc & dcache_s2_data_error ==1'h0; 
    wire dcache_s2_valid_miss = dcache_s2_valid_masked & dcache_s2_readwrite & dcache_s2_meta_error ==1'h0& dcache_s2_hit ==1'h0; 
    wire dcache_s2_uncached = dcache_s2_pma_cacheable ==1'h0| dcache_s2_req_no_alloc & dcache_s2_pma_must_alloc ==1'h0& dcache_s2_hit_valid ==1'h0; 
    wire dcache_s2_valid_cached_miss = dcache_s2_valid_miss & dcache_s2_uncached ==1'h0&(| dcache_uncachedInFlight_0 )==1'h0; 
    wire dcache_s2_want_victimize =( dcache_s2_valid_cached_miss | dcache_s2_valid_flush_line | dcache_s2_valid_data_error | dcache_s2_flush_valid )&1'h1; 
    wire dcache_s2_cannot_victimize = dcache_s2_flush_valid ==1'h0& dcache_io_cpu_s2_kill ; 
    wire dcache_s2_victimize = dcache_s2_want_victimize & dcache_s2_cannot_victimize ==1'h0; 
    wire dcache_s2_valid_uncached_pending = dcache_s2_valid_miss & dcache_s2_uncached &(& dcache_uncachedInFlight_0 )==1'h0; 
    wire dcache__GEN_135 = dcache_s1_valid_not_nacked | dcache_s1_flush_valid ; 
    reg dcache_s2_victim_way_r ; 
    wire[1:0] dcache_s2_victim_way =2'h1<< dcache_s2_victim_way_r ; 
    wire[1:0] dcache_s2_victim_or_hit_way = dcache_s2_hit_valid  ? {1'h0, dcache_s2_hit_way }: dcache_s2_victim_way ; 
    wire[19:0] dcache_s2_victim_tag = dcache_s2_valid_data_error | dcache_s2_valid_flush_line  ?  dcache_s2_req_addr [31:12]: dcache_s2_meta_corrected_0_tag ; 
    wire[1:0] dcache_s2_victim_state_state = dcache_s2_hit_valid  ?  dcache_s2_hit_state_state : dcache_s2_meta_corrected_0_coh_state ; 
    wire[3:0] dcache__GEN_136 ={ dcache_probe_bits_param , dcache_s2_probe_state_state }; 
    wire dcache__GEN_137 =4'h8== dcache__GEN_136 ; 
    wire dcache__GEN_138 =4'h9== dcache__GEN_136 ; 
    wire dcache__GEN_139 =4'hA== dcache__GEN_136 ; 
    wire dcache__GEN_140 =4'hB== dcache__GEN_136 ; 
    wire dcache__GEN_141 =4'h4== dcache__GEN_136 ; 
    wire dcache__GEN_142 =4'h5== dcache__GEN_136 ; 
    wire dcache__GEN_143 =4'h6== dcache__GEN_136 ; 
    wire dcache__GEN_144 =4'h7== dcache__GEN_136 ; 
    wire dcache__GEN_145 =4'h0== dcache__GEN_136 ; 
    wire dcache__GEN_146 =4'h1== dcache__GEN_136 ; 
    wire dcache__GEN_147 =4'h2== dcache__GEN_136 ; 
    wire dcache__GEN_148 =4'h3== dcache__GEN_136 ; 
    wire dcache_s2_prb_ack_data = dcache__GEN_148  ? 1'h1: dcache__GEN_147  ? 1'h0: dcache__GEN_146  ? 1'h0: dcache__GEN_145  ? 1'h0: dcache__GEN_144  ? 1'h1: dcache__GEN_143  ? 1'h0: dcache__GEN_142  ? 1'h0: dcache__GEN_141  ? 1'h0: dcache__GEN_140 ; 
    wire[2:0] dcache_s2_report_param = dcache__GEN_148  ? 3'h3: dcache__GEN_147  ? 3'h3: dcache__GEN_146  ? 3'h4: dcache__GEN_145  ? 3'h5: dcache__GEN_144  ? 3'h0: dcache__GEN_143  ? 3'h0: dcache__GEN_142  ? 3'h4: dcache__GEN_141  ? 3'h5: dcache__GEN_140  ? 3'h1: dcache__GEN_139  ? 3'h1: dcache__GEN_138  ? 3'h2: dcache__GEN_137  ? 3'h5:3'h0; 
    wire[2:0] dcache_cleanReleaseMessage_param = dcache_s2_report_param ; 
    wire[2:0] dcache_dirtyReleaseMessage_param = dcache_s2_report_param ; 
    wire[1:0] dcache_probeNewCoh_state = dcache__GEN_148  ? 2'h2: dcache__GEN_147  ? 2'h2: dcache__GEN_146  ? 2'h1: dcache__GEN_145  ? 2'h0: dcache__GEN_144  ? 2'h1: dcache__GEN_143  ? 2'h1: dcache__GEN_142  ? 2'h1: dcache__GEN_141  ? 2'h0: dcache__GEN_140  ? 2'h0: dcache__GEN_139  ? 2'h0: dcache__GEN_138  ? 2'h0: dcache__GEN_137  ? 2'h0:2'h0; 
    wire[3:0] dcache__GEN_149 ={2'h2, dcache_s2_victim_state_state }; 
    wire dcache__GEN_150 =4'h8== dcache__GEN_149 ; 
    wire dcache__GEN_151 =4'h9== dcache__GEN_149 ; 
    wire dcache__GEN_152 =4'hA== dcache__GEN_149 ; 
    wire dcache__GEN_153 =4'hB== dcache__GEN_149 ; 
    wire dcache__GEN_154 =4'h4== dcache__GEN_149 ; 
    wire dcache__GEN_155 =4'h5== dcache__GEN_149 ; 
    wire dcache__GEN_156 =4'h6== dcache__GEN_149 ; 
    wire dcache__GEN_157 =4'h7== dcache__GEN_149 ; 
    wire dcache__GEN_158 =4'h0== dcache__GEN_149 ; 
    wire dcache__GEN_159 =4'h1== dcache__GEN_149 ; 
    wire dcache__GEN_160 =4'h2== dcache__GEN_149 ; 
    wire dcache__GEN_161 =4'h3== dcache__GEN_149 ; 
    wire dcache_s2_victim_dirty = dcache__GEN_161  ? 1'h1: dcache__GEN_160  ? 1'h0: dcache__GEN_159  ? 1'h0: dcache__GEN_158  ? 1'h0: dcache__GEN_157  ? 1'h1: dcache__GEN_156  ? 1'h0: dcache__GEN_155  ? 1'h0: dcache__GEN_154  ? 1'h0: dcache__GEN_153 ; 
    wire[2:0] dcache_s2_shrink_param = dcache__GEN_161  ? 3'h3: dcache__GEN_160  ? 3'h3: dcache__GEN_159  ? 3'h4: dcache__GEN_158  ? 3'h5: dcache__GEN_157  ? 3'h0: dcache__GEN_156  ? 3'h0: dcache__GEN_155  ? 3'h4: dcache__GEN_154  ? 3'h5: dcache__GEN_153  ? 3'h1: dcache__GEN_152  ? 3'h1: dcache__GEN_151  ? 3'h2: dcache__GEN_150  ? 3'h5:3'h0; 
    wire[2:0] dcache_nodeOut_c_bits_c_param = dcache_s2_shrink_param ; 
    wire[2:0] dcache_nodeOut_c_bits_c_1_param = dcache_s2_shrink_param ; 
    wire[1:0] dcache_voluntaryNewCoh_state = dcache__GEN_161  ? 2'h2: dcache__GEN_160  ? 2'h2: dcache__GEN_159  ? 2'h1: dcache__GEN_158  ? 2'h0: dcache__GEN_157  ? 2'h1: dcache__GEN_156  ? 2'h1: dcache__GEN_155  ? 2'h1: dcache__GEN_154  ? 2'h0: dcache__GEN_153  ? 2'h0: dcache__GEN_152  ? 2'h0: dcache__GEN_151  ? 2'h0: dcache__GEN_150  ? 2'h0:2'h0; 
    wire dcache_s2_update_meta = dcache_s2_hit_state_state == dcache_s2_new_hit_state_state ==1'h0; 
    wire dcache_s2_dont_nack_uncached = dcache_s2_valid_uncached_pending & dcache_tl_out_a_ready ; 
    wire dcache_s2_dont_nack_misc = dcache_s2_valid_masked & dcache_s2_meta_error ==1'h0&( dcache_s2_req_cmd ==5'h17|1'h0); 
    wire dcache__io_cpu_s2_nack_output = dcache_s2_valid_no_xcpt & dcache_s2_dont_nack_uncached ==1'h0& dcache_s2_dont_nack_misc ==1'h0& dcache_s2_valid_hit ==1'h0; 
  assign  dcache_metaArb_io_in_1_valid = dcache_s2_meta_error &( dcache_s2_valid_masked | dcache_s2_flush_valid_pre_tag_ecc | dcache_s2_probe ); 
  assign  dcache_metaArb_io_in_1_bits_way_en = dcache_s2_meta_uncorrectable_errors |( dcache_s2_meta_error_uncorrectable  ? 1'h0: dcache_s2_meta_correctable_errors ); 
  assign  dcache_metaArb_io_in_1_bits_idx = dcache_s2_probe  ?  dcache_probe_bits_address [11:6]: dcache_s2_vaddr [11:6]; 
  assign  dcache_metaArb_io_in_1_bits_addr ={ dcache_io_cpu_req_bits_addr [33:12],{ dcache_metaArb_io_in_1_bits_idx ,6'h0}}; 
    wire[1:0] dcache_metaArb_io_in_1_bits_data_new_meta_coh_state = dcache_s2_meta_error_uncorrectable  ?  dcache_metaArb_io_in_1_bits_data_new_meta_coh_meta_state : dcache_s2_meta_corrected_0_coh_state ; 
  assign  dcache_metaArb_io_in_1_bits_data ={ dcache_metaArb_io_in_1_bits_data_new_meta_coh_state , dcache_metaArb_io_in_1_bits_data_new_meta_tag }; 
  assign  dcache_metaArb_io_in_2_valid = dcache_s2_valid_hit_pre_data_ecc_and_waw & dcache_s2_update_meta ; 
  assign  dcache_metaArb_io_in_2_bits_write = dcache_io_cpu_s2_kill ==1'h0; 
  assign  dcache_metaArb_io_in_2_bits_way_en = dcache_s2_victim_or_hit_way [0]; 
  assign  dcache_metaArb_io_in_2_bits_idx = dcache_s2_vaddr [11:6]; 
  assign  dcache_metaArb_io_in_2_bits_addr ={ dcache_io_cpu_req_bits_addr [33:12], dcache_s2_vaddr [11:0]}; 
    wire[21:0] dcache__s2_req_addr_33to12 = dcache_s2_req_addr [33:12]; 
    wire[19:0] dcache_metaArb_io_in_2_bits_data_meta_tag = dcache__s2_req_addr_33to12 [19:0]; 
  assign  dcache_metaArb_io_in_2_bits_data ={ dcache_metaArb_io_in_2_bits_data_meta_coh_state , dcache_metaArb_io_in_2_bits_data_meta_tag }; 
    wire dcache_s2_lr = dcache_s2_req_cmd ==5'h6&1'h1; 
    wire dcache_s2_sc = dcache_s2_req_cmd ==5'h7&1'h1; reg[6:0] dcache_lrscCount ; 
    wire dcache_lrscValid = dcache_lrscCount >7'h3; 
    wire dcache_lrscBackingOff = dcache_lrscCount >7'h0& dcache_lrscValid ==1'h0; reg[27:0] dcache_lrscAddr ; 
    wire dcache_lrscAddrMatch = dcache_lrscAddr == dcache_s2_req_addr [33:6]; 
    wire dcache_s2_sc_fail = dcache_s2_sc &( dcache_lrscValid & dcache_lrscAddrMatch )==1'h0; 
    wire dcache__GEN_162 =( dcache_s2_valid_hit & dcache_s2_lr & dcache_cached_grant_wait ==1'h0| dcache_s2_valid_cached_miss )& dcache_io_cpu_s2_kill ==1'h0; 
    wire[6:0] dcache__GEN_163 = dcache_s2_hit  ? 7'h4F:7'h0; 
    wire dcache__GEN_164 = dcache_lrscCount >7'h0; 
    wire[7:0] dcache__GEN_165 ={1'h0, dcache_lrscCount }-8'h1; 
    wire dcache__GEN_166 = dcache_s2_valid_not_killed & dcache_lrscValid ; 
    wire dcache_any_pstore_valid ; 
    reg dcache_s2_correct_REG ; 
    wire dcache_s2_valid_correct = dcache_s2_valid_hit_pre_data_ecc_and_waw & dcache_s2_correct & dcache_io_cpu_s2_kill ==1'h0; 
    wire dcache__GEN_167 = dcache_s1_valid_not_nacked & dcache_s1_write ; reg[4:0] dcache_pstore1_cmd ; 
    wire dcache__GEN_168 = dcache_s1_valid_not_nacked & dcache_s1_write ; reg[33:0] dcache_pstore1_addr ; 
    wire dcache__GEN_169 = dcache_s1_valid_not_nacked & dcache_s1_write ; reg[63:0] dcache_pstore1_data ; 
    wire[63:0] dcache_put_data = dcache_pstore1_data ; 
    wire[63:0] dcache_putpartial_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_1_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_2_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_3_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_4_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_5_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_6_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_7_data = dcache_pstore1_data ; 
    wire[63:0] dcache_atomics_a_8_data = dcache_pstore1_data ; 
    wire dcache__GEN_170 = dcache_s1_valid_not_nacked & dcache_s1_write ; 
    reg dcache_pstore1_way ; 
    wire dcache__GEN_171 = dcache_s1_valid_not_nacked & dcache_s1_write ; reg[7:0] dcache_pstore1_mask ; 
    wire dcache__GEN_172 = dcache_s1_req_cmd ==5'h0| dcache_s1_req_cmd ==5'h10| dcache_s1_req_cmd ==5'h6| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF|( dcache_s1_req_cmd ==5'h1| dcache_s1_req_cmd ==5'h11| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF)&( dcache_s1_req_cmd ==5'h11| dcache_s1_req_size <2'h0); 
    wire dcache__GEN_173 = dcache_s1_valid_not_nacked & dcache_s1_write ; 
    reg dcache_pstore1_rmw_r ; 
    wire dcache_pstore1_rmw = dcache_pstore1_rmw_r &1'h1; 
    wire dcache_pstore1_merge_likely = dcache_s2_valid_not_nacked_in_s1 & dcache_s2_write & dcache_s2_store_merge ; 
    wire dcache_pstore1_merge = dcache_s2_valid_hit & dcache_s2_write & dcache_s2_sc_fail ==1'h0& dcache_io_cpu_s2_kill ==1'h0& dcache_s2_store_merge ; 
    reg dcache_pstore2_valid ; 
    wire dcache_pstore_drain_opportunistic_res =( dcache_io_cpu_req_bits_cmd ==5'h1| dcache_io_cpu_req_bits_cmd ==5'h3)==1'h0| dcache_io_cpu_req_bits_size <2'h0; 
    wire dcache__GEN_174 =(( dcache_io_cpu_req_bits_cmd ==5'h0| dcache_io_cpu_req_bits_cmd ==5'h10| dcache_io_cpu_req_bits_cmd ==5'h6| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF|( dcache_io_cpu_req_bits_cmd ==5'h1| dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_cmd ==5'h7| dcache_io_cpu_req_bits_cmd ==5'h4| dcache_io_cpu_req_bits_cmd ==5'h9| dcache_io_cpu_req_bits_cmd ==5'hA| dcache_io_cpu_req_bits_cmd ==5'hB| dcache_io_cpu_req_bits_cmd ==5'h8| dcache_io_cpu_req_bits_cmd ==5'hC| dcache_io_cpu_req_bits_cmd ==5'hD| dcache_io_cpu_req_bits_cmd ==5'hE| dcache_io_cpu_req_bits_cmd ==5'hF)&( dcache_io_cpu_req_bits_cmd ==5'h11| dcache_io_cpu_req_bits_size <2'h0))==1'h0| dcache_pstore_drain_opportunistic_res )==1'h0; 
    wire dcache_pstore_drain_opportunistic =( dcache_io_cpu_req_valid & dcache_pstore_drain_opportunistic_res )==1'h0&( dcache_s1_valid & dcache_s1_waw_hazard )==1'h0; 
    reg dcache_pstore_drain_on_miss_REG ; 
    wire dcache_pstore_drain_on_miss = dcache_releaseInFlight | dcache_pstore_drain_on_miss_REG ; 
    reg dcache_pstore1_held ; 
    wire dcache_pstore1_valid_likely = dcache_s2_valid & dcache_s2_write | dcache_pstore1_held ; 
    wire dcache_pstore1_valid = dcache_s2_valid_hit & dcache_s2_write & dcache_s2_sc_fail ==1'h0& dcache_io_cpu_s2_kill ==1'h0| dcache_pstore1_held ; 
  assign  dcache_any_pstore_valid = dcache_pstore1_held | dcache_pstore2_valid ; 
    wire dcache_pstore_drain_structural = dcache_pstore1_valid_likely & dcache_pstore2_valid &( dcache_s1_valid & dcache_s1_write | dcache_pstore1_rmw ); 
    wire dcache__GEN_175 =( dcache_pstore1_rmw |( dcache_s2_valid_hit_pre_data_ecc & dcache_s2_write & dcache_io_cpu_s2_kill ==1'h0| dcache_pstore1_held )== dcache_pstore1_valid )==1'h0; 
    wire dcache_pstore_drain_s2_kill = dcache_io_cpu_s2_kill &1'h1; 
  assign  dcache_pstore_drain = dcache_pstore1_merge_likely ==1'h0&( dcache_pstore_drain_structural &1'h1|(( dcache_s2_valid_hit_pre_data_ecc & dcache_s2_write & dcache_pstore_drain_s2_kill ==1'h0| dcache_pstore1_held )& dcache_pstore1_rmw ==1'h0| dcache_pstore2_valid )&( dcache_pstore_drain_opportunistic | dcache_pstore_drain_on_miss )); 
  assign  dcache_dataArb_io_in_0_bits_write = dcache_pstore_drain ; 
    wire dcache_advance_pstore1 =( dcache_pstore1_valid | dcache_s2_valid_correct )& dcache_pstore2_valid == dcache_pstore_drain ; 
    wire[33:0] dcache__GEN_176 = dcache_s2_correct  ?  dcache_s2_vaddr : dcache_pstore1_addr ; reg[33:0] dcache_pstore2_addr ; 
    wire dcache__GEN_177 = dcache_s2_correct  ?  dcache_s2_hit_way : dcache_pstore1_way ; 
    reg dcache_pstore2_way ; 
    wire[63:0] dcache_pstore1_storegen_data ; 
    wire dcache__GEN_178 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [0]; reg[7:0] dcache_pstore2_storegen_data_r ; 
    wire dcache__GEN_179 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [1]; reg[7:0] dcache_pstore2_storegen_data_r_1 ; 
    wire dcache__GEN_180 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [2]; reg[7:0] dcache_pstore2_storegen_data_r_2 ; 
    wire dcache__GEN_181 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [3]; reg[7:0] dcache_pstore2_storegen_data_r_3 ; 
    wire dcache__GEN_182 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [4]; reg[7:0] dcache_pstore2_storegen_data_r_4 ; 
    wire dcache__GEN_183 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [5]; reg[7:0] dcache_pstore2_storegen_data_r_5 ; 
    wire dcache__GEN_184 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [6]; reg[7:0] dcache_pstore2_storegen_data_r_6 ; 
    wire dcache__GEN_185 = dcache_advance_pstore1 | dcache_pstore1_merge & dcache_pstore1_mask [7]; reg[7:0] dcache_pstore2_storegen_data_r_7 ; 
    wire[15:0] dcache_pstore2_storegen_data_lo_lo ={ dcache_pstore2_storegen_data_r_1 , dcache_pstore2_storegen_data_r }; 
    wire[15:0] dcache_pstore2_storegen_data_lo_hi ={ dcache_pstore2_storegen_data_r_3 , dcache_pstore2_storegen_data_r_2 }; 
    wire[31:0] dcache_pstore2_storegen_data_lo ={ dcache_pstore2_storegen_data_lo_hi , dcache_pstore2_storegen_data_lo_lo }; 
    wire[15:0] dcache_pstore2_storegen_data_hi_lo ={ dcache_pstore2_storegen_data_r_5 , dcache_pstore2_storegen_data_r_4 }; 
    wire[15:0] dcache_pstore2_storegen_data_hi_hi ={ dcache_pstore2_storegen_data_r_7 , dcache_pstore2_storegen_data_r_6 }; 
    wire[31:0] dcache_pstore2_storegen_data_hi ={ dcache_pstore2_storegen_data_hi_hi , dcache_pstore2_storegen_data_hi_lo }; 
    wire[63:0] dcache_pstore2_storegen_data ={ dcache_pstore2_storegen_data_hi , dcache_pstore2_storegen_data_lo }; reg[7:0] dcache_pstore2_storegen_mask ; 
    wire dcache__GEN_186 = dcache_advance_pstore1 | dcache_pstore1_merge ; 
    wire[7:0] dcache_pstore2_storegen_mask_mergedMask = dcache_pstore1_mask |( dcache_pstore1_merge  ?  dcache_pstore2_storegen_mask :8'h0); 
    wire[7:0] dcache__GEN_187 =~( dcache_s2_correct  ? 8'h0:~ dcache_pstore2_storegen_mask_mergedMask ); 
  assign  dcache_dataArb_io_in_0_valid = dcache_pstore1_merge_likely ==1'h0&( dcache_pstore_drain_structural &1'h1|(( dcache_s2_valid_hit_pre_data_ecc & dcache_s2_write & dcache_dataArb_io_in_0_valid_s2_kill ==1'h0| dcache_pstore1_held )& dcache_pstore1_rmw ==1'h0| dcache_pstore2_valid )&( dcache_pstore_drain_opportunistic | dcache_pstore_drain_on_miss )); 
    wire[33:0] dcache__GEN_188 = dcache_pstore2_valid  ?  dcache_pstore2_addr : dcache_pstore1_addr ; 
  assign  dcache_dataArb_io_in_0_bits_addr = dcache__GEN_188 [11:0]; 
  assign  dcache_dataArb_io_in_0_bits_way_en = dcache_pstore2_valid  ?  dcache_pstore2_way : dcache_pstore1_way ; 
    wire[63:0] dcache__GEN_189 = dcache_pstore2_valid  ?  dcache_pstore2_storegen_data : dcache_pstore1_data ; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_lo_lo ={ dcache__GEN_189 [15:8], dcache__GEN_189 [7:0]}; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_lo_hi ={ dcache__GEN_189 [31:24], dcache__GEN_189 [23:16]}; 
    wire[31:0] dcache_dataArb_io_in_0_bits_wdata_lo ={ dcache_dataArb_io_in_0_bits_wdata_lo_hi , dcache_dataArb_io_in_0_bits_wdata_lo_lo }; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_hi_lo ={ dcache__GEN_189 [47:40], dcache__GEN_189 [39:32]}; 
    wire[15:0] dcache_dataArb_io_in_0_bits_wdata_hi_hi ={ dcache__GEN_189 [63:56], dcache__GEN_189 [55:48]}; 
    wire[31:0] dcache_dataArb_io_in_0_bits_wdata_hi ={ dcache_dataArb_io_in_0_bits_wdata_hi_hi , dcache_dataArb_io_in_0_bits_wdata_hi_lo }; 
  assign  dcache_dataArb_io_in_0_bits_wdata ={ dcache_dataArb_io_in_0_bits_wdata_hi , dcache_dataArb_io_in_0_bits_wdata_lo }; 
    wire dcache_dataArb_io_in_0_bits_wordMask_eccMask = dcache_dataArb_io_in_0_bits_eccMask [0]| dcache_dataArb_io_in_0_bits_eccMask [1]| dcache_dataArb_io_in_0_bits_eccMask [2]| dcache_dataArb_io_in_0_bits_eccMask [3]| dcache_dataArb_io_in_0_bits_eccMask [4]| dcache_dataArb_io_in_0_bits_eccMask [5]| dcache_dataArb_io_in_0_bits_eccMask [6]| dcache_dataArb_io_in_0_bits_eccMask [7]; 
    wire[1:0] dcache_dataArb_io_in_0_bits_wordMask_wordMask =2'h1; 
    wire[1:0] dcache__GEN_190 ={ dcache_dataArb_io_in_0_bits_wordMask_wordMask [1], dcache_dataArb_io_in_0_bits_wordMask_wordMask [0]}&{1'h0, dcache_dataArb_io_in_0_bits_wordMask_eccMask }; 
  assign  dcache_dataArb_io_in_0_bits_wordMask = dcache__GEN_190 [0]; 
    wire[7:0] dcache__GEN_191 = dcache_pstore2_valid  ?  dcache_pstore2_storegen_mask : dcache_pstore1_mask ; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_lo_lo ={|( dcache__GEN_191 [1]),|( dcache__GEN_191 [0])}; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_lo_hi ={|( dcache__GEN_191 [3]),|( dcache__GEN_191 [2])}; 
    wire[3:0] dcache_dataArb_io_in_0_bits_eccMask_lo ={ dcache_dataArb_io_in_0_bits_eccMask_lo_hi , dcache_dataArb_io_in_0_bits_eccMask_lo_lo }; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_hi_lo ={|( dcache__GEN_191 [5]),|( dcache__GEN_191 [4])}; 
    wire[1:0] dcache_dataArb_io_in_0_bits_eccMask_hi_hi ={|( dcache__GEN_191 [7]),|( dcache__GEN_191 [6])}; 
    wire[3:0] dcache_dataArb_io_in_0_bits_eccMask_hi ={ dcache_dataArb_io_in_0_bits_eccMask_hi_hi , dcache_dataArb_io_in_0_bits_eccMask_hi_lo }; 
  assign  dcache_dataArb_io_in_0_bits_eccMask ={ dcache_dataArb_io_in_0_bits_eccMask_hi , dcache_dataArb_io_in_0_bits_eccMask_lo }; 
    wire[1:0] dcache_s1_hazard_lo_lo ={|( dcache_pstore1_mask [1]),|( dcache_pstore1_mask [0])}; 
    wire[1:0] dcache_s1_hazard_lo_hi ={|( dcache_pstore1_mask [3]),|( dcache_pstore1_mask [2])}; 
    wire[3:0] dcache_s1_hazard_lo ={ dcache_s1_hazard_lo_hi , dcache_s1_hazard_lo_lo }; 
    wire[1:0] dcache_s1_hazard_hi_lo ={|( dcache_pstore1_mask [5]),|( dcache_pstore1_mask [4])}; 
    wire[1:0] dcache_s1_hazard_hi_hi ={|( dcache_pstore1_mask [7]),|( dcache_pstore1_mask [6])}; 
    wire[3:0] dcache_s1_hazard_hi ={ dcache_s1_hazard_hi_hi , dcache_s1_hazard_hi_lo }; 
    wire[7:0] dcache__GEN_192 ={ dcache_s1_hazard_hi , dcache_s1_hazard_lo }; 
    wire[1:0] dcache_s1_hazard_lo_lo_1 ={ dcache__GEN_192 [1], dcache__GEN_192 [0]}; 
    wire[1:0] dcache_s1_hazard_lo_hi_1 ={ dcache__GEN_192 [3], dcache__GEN_192 [2]}; 
    wire[3:0] dcache_s1_hazard_lo_1 ={ dcache_s1_hazard_lo_hi_1 , dcache_s1_hazard_lo_lo_1 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_1 ={ dcache__GEN_192 [5], dcache__GEN_192 [4]}; 
    wire[1:0] dcache_s1_hazard_hi_hi_1 ={ dcache__GEN_192 [7], dcache__GEN_192 [6]}; 
    wire[3:0] dcache_s1_hazard_hi_1 ={ dcache_s1_hazard_hi_hi_1 , dcache_s1_hazard_hi_lo_1 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_2 ={|( dcache_s1_mask_xwr [1]),|( dcache_s1_mask_xwr [0])}; 
    wire[1:0] dcache_s1_hazard_lo_hi_2 ={|( dcache_s1_mask_xwr [3]),|( dcache_s1_mask_xwr [2])}; 
    wire[3:0] dcache_s1_hazard_lo_2 ={ dcache_s1_hazard_lo_hi_2 , dcache_s1_hazard_lo_lo_2 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_2 ={|( dcache_s1_mask_xwr [5]),|( dcache_s1_mask_xwr [4])}; 
    wire[1:0] dcache_s1_hazard_hi_hi_2 ={|( dcache_s1_mask_xwr [7]),|( dcache_s1_mask_xwr [6])}; 
    wire[3:0] dcache_s1_hazard_hi_2 ={ dcache_s1_hazard_hi_hi_2 , dcache_s1_hazard_hi_lo_2 }; 
    wire[7:0] dcache__GEN_193 ={ dcache_s1_hazard_hi_2 , dcache_s1_hazard_lo_2 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_3 ={ dcache__GEN_193 [1], dcache__GEN_193 [0]}; 
    wire[1:0] dcache_s1_hazard_lo_hi_3 ={ dcache__GEN_193 [3], dcache__GEN_193 [2]}; 
    wire[3:0] dcache_s1_hazard_lo_3 ={ dcache_s1_hazard_lo_hi_3 , dcache_s1_hazard_lo_lo_3 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_3 ={ dcache__GEN_193 [5], dcache__GEN_193 [4]}; 
    wire[1:0] dcache_s1_hazard_hi_hi_3 ={ dcache__GEN_193 [7], dcache__GEN_193 [6]}; 
    wire[3:0] dcache_s1_hazard_hi_3 ={ dcache_s1_hazard_hi_hi_3 , dcache_s1_hazard_hi_lo_3 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_4 ={|( dcache_pstore2_storegen_mask [1]),|( dcache_pstore2_storegen_mask [0])}; 
    wire[1:0] dcache_s1_hazard_lo_hi_4 ={|( dcache_pstore2_storegen_mask [3]),|( dcache_pstore2_storegen_mask [2])}; 
    wire[3:0] dcache_s1_hazard_lo_4 ={ dcache_s1_hazard_lo_hi_4 , dcache_s1_hazard_lo_lo_4 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_4 ={|( dcache_pstore2_storegen_mask [5]),|( dcache_pstore2_storegen_mask [4])}; 
    wire[1:0] dcache_s1_hazard_hi_hi_4 ={|( dcache_pstore2_storegen_mask [7]),|( dcache_pstore2_storegen_mask [6])}; 
    wire[3:0] dcache_s1_hazard_hi_4 ={ dcache_s1_hazard_hi_hi_4 , dcache_s1_hazard_hi_lo_4 }; 
    wire[7:0] dcache__GEN_194 ={ dcache_s1_hazard_hi_4 , dcache_s1_hazard_lo_4 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_5 ={ dcache__GEN_194 [1], dcache__GEN_194 [0]}; 
    wire[1:0] dcache_s1_hazard_lo_hi_5 ={ dcache__GEN_194 [3], dcache__GEN_194 [2]}; 
    wire[3:0] dcache_s1_hazard_lo_5 ={ dcache_s1_hazard_lo_hi_5 , dcache_s1_hazard_lo_lo_5 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_5 ={ dcache__GEN_194 [5], dcache__GEN_194 [4]}; 
    wire[1:0] dcache_s1_hazard_hi_hi_5 ={ dcache__GEN_194 [7], dcache__GEN_194 [6]}; 
    wire[3:0] dcache_s1_hazard_hi_5 ={ dcache_s1_hazard_hi_hi_5 , dcache_s1_hazard_hi_lo_5 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_6 ={|( dcache_s1_mask_xwr [1]),|( dcache_s1_mask_xwr [0])}; 
    wire[1:0] dcache_s1_hazard_lo_hi_6 ={|( dcache_s1_mask_xwr [3]),|( dcache_s1_mask_xwr [2])}; 
    wire[3:0] dcache_s1_hazard_lo_6 ={ dcache_s1_hazard_lo_hi_6 , dcache_s1_hazard_lo_lo_6 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_6 ={|( dcache_s1_mask_xwr [5]),|( dcache_s1_mask_xwr [4])}; 
    wire[1:0] dcache_s1_hazard_hi_hi_6 ={|( dcache_s1_mask_xwr [7]),|( dcache_s1_mask_xwr [6])}; 
    wire[3:0] dcache_s1_hazard_hi_6 ={ dcache_s1_hazard_hi_hi_6 , dcache_s1_hazard_hi_lo_6 }; 
    wire[7:0] dcache__GEN_195 ={ dcache_s1_hazard_hi_6 , dcache_s1_hazard_lo_6 }; 
    wire[1:0] dcache_s1_hazard_lo_lo_7 ={ dcache__GEN_195 [1], dcache__GEN_195 [0]}; 
    wire[1:0] dcache_s1_hazard_lo_hi_7 ={ dcache__GEN_195 [3], dcache__GEN_195 [2]}; 
    wire[3:0] dcache_s1_hazard_lo_7 ={ dcache_s1_hazard_lo_hi_7 , dcache_s1_hazard_lo_lo_7 }; 
    wire[1:0] dcache_s1_hazard_hi_lo_7 ={ dcache__GEN_195 [5], dcache__GEN_195 [4]}; 
    wire[1:0] dcache_s1_hazard_hi_hi_7 ={ dcache__GEN_195 [7], dcache__GEN_195 [6]}; 
    wire[3:0] dcache_s1_hazard_hi_7 ={ dcache_s1_hazard_hi_hi_7 , dcache_s1_hazard_hi_lo_7 }; 
    wire dcache_s1_hazard = dcache_pstore1_valid_likely & dcache_pstore1_addr [11:3]== dcache_s1_vaddr [11:3]&( dcache_s1_write  ? (|({ dcache_s1_hazard_hi_1 , dcache_s1_hazard_lo_1 }&{ dcache_s1_hazard_hi_3 , dcache_s1_hazard_lo_3 })):(|( dcache_pstore1_mask & dcache_s1_mask_xwr )))| dcache_pstore2_valid & dcache_pstore2_addr [11:3]== dcache_s1_vaddr [11:3]&( dcache_s1_write  ? (|({ dcache_s1_hazard_hi_5 , dcache_s1_hazard_lo_5 }&{ dcache_s1_hazard_hi_7 , dcache_s1_hazard_lo_7 })):(|( dcache_pstore2_storegen_mask & dcache_s1_mask_xwr ))); 
    wire dcache_s1_raw_hazard = dcache_s1_read & dcache_s1_hazard ; 
    wire dcache__GEN_196 = dcache_s1_valid & dcache_s1_raw_hazard  ? 1'h1: dcache__io_cpu_s2_nack_output | dcache_s2_valid_hit_pre_data_ecc_and_waw & dcache_s2_update_meta  ? 1'h1: dcache_s1_tlb_req_valid & dcache_s1_valid &( dcache_s1_req_phys & dcache_s1_req_no_xcpt )==1'h0 ? 1'h1: dcache_s1_tlb_req_valid ==1'h0& dcache_s1_valid & dcache_s1_cmd_uses_tlb & dcache_tlb_io_resp_miss ; 
    reg dcache_io_cpu_s2_nack_cause_raw_REG ; 
    wire[1:0] dcache__GEN_197 ={~ dcache_uncachedInFlight_0 ,1'h0}; 
    wire dcache_a_source = dcache__GEN_197 [0] ? 1'h0:1'h1; 
    wire dcache_get_source = dcache_a_source ; 
    wire dcache_put_source = dcache_a_source ; 
    wire dcache_putpartial_source = dcache_a_source ; 
    wire dcache_atomics_a_source = dcache_a_source ; 
    wire dcache_atomics_a_1_source = dcache_a_source ; 
    wire dcache_atomics_a_2_source = dcache_a_source ; 
    wire dcache_atomics_a_3_source = dcache_a_source ; 
    wire dcache_atomics_a_4_source = dcache_a_source ; 
    wire dcache_atomics_a_5_source = dcache_a_source ; 
    wire dcache_atomics_a_6_source = dcache_a_source ; 
    wire dcache_atomics_a_7_source = dcache_a_source ; 
    wire dcache_atomics_a_8_source = dcache_a_source ; 
    wire dcache_a_sel_shiftAmount = dcache_a_source ; 
    wire[33:0] dcache_acquire_address ={ dcache_s2_req_addr [33:6],6'h0}; 
    wire[22:0] dcache_a_mask ={15'h0, dcache_pstore1_mask }; 
    wire dcache_get_legal =(2'h0<= dcache_s2_req_size &{2'h0, dcache_s2_req_size }<=4'hC|1'h0)&({1'h0, dcache_s2_req_addr ^34'h2000}&35'hCA012000)==35'h0|1'h0|(2'h0<= dcache_s2_req_size &{1'h0, dcache_s2_req_size }<=3'h6|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hCA012000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h10000}&35'hCA010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h80000000}&35'hC0000000)==35'h0); 
    wire[2:0] dcache_get_param =3'h0; 
    wire[3:0] dcache_get_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_get_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_198 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_get_a_mask_sizeOH_shiftAmount = dcache__GEN_198 [1:0]; 
    wire[3:0] dcache__GEN_199 =4'h1<< dcache_get_a_mask_sizeOH_shiftAmount ; 
    wire[2:0] dcache_get_a_mask_sizeOH = dcache__GEN_199 [2:0]|3'h1; 
    wire dcache__GEN_200 = dcache_s2_req_size >=2'h3; 
    wire dcache_get_a_mask_size = dcache_get_a_mask_sizeOH [2]; 
    wire dcache_get_a_mask_bit = dcache_s2_req_addr [2]; 
    wire dcache_get_a_mask_nbit = dcache_get_a_mask_bit ==1'h0; 
    wire dcache_get_a_mask_eq = dcache_get_a_mask_nbit &1'h1; 
    wire dcache_get_a_mask_acc = dcache__GEN_200 | dcache_get_a_mask_size & dcache_get_a_mask_eq ; 
    wire dcache_get_a_mask_eq_1 = dcache_get_a_mask_bit &1'h1; 
    wire dcache_get_a_mask_acc_1 = dcache__GEN_200 | dcache_get_a_mask_size & dcache_get_a_mask_eq_1 ; 
    wire dcache_get_a_mask_size_1 = dcache_get_a_mask_sizeOH [1]; 
    wire dcache_get_a_mask_bit_1 = dcache_s2_req_addr [1]; 
    wire dcache_get_a_mask_nbit_1 = dcache_get_a_mask_bit_1 ==1'h0; 
    wire dcache_get_a_mask_eq_2 = dcache_get_a_mask_eq & dcache_get_a_mask_nbit_1 ; 
    wire dcache_get_a_mask_acc_2 = dcache_get_a_mask_acc | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_2 ; 
    wire dcache_get_a_mask_eq_3 = dcache_get_a_mask_eq & dcache_get_a_mask_bit_1 ; 
    wire dcache_get_a_mask_acc_3 = dcache_get_a_mask_acc | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_3 ; 
    wire dcache_get_a_mask_eq_4 = dcache_get_a_mask_eq_1 & dcache_get_a_mask_nbit_1 ; 
    wire dcache_get_a_mask_acc_4 = dcache_get_a_mask_acc_1 | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_4 ; 
    wire dcache_get_a_mask_eq_5 = dcache_get_a_mask_eq_1 & dcache_get_a_mask_bit_1 ; 
    wire dcache_get_a_mask_acc_5 = dcache_get_a_mask_acc_1 | dcache_get_a_mask_size_1 & dcache_get_a_mask_eq_5 ; 
    wire dcache_get_a_mask_size_2 = dcache_get_a_mask_sizeOH [0]; 
    wire dcache_get_a_mask_bit_2 = dcache_s2_req_addr [0]; 
    wire dcache_get_a_mask_nbit_2 = dcache_get_a_mask_bit_2 ==1'h0; 
    wire dcache_get_a_mask_eq_6 = dcache_get_a_mask_eq_2 & dcache_get_a_mask_nbit_2 ; 
    wire dcache_get_a_mask_acc_6 = dcache_get_a_mask_acc_2 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_6 ; 
    wire dcache_get_a_mask_eq_7 = dcache_get_a_mask_eq_2 & dcache_get_a_mask_bit_2 ; 
    wire dcache_get_a_mask_acc_7 = dcache_get_a_mask_acc_2 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_7 ; 
    wire dcache_get_a_mask_eq_8 = dcache_get_a_mask_eq_3 & dcache_get_a_mask_nbit_2 ; 
    wire dcache_get_a_mask_acc_8 = dcache_get_a_mask_acc_3 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_8 ; 
    wire dcache_get_a_mask_eq_9 = dcache_get_a_mask_eq_3 & dcache_get_a_mask_bit_2 ; 
    wire dcache_get_a_mask_acc_9 = dcache_get_a_mask_acc_3 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_9 ; 
    wire dcache_get_a_mask_eq_10 = dcache_get_a_mask_eq_4 & dcache_get_a_mask_nbit_2 ; 
    wire dcache_get_a_mask_acc_10 = dcache_get_a_mask_acc_4 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_10 ; 
    wire dcache_get_a_mask_eq_11 = dcache_get_a_mask_eq_4 & dcache_get_a_mask_bit_2 ; 
    wire dcache_get_a_mask_acc_11 = dcache_get_a_mask_acc_4 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_11 ; 
    wire dcache_get_a_mask_eq_12 = dcache_get_a_mask_eq_5 & dcache_get_a_mask_nbit_2 ; 
    wire dcache_get_a_mask_acc_12 = dcache_get_a_mask_acc_5 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_12 ; 
    wire dcache_get_a_mask_eq_13 = dcache_get_a_mask_eq_5 & dcache_get_a_mask_bit_2 ; 
    wire dcache_get_a_mask_acc_13 = dcache_get_a_mask_acc_5 | dcache_get_a_mask_size_2 & dcache_get_a_mask_eq_13 ; 
    wire[1:0] dcache_get_a_mask_lo_lo ={ dcache_get_a_mask_acc_7 , dcache_get_a_mask_acc_6 }; 
    wire[1:0] dcache_get_a_mask_lo_hi ={ dcache_get_a_mask_acc_9 , dcache_get_a_mask_acc_8 }; 
    wire[3:0] dcache_get_a_mask_lo ={ dcache_get_a_mask_lo_hi , dcache_get_a_mask_lo_lo }; 
    wire[1:0] dcache_get_a_mask_hi_lo ={ dcache_get_a_mask_acc_11 , dcache_get_a_mask_acc_10 }; 
    wire[1:0] dcache_get_a_mask_hi_hi ={ dcache_get_a_mask_acc_13 , dcache_get_a_mask_acc_12 }; 
    wire[3:0] dcache_get_a_mask_hi ={ dcache_get_a_mask_hi_hi , dcache_get_a_mask_hi_lo }; 
    wire[7:0] dcache_get_mask ={ dcache_get_a_mask_hi , dcache_get_a_mask_lo }; 
    wire[63:0] dcache_get_data =64'h0; 
    wire dcache_put_legal =(2'h0<= dcache_s2_req_size &{2'h0, dcache_s2_req_size }<=4'hC|1'h0)&({1'h0, dcache_s2_req_addr ^34'h2000}&35'hCA012000)==35'h0|1'h0|(2'h0<= dcache_s2_req_size &{1'h0, dcache_s2_req_size }<=3'h6|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hCA012000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h80000000}&35'hC0000000)==35'h0)|(2'h0<= dcache_s2_req_size &{2'h0, dcache_s2_req_size }<=4'h8|1'h0)&({1'h0, dcache_s2_req_addr ^34'h40000000}&35'hC0000000)==35'h0; 
    wire[2:0] dcache_put_opcode =3'h0; 
    wire[2:0] dcache_put_param =3'h0; 
    wire[3:0] dcache_put_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_put_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_201 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_put_a_mask_sizeOH_shiftAmount = dcache__GEN_201 [1:0]; 
    wire[3:0] dcache__GEN_202 =4'h1<< dcache_put_a_mask_sizeOH_shiftAmount ; 
    wire[2:0] dcache_put_a_mask_sizeOH = dcache__GEN_202 [2:0]|3'h1; 
    wire dcache__GEN_203 = dcache_s2_req_size >=2'h3; 
    wire dcache_put_a_mask_size = dcache_put_a_mask_sizeOH [2]; 
    wire dcache_put_a_mask_bit = dcache_s2_req_addr [2]; 
    wire dcache_put_a_mask_nbit = dcache_put_a_mask_bit ==1'h0; 
    wire dcache_put_a_mask_eq = dcache_put_a_mask_nbit &1'h1; 
    wire dcache_put_a_mask_acc = dcache__GEN_203 | dcache_put_a_mask_size & dcache_put_a_mask_eq ; 
    wire dcache_put_a_mask_eq_1 = dcache_put_a_mask_bit &1'h1; 
    wire dcache_put_a_mask_acc_1 = dcache__GEN_203 | dcache_put_a_mask_size & dcache_put_a_mask_eq_1 ; 
    wire dcache_put_a_mask_size_1 = dcache_put_a_mask_sizeOH [1]; 
    wire dcache_put_a_mask_bit_1 = dcache_s2_req_addr [1]; 
    wire dcache_put_a_mask_nbit_1 = dcache_put_a_mask_bit_1 ==1'h0; 
    wire dcache_put_a_mask_eq_2 = dcache_put_a_mask_eq & dcache_put_a_mask_nbit_1 ; 
    wire dcache_put_a_mask_acc_2 = dcache_put_a_mask_acc | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_2 ; 
    wire dcache_put_a_mask_eq_3 = dcache_put_a_mask_eq & dcache_put_a_mask_bit_1 ; 
    wire dcache_put_a_mask_acc_3 = dcache_put_a_mask_acc | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_3 ; 
    wire dcache_put_a_mask_eq_4 = dcache_put_a_mask_eq_1 & dcache_put_a_mask_nbit_1 ; 
    wire dcache_put_a_mask_acc_4 = dcache_put_a_mask_acc_1 | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_4 ; 
    wire dcache_put_a_mask_eq_5 = dcache_put_a_mask_eq_1 & dcache_put_a_mask_bit_1 ; 
    wire dcache_put_a_mask_acc_5 = dcache_put_a_mask_acc_1 | dcache_put_a_mask_size_1 & dcache_put_a_mask_eq_5 ; 
    wire dcache_put_a_mask_size_2 = dcache_put_a_mask_sizeOH [0]; 
    wire dcache_put_a_mask_bit_2 = dcache_s2_req_addr [0]; 
    wire dcache_put_a_mask_nbit_2 = dcache_put_a_mask_bit_2 ==1'h0; 
    wire dcache_put_a_mask_eq_6 = dcache_put_a_mask_eq_2 & dcache_put_a_mask_nbit_2 ; 
    wire dcache_put_a_mask_acc_6 = dcache_put_a_mask_acc_2 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_6 ; 
    wire dcache_put_a_mask_eq_7 = dcache_put_a_mask_eq_2 & dcache_put_a_mask_bit_2 ; 
    wire dcache_put_a_mask_acc_7 = dcache_put_a_mask_acc_2 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_7 ; 
    wire dcache_put_a_mask_eq_8 = dcache_put_a_mask_eq_3 & dcache_put_a_mask_nbit_2 ; 
    wire dcache_put_a_mask_acc_8 = dcache_put_a_mask_acc_3 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_8 ; 
    wire dcache_put_a_mask_eq_9 = dcache_put_a_mask_eq_3 & dcache_put_a_mask_bit_2 ; 
    wire dcache_put_a_mask_acc_9 = dcache_put_a_mask_acc_3 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_9 ; 
    wire dcache_put_a_mask_eq_10 = dcache_put_a_mask_eq_4 & dcache_put_a_mask_nbit_2 ; 
    wire dcache_put_a_mask_acc_10 = dcache_put_a_mask_acc_4 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_10 ; 
    wire dcache_put_a_mask_eq_11 = dcache_put_a_mask_eq_4 & dcache_put_a_mask_bit_2 ; 
    wire dcache_put_a_mask_acc_11 = dcache_put_a_mask_acc_4 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_11 ; 
    wire dcache_put_a_mask_eq_12 = dcache_put_a_mask_eq_5 & dcache_put_a_mask_nbit_2 ; 
    wire dcache_put_a_mask_acc_12 = dcache_put_a_mask_acc_5 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_12 ; 
    wire dcache_put_a_mask_eq_13 = dcache_put_a_mask_eq_5 & dcache_put_a_mask_bit_2 ; 
    wire dcache_put_a_mask_acc_13 = dcache_put_a_mask_acc_5 | dcache_put_a_mask_size_2 & dcache_put_a_mask_eq_13 ; 
    wire[1:0] dcache_put_a_mask_lo_lo ={ dcache_put_a_mask_acc_7 , dcache_put_a_mask_acc_6 }; 
    wire[1:0] dcache_put_a_mask_lo_hi ={ dcache_put_a_mask_acc_9 , dcache_put_a_mask_acc_8 }; 
    wire[3:0] dcache_put_a_mask_lo ={ dcache_put_a_mask_lo_hi , dcache_put_a_mask_lo_lo }; 
    wire[1:0] dcache_put_a_mask_hi_lo ={ dcache_put_a_mask_acc_11 , dcache_put_a_mask_acc_10 }; 
    wire[1:0] dcache_put_a_mask_hi_hi ={ dcache_put_a_mask_acc_13 , dcache_put_a_mask_acc_12 }; 
    wire[3:0] dcache_put_a_mask_hi ={ dcache_put_a_mask_hi_hi , dcache_put_a_mask_hi_lo }; 
    wire[7:0] dcache_put_mask ={ dcache_put_a_mask_hi , dcache_put_a_mask_lo }; 
    wire dcache_putpartial_legal =(2'h0<= dcache_s2_req_size &{2'h0, dcache_s2_req_size }<=4'hC|1'h0)&({1'h0, dcache_s2_req_addr ^34'h2000}&35'hCA012000)==35'h0|1'h0|(2'h0<= dcache_s2_req_size &{1'h0, dcache_s2_req_size }<=3'h6|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hCA012000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h80000000}&35'hC0000000)==35'h0)|(2'h0<= dcache_s2_req_size &{2'h0, dcache_s2_req_size }<=4'h8|1'h0)&({1'h0, dcache_s2_req_addr ^34'h40000000}&35'hC0000000)==35'h0; 
    wire[2:0] dcache_putpartial_opcode =3'h1; 
    wire[2:0] dcache_putpartial_param =3'h0; 
    wire[3:0] dcache_putpartial_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_putpartial_address = dcache_s2_req_addr [31:0]; 
    wire[7:0] dcache_putpartial_mask = dcache_a_mask [7:0]; 
    wire[2:0] dcache__atomics_WIRE_1_opcode = dcache__atomics_WIRE_opcode ; 
    wire[2:0] dcache__atomics_WIRE_1_param = dcache__atomics_WIRE_param ; 
    wire[3:0] dcache__atomics_WIRE_1_size = dcache__atomics_WIRE_size ; 
    wire dcache__atomics_WIRE_1_source = dcache__atomics_WIRE_source ; 
    wire[31:0] dcache__atomics_WIRE_1_address = dcache__atomics_WIRE_address ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_bufferable = dcache__atomics_WIRE_user_amba_prot_bufferable ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_modifiable = dcache__atomics_WIRE_user_amba_prot_modifiable ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_readalloc = dcache__atomics_WIRE_user_amba_prot_readalloc ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_writealloc = dcache__atomics_WIRE_user_amba_prot_writealloc ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_privileged = dcache__atomics_WIRE_user_amba_prot_privileged ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_secure = dcache__atomics_WIRE_user_amba_prot_secure ; 
    wire dcache__atomics_WIRE_1_user_amba_prot_fetch = dcache__atomics_WIRE_user_amba_prot_fetch ; 
    wire[7:0] dcache__atomics_WIRE_1_mask = dcache__atomics_WIRE_mask ; 
    wire[63:0] dcache__atomics_WIRE_1_data = dcache__atomics_WIRE_data ; 
    wire dcache__atomics_WIRE_1_corrupt = dcache__atomics_WIRE_corrupt ; 
    wire dcache_atomics_legal =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_opcode =3'h3; 
    wire[3:0] dcache_atomics_a_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_204 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount = dcache__GEN_204 [1:0]; 
    wire[3:0] dcache__GEN_205 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH = dcache__GEN_205 [2:0]|3'h1; 
    wire dcache__GEN_206 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size = dcache_atomics_a_mask_sizeOH [2]; 
    wire dcache_atomics_a_mask_bit = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit = dcache_atomics_a_mask_bit ==1'h0; 
    wire dcache_atomics_a_mask_eq = dcache_atomics_a_mask_nbit &1'h1; 
    wire dcache_atomics_a_mask_acc = dcache__GEN_206 | dcache_atomics_a_mask_size & dcache_atomics_a_mask_eq ; 
    wire dcache_atomics_a_mask_eq_1 = dcache_atomics_a_mask_bit &1'h1; 
    wire dcache_atomics_a_mask_acc_1 = dcache__GEN_206 | dcache_atomics_a_mask_size & dcache_atomics_a_mask_eq_1 ; 
    wire dcache_atomics_a_mask_size_1 = dcache_atomics_a_mask_sizeOH [1]; 
    wire dcache_atomics_a_mask_bit_1 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_1 = dcache_atomics_a_mask_bit_1 ==1'h0; 
    wire dcache_atomics_a_mask_eq_2 = dcache_atomics_a_mask_eq & dcache_atomics_a_mask_nbit_1 ; 
    wire dcache_atomics_a_mask_acc_2 = dcache_atomics_a_mask_acc | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_2 ; 
    wire dcache_atomics_a_mask_eq_3 = dcache_atomics_a_mask_eq & dcache_atomics_a_mask_bit_1 ; 
    wire dcache_atomics_a_mask_acc_3 = dcache_atomics_a_mask_acc | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_3 ; 
    wire dcache_atomics_a_mask_eq_4 = dcache_atomics_a_mask_eq_1 & dcache_atomics_a_mask_nbit_1 ; 
    wire dcache_atomics_a_mask_acc_4 = dcache_atomics_a_mask_acc_1 | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_4 ; 
    wire dcache_atomics_a_mask_eq_5 = dcache_atomics_a_mask_eq_1 & dcache_atomics_a_mask_bit_1 ; 
    wire dcache_atomics_a_mask_acc_5 = dcache_atomics_a_mask_acc_1 | dcache_atomics_a_mask_size_1 & dcache_atomics_a_mask_eq_5 ; 
    wire dcache_atomics_a_mask_size_2 = dcache_atomics_a_mask_sizeOH [0]; 
    wire dcache_atomics_a_mask_bit_2 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_2 = dcache_atomics_a_mask_bit_2 ==1'h0; 
    wire dcache_atomics_a_mask_eq_6 = dcache_atomics_a_mask_eq_2 & dcache_atomics_a_mask_nbit_2 ; 
    wire dcache_atomics_a_mask_acc_6 = dcache_atomics_a_mask_acc_2 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_6 ; 
    wire dcache_atomics_a_mask_eq_7 = dcache_atomics_a_mask_eq_2 & dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_acc_7 = dcache_atomics_a_mask_acc_2 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_7 ; 
    wire dcache_atomics_a_mask_eq_8 = dcache_atomics_a_mask_eq_3 & dcache_atomics_a_mask_nbit_2 ; 
    wire dcache_atomics_a_mask_acc_8 = dcache_atomics_a_mask_acc_3 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_8 ; 
    wire dcache_atomics_a_mask_eq_9 = dcache_atomics_a_mask_eq_3 & dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_acc_9 = dcache_atomics_a_mask_acc_3 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_9 ; 
    wire dcache_atomics_a_mask_eq_10 = dcache_atomics_a_mask_eq_4 & dcache_atomics_a_mask_nbit_2 ; 
    wire dcache_atomics_a_mask_acc_10 = dcache_atomics_a_mask_acc_4 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_10 ; 
    wire dcache_atomics_a_mask_eq_11 = dcache_atomics_a_mask_eq_4 & dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_acc_11 = dcache_atomics_a_mask_acc_4 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_11 ; 
    wire dcache_atomics_a_mask_eq_12 = dcache_atomics_a_mask_eq_5 & dcache_atomics_a_mask_nbit_2 ; 
    wire dcache_atomics_a_mask_acc_12 = dcache_atomics_a_mask_acc_5 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_12 ; 
    wire dcache_atomics_a_mask_eq_13 = dcache_atomics_a_mask_eq_5 & dcache_atomics_a_mask_bit_2 ; 
    wire dcache_atomics_a_mask_acc_13 = dcache_atomics_a_mask_acc_5 | dcache_atomics_a_mask_size_2 & dcache_atomics_a_mask_eq_13 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo ={ dcache_atomics_a_mask_acc_7 , dcache_atomics_a_mask_acc_6 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi ={ dcache_atomics_a_mask_acc_9 , dcache_atomics_a_mask_acc_8 }; 
    wire[3:0] dcache_atomics_a_mask_lo ={ dcache_atomics_a_mask_lo_hi , dcache_atomics_a_mask_lo_lo }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo ={ dcache_atomics_a_mask_acc_11 , dcache_atomics_a_mask_acc_10 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi ={ dcache_atomics_a_mask_acc_13 , dcache_atomics_a_mask_acc_12 }; 
    wire[3:0] dcache_atomics_a_mask_hi ={ dcache_atomics_a_mask_hi_hi , dcache_atomics_a_mask_hi_lo }; 
    wire[7:0] dcache_atomics_a_mask ={ dcache_atomics_a_mask_hi , dcache_atomics_a_mask_lo }; 
    wire dcache_atomics_legal_1 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_1_opcode =3'h3; 
    wire[3:0] dcache_atomics_a_1_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_1_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_207 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_1 = dcache__GEN_207 [1:0]; 
    wire[3:0] dcache__GEN_208 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_1 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_1 = dcache__GEN_208 [2:0]|3'h1; 
    wire dcache__GEN_209 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_3 = dcache_atomics_a_mask_sizeOH_1 [2]; 
    wire dcache_atomics_a_mask_bit_3 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_3 = dcache_atomics_a_mask_bit_3 ==1'h0; 
    wire dcache_atomics_a_mask_eq_14 = dcache_atomics_a_mask_nbit_3 &1'h1; 
    wire dcache_atomics_a_mask_acc_14 = dcache__GEN_209 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_14 ; 
    wire dcache_atomics_a_mask_eq_15 = dcache_atomics_a_mask_bit_3 &1'h1; 
    wire dcache_atomics_a_mask_acc_15 = dcache__GEN_209 | dcache_atomics_a_mask_size_3 & dcache_atomics_a_mask_eq_15 ; 
    wire dcache_atomics_a_mask_size_4 = dcache_atomics_a_mask_sizeOH_1 [1]; 
    wire dcache_atomics_a_mask_bit_4 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_4 = dcache_atomics_a_mask_bit_4 ==1'h0; 
    wire dcache_atomics_a_mask_eq_16 = dcache_atomics_a_mask_eq_14 & dcache_atomics_a_mask_nbit_4 ; 
    wire dcache_atomics_a_mask_acc_16 = dcache_atomics_a_mask_acc_14 | dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_16 ; 
    wire dcache_atomics_a_mask_eq_17 = dcache_atomics_a_mask_eq_14 & dcache_atomics_a_mask_bit_4 ; 
    wire dcache_atomics_a_mask_acc_17 = dcache_atomics_a_mask_acc_14 | dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_17 ; 
    wire dcache_atomics_a_mask_eq_18 = dcache_atomics_a_mask_eq_15 & dcache_atomics_a_mask_nbit_4 ; 
    wire dcache_atomics_a_mask_acc_18 = dcache_atomics_a_mask_acc_15 | dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_18 ; 
    wire dcache_atomics_a_mask_eq_19 = dcache_atomics_a_mask_eq_15 & dcache_atomics_a_mask_bit_4 ; 
    wire dcache_atomics_a_mask_acc_19 = dcache_atomics_a_mask_acc_15 | dcache_atomics_a_mask_size_4 & dcache_atomics_a_mask_eq_19 ; 
    wire dcache_atomics_a_mask_size_5 = dcache_atomics_a_mask_sizeOH_1 [0]; 
    wire dcache_atomics_a_mask_bit_5 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_5 = dcache_atomics_a_mask_bit_5 ==1'h0; 
    wire dcache_atomics_a_mask_eq_20 = dcache_atomics_a_mask_eq_16 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_20 = dcache_atomics_a_mask_acc_16 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_20 ; 
    wire dcache_atomics_a_mask_eq_21 = dcache_atomics_a_mask_eq_16 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_21 = dcache_atomics_a_mask_acc_16 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_21 ; 
    wire dcache_atomics_a_mask_eq_22 = dcache_atomics_a_mask_eq_17 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_22 = dcache_atomics_a_mask_acc_17 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_22 ; 
    wire dcache_atomics_a_mask_eq_23 = dcache_atomics_a_mask_eq_17 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_23 = dcache_atomics_a_mask_acc_17 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_23 ; 
    wire dcache_atomics_a_mask_eq_24 = dcache_atomics_a_mask_eq_18 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_24 = dcache_atomics_a_mask_acc_18 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_24 ; 
    wire dcache_atomics_a_mask_eq_25 = dcache_atomics_a_mask_eq_18 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_25 = dcache_atomics_a_mask_acc_18 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_25 ; 
    wire dcache_atomics_a_mask_eq_26 = dcache_atomics_a_mask_eq_19 & dcache_atomics_a_mask_nbit_5 ; 
    wire dcache_atomics_a_mask_acc_26 = dcache_atomics_a_mask_acc_19 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_26 ; 
    wire dcache_atomics_a_mask_eq_27 = dcache_atomics_a_mask_eq_19 & dcache_atomics_a_mask_bit_5 ; 
    wire dcache_atomics_a_mask_acc_27 = dcache_atomics_a_mask_acc_19 | dcache_atomics_a_mask_size_5 & dcache_atomics_a_mask_eq_27 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_1 ={ dcache_atomics_a_mask_acc_21 , dcache_atomics_a_mask_acc_20 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_1 ={ dcache_atomics_a_mask_acc_23 , dcache_atomics_a_mask_acc_22 }; 
    wire[3:0] dcache_atomics_a_mask_lo_1 ={ dcache_atomics_a_mask_lo_hi_1 , dcache_atomics_a_mask_lo_lo_1 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_1 ={ dcache_atomics_a_mask_acc_25 , dcache_atomics_a_mask_acc_24 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_1 ={ dcache_atomics_a_mask_acc_27 , dcache_atomics_a_mask_acc_26 }; 
    wire[3:0] dcache_atomics_a_mask_hi_1 ={ dcache_atomics_a_mask_hi_hi_1 , dcache_atomics_a_mask_hi_lo_1 }; 
    wire[7:0] dcache_atomics_a_1_mask ={ dcache_atomics_a_mask_hi_1 , dcache_atomics_a_mask_lo_1 }; 
    wire dcache_atomics_legal_2 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_2_opcode =3'h3; 
    wire[3:0] dcache_atomics_a_2_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_2_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_210 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_2 = dcache__GEN_210 [1:0]; 
    wire[3:0] dcache__GEN_211 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_2 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_2 = dcache__GEN_211 [2:0]|3'h1; 
    wire dcache__GEN_212 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_6 = dcache_atomics_a_mask_sizeOH_2 [2]; 
    wire dcache_atomics_a_mask_bit_6 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_6 = dcache_atomics_a_mask_bit_6 ==1'h0; 
    wire dcache_atomics_a_mask_eq_28 = dcache_atomics_a_mask_nbit_6 &1'h1; 
    wire dcache_atomics_a_mask_acc_28 = dcache__GEN_212 | dcache_atomics_a_mask_size_6 & dcache_atomics_a_mask_eq_28 ; 
    wire dcache_atomics_a_mask_eq_29 = dcache_atomics_a_mask_bit_6 &1'h1; 
    wire dcache_atomics_a_mask_acc_29 = dcache__GEN_212 | dcache_atomics_a_mask_size_6 & dcache_atomics_a_mask_eq_29 ; 
    wire dcache_atomics_a_mask_size_7 = dcache_atomics_a_mask_sizeOH_2 [1]; 
    wire dcache_atomics_a_mask_bit_7 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_7 = dcache_atomics_a_mask_bit_7 ==1'h0; 
    wire dcache_atomics_a_mask_eq_30 = dcache_atomics_a_mask_eq_28 & dcache_atomics_a_mask_nbit_7 ; 
    wire dcache_atomics_a_mask_acc_30 = dcache_atomics_a_mask_acc_28 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_30 ; 
    wire dcache_atomics_a_mask_eq_31 = dcache_atomics_a_mask_eq_28 & dcache_atomics_a_mask_bit_7 ; 
    wire dcache_atomics_a_mask_acc_31 = dcache_atomics_a_mask_acc_28 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_31 ; 
    wire dcache_atomics_a_mask_eq_32 = dcache_atomics_a_mask_eq_29 & dcache_atomics_a_mask_nbit_7 ; 
    wire dcache_atomics_a_mask_acc_32 = dcache_atomics_a_mask_acc_29 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_32 ; 
    wire dcache_atomics_a_mask_eq_33 = dcache_atomics_a_mask_eq_29 & dcache_atomics_a_mask_bit_7 ; 
    wire dcache_atomics_a_mask_acc_33 = dcache_atomics_a_mask_acc_29 | dcache_atomics_a_mask_size_7 & dcache_atomics_a_mask_eq_33 ; 
    wire dcache_atomics_a_mask_size_8 = dcache_atomics_a_mask_sizeOH_2 [0]; 
    wire dcache_atomics_a_mask_bit_8 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_8 = dcache_atomics_a_mask_bit_8 ==1'h0; 
    wire dcache_atomics_a_mask_eq_34 = dcache_atomics_a_mask_eq_30 & dcache_atomics_a_mask_nbit_8 ; 
    wire dcache_atomics_a_mask_acc_34 = dcache_atomics_a_mask_acc_30 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_34 ; 
    wire dcache_atomics_a_mask_eq_35 = dcache_atomics_a_mask_eq_30 & dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_acc_35 = dcache_atomics_a_mask_acc_30 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_35 ; 
    wire dcache_atomics_a_mask_eq_36 = dcache_atomics_a_mask_eq_31 & dcache_atomics_a_mask_nbit_8 ; 
    wire dcache_atomics_a_mask_acc_36 = dcache_atomics_a_mask_acc_31 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_36 ; 
    wire dcache_atomics_a_mask_eq_37 = dcache_atomics_a_mask_eq_31 & dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_acc_37 = dcache_atomics_a_mask_acc_31 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_37 ; 
    wire dcache_atomics_a_mask_eq_38 = dcache_atomics_a_mask_eq_32 & dcache_atomics_a_mask_nbit_8 ; 
    wire dcache_atomics_a_mask_acc_38 = dcache_atomics_a_mask_acc_32 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_38 ; 
    wire dcache_atomics_a_mask_eq_39 = dcache_atomics_a_mask_eq_32 & dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_acc_39 = dcache_atomics_a_mask_acc_32 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_39 ; 
    wire dcache_atomics_a_mask_eq_40 = dcache_atomics_a_mask_eq_33 & dcache_atomics_a_mask_nbit_8 ; 
    wire dcache_atomics_a_mask_acc_40 = dcache_atomics_a_mask_acc_33 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_40 ; 
    wire dcache_atomics_a_mask_eq_41 = dcache_atomics_a_mask_eq_33 & dcache_atomics_a_mask_bit_8 ; 
    wire dcache_atomics_a_mask_acc_41 = dcache_atomics_a_mask_acc_33 | dcache_atomics_a_mask_size_8 & dcache_atomics_a_mask_eq_41 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_2 ={ dcache_atomics_a_mask_acc_35 , dcache_atomics_a_mask_acc_34 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_2 ={ dcache_atomics_a_mask_acc_37 , dcache_atomics_a_mask_acc_36 }; 
    wire[3:0] dcache_atomics_a_mask_lo_2 ={ dcache_atomics_a_mask_lo_hi_2 , dcache_atomics_a_mask_lo_lo_2 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_2 ={ dcache_atomics_a_mask_acc_39 , dcache_atomics_a_mask_acc_38 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_2 ={ dcache_atomics_a_mask_acc_41 , dcache_atomics_a_mask_acc_40 }; 
    wire[3:0] dcache_atomics_a_mask_hi_2 ={ dcache_atomics_a_mask_hi_hi_2 , dcache_atomics_a_mask_hi_lo_2 }; 
    wire[7:0] dcache_atomics_a_2_mask ={ dcache_atomics_a_mask_hi_2 , dcache_atomics_a_mask_lo_2 }; 
    wire dcache_atomics_legal_3 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_3_opcode =3'h3; 
    wire[3:0] dcache_atomics_a_3_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_3_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_213 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_3 = dcache__GEN_213 [1:0]; 
    wire[3:0] dcache__GEN_214 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_3 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_3 = dcache__GEN_214 [2:0]|3'h1; 
    wire dcache__GEN_215 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_9 = dcache_atomics_a_mask_sizeOH_3 [2]; 
    wire dcache_atomics_a_mask_bit_9 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_9 = dcache_atomics_a_mask_bit_9 ==1'h0; 
    wire dcache_atomics_a_mask_eq_42 = dcache_atomics_a_mask_nbit_9 &1'h1; 
    wire dcache_atomics_a_mask_acc_42 = dcache__GEN_215 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_42 ; 
    wire dcache_atomics_a_mask_eq_43 = dcache_atomics_a_mask_bit_9 &1'h1; 
    wire dcache_atomics_a_mask_acc_43 = dcache__GEN_215 | dcache_atomics_a_mask_size_9 & dcache_atomics_a_mask_eq_43 ; 
    wire dcache_atomics_a_mask_size_10 = dcache_atomics_a_mask_sizeOH_3 [1]; 
    wire dcache_atomics_a_mask_bit_10 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_10 = dcache_atomics_a_mask_bit_10 ==1'h0; 
    wire dcache_atomics_a_mask_eq_44 = dcache_atomics_a_mask_eq_42 & dcache_atomics_a_mask_nbit_10 ; 
    wire dcache_atomics_a_mask_acc_44 = dcache_atomics_a_mask_acc_42 | dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_44 ; 
    wire dcache_atomics_a_mask_eq_45 = dcache_atomics_a_mask_eq_42 & dcache_atomics_a_mask_bit_10 ; 
    wire dcache_atomics_a_mask_acc_45 = dcache_atomics_a_mask_acc_42 | dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_45 ; 
    wire dcache_atomics_a_mask_eq_46 = dcache_atomics_a_mask_eq_43 & dcache_atomics_a_mask_nbit_10 ; 
    wire dcache_atomics_a_mask_acc_46 = dcache_atomics_a_mask_acc_43 | dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_46 ; 
    wire dcache_atomics_a_mask_eq_47 = dcache_atomics_a_mask_eq_43 & dcache_atomics_a_mask_bit_10 ; 
    wire dcache_atomics_a_mask_acc_47 = dcache_atomics_a_mask_acc_43 | dcache_atomics_a_mask_size_10 & dcache_atomics_a_mask_eq_47 ; 
    wire dcache_atomics_a_mask_size_11 = dcache_atomics_a_mask_sizeOH_3 [0]; 
    wire dcache_atomics_a_mask_bit_11 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_11 = dcache_atomics_a_mask_bit_11 ==1'h0; 
    wire dcache_atomics_a_mask_eq_48 = dcache_atomics_a_mask_eq_44 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_48 = dcache_atomics_a_mask_acc_44 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_48 ; 
    wire dcache_atomics_a_mask_eq_49 = dcache_atomics_a_mask_eq_44 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_49 = dcache_atomics_a_mask_acc_44 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_49 ; 
    wire dcache_atomics_a_mask_eq_50 = dcache_atomics_a_mask_eq_45 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_50 = dcache_atomics_a_mask_acc_45 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_50 ; 
    wire dcache_atomics_a_mask_eq_51 = dcache_atomics_a_mask_eq_45 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_51 = dcache_atomics_a_mask_acc_45 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_51 ; 
    wire dcache_atomics_a_mask_eq_52 = dcache_atomics_a_mask_eq_46 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_52 = dcache_atomics_a_mask_acc_46 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_52 ; 
    wire dcache_atomics_a_mask_eq_53 = dcache_atomics_a_mask_eq_46 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_53 = dcache_atomics_a_mask_acc_46 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_53 ; 
    wire dcache_atomics_a_mask_eq_54 = dcache_atomics_a_mask_eq_47 & dcache_atomics_a_mask_nbit_11 ; 
    wire dcache_atomics_a_mask_acc_54 = dcache_atomics_a_mask_acc_47 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_54 ; 
    wire dcache_atomics_a_mask_eq_55 = dcache_atomics_a_mask_eq_47 & dcache_atomics_a_mask_bit_11 ; 
    wire dcache_atomics_a_mask_acc_55 = dcache_atomics_a_mask_acc_47 | dcache_atomics_a_mask_size_11 & dcache_atomics_a_mask_eq_55 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_3 ={ dcache_atomics_a_mask_acc_49 , dcache_atomics_a_mask_acc_48 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_3 ={ dcache_atomics_a_mask_acc_51 , dcache_atomics_a_mask_acc_50 }; 
    wire[3:0] dcache_atomics_a_mask_lo_3 ={ dcache_atomics_a_mask_lo_hi_3 , dcache_atomics_a_mask_lo_lo_3 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_3 ={ dcache_atomics_a_mask_acc_53 , dcache_atomics_a_mask_acc_52 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_3 ={ dcache_atomics_a_mask_acc_55 , dcache_atomics_a_mask_acc_54 }; 
    wire[3:0] dcache_atomics_a_mask_hi_3 ={ dcache_atomics_a_mask_hi_hi_3 , dcache_atomics_a_mask_hi_lo_3 }; 
    wire[7:0] dcache_atomics_a_3_mask ={ dcache_atomics_a_mask_hi_3 , dcache_atomics_a_mask_lo_3 }; 
    wire dcache_atomics_legal_4 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_4_opcode =3'h2; 
    wire[3:0] dcache_atomics_a_4_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_4_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_216 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_4 = dcache__GEN_216 [1:0]; 
    wire[3:0] dcache__GEN_217 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_4 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_4 = dcache__GEN_217 [2:0]|3'h1; 
    wire dcache__GEN_218 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_12 = dcache_atomics_a_mask_sizeOH_4 [2]; 
    wire dcache_atomics_a_mask_bit_12 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_12 = dcache_atomics_a_mask_bit_12 ==1'h0; 
    wire dcache_atomics_a_mask_eq_56 = dcache_atomics_a_mask_nbit_12 &1'h1; 
    wire dcache_atomics_a_mask_acc_56 = dcache__GEN_218 | dcache_atomics_a_mask_size_12 & dcache_atomics_a_mask_eq_56 ; 
    wire dcache_atomics_a_mask_eq_57 = dcache_atomics_a_mask_bit_12 &1'h1; 
    wire dcache_atomics_a_mask_acc_57 = dcache__GEN_218 | dcache_atomics_a_mask_size_12 & dcache_atomics_a_mask_eq_57 ; 
    wire dcache_atomics_a_mask_size_13 = dcache_atomics_a_mask_sizeOH_4 [1]; 
    wire dcache_atomics_a_mask_bit_13 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_13 = dcache_atomics_a_mask_bit_13 ==1'h0; 
    wire dcache_atomics_a_mask_eq_58 = dcache_atomics_a_mask_eq_56 & dcache_atomics_a_mask_nbit_13 ; 
    wire dcache_atomics_a_mask_acc_58 = dcache_atomics_a_mask_acc_56 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_58 ; 
    wire dcache_atomics_a_mask_eq_59 = dcache_atomics_a_mask_eq_56 & dcache_atomics_a_mask_bit_13 ; 
    wire dcache_atomics_a_mask_acc_59 = dcache_atomics_a_mask_acc_56 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_59 ; 
    wire dcache_atomics_a_mask_eq_60 = dcache_atomics_a_mask_eq_57 & dcache_atomics_a_mask_nbit_13 ; 
    wire dcache_atomics_a_mask_acc_60 = dcache_atomics_a_mask_acc_57 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_60 ; 
    wire dcache_atomics_a_mask_eq_61 = dcache_atomics_a_mask_eq_57 & dcache_atomics_a_mask_bit_13 ; 
    wire dcache_atomics_a_mask_acc_61 = dcache_atomics_a_mask_acc_57 | dcache_atomics_a_mask_size_13 & dcache_atomics_a_mask_eq_61 ; 
    wire dcache_atomics_a_mask_size_14 = dcache_atomics_a_mask_sizeOH_4 [0]; 
    wire dcache_atomics_a_mask_bit_14 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_14 = dcache_atomics_a_mask_bit_14 ==1'h0; 
    wire dcache_atomics_a_mask_eq_62 = dcache_atomics_a_mask_eq_58 & dcache_atomics_a_mask_nbit_14 ; 
    wire dcache_atomics_a_mask_acc_62 = dcache_atomics_a_mask_acc_58 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_62 ; 
    wire dcache_atomics_a_mask_eq_63 = dcache_atomics_a_mask_eq_58 & dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_acc_63 = dcache_atomics_a_mask_acc_58 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_63 ; 
    wire dcache_atomics_a_mask_eq_64 = dcache_atomics_a_mask_eq_59 & dcache_atomics_a_mask_nbit_14 ; 
    wire dcache_atomics_a_mask_acc_64 = dcache_atomics_a_mask_acc_59 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_64 ; 
    wire dcache_atomics_a_mask_eq_65 = dcache_atomics_a_mask_eq_59 & dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_acc_65 = dcache_atomics_a_mask_acc_59 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_65 ; 
    wire dcache_atomics_a_mask_eq_66 = dcache_atomics_a_mask_eq_60 & dcache_atomics_a_mask_nbit_14 ; 
    wire dcache_atomics_a_mask_acc_66 = dcache_atomics_a_mask_acc_60 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_66 ; 
    wire dcache_atomics_a_mask_eq_67 = dcache_atomics_a_mask_eq_60 & dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_acc_67 = dcache_atomics_a_mask_acc_60 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_67 ; 
    wire dcache_atomics_a_mask_eq_68 = dcache_atomics_a_mask_eq_61 & dcache_atomics_a_mask_nbit_14 ; 
    wire dcache_atomics_a_mask_acc_68 = dcache_atomics_a_mask_acc_61 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_68 ; 
    wire dcache_atomics_a_mask_eq_69 = dcache_atomics_a_mask_eq_61 & dcache_atomics_a_mask_bit_14 ; 
    wire dcache_atomics_a_mask_acc_69 = dcache_atomics_a_mask_acc_61 | dcache_atomics_a_mask_size_14 & dcache_atomics_a_mask_eq_69 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_4 ={ dcache_atomics_a_mask_acc_63 , dcache_atomics_a_mask_acc_62 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_4 ={ dcache_atomics_a_mask_acc_65 , dcache_atomics_a_mask_acc_64 }; 
    wire[3:0] dcache_atomics_a_mask_lo_4 ={ dcache_atomics_a_mask_lo_hi_4 , dcache_atomics_a_mask_lo_lo_4 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_4 ={ dcache_atomics_a_mask_acc_67 , dcache_atomics_a_mask_acc_66 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_4 ={ dcache_atomics_a_mask_acc_69 , dcache_atomics_a_mask_acc_68 }; 
    wire[3:0] dcache_atomics_a_mask_hi_4 ={ dcache_atomics_a_mask_hi_hi_4 , dcache_atomics_a_mask_hi_lo_4 }; 
    wire[7:0] dcache_atomics_a_4_mask ={ dcache_atomics_a_mask_hi_4 , dcache_atomics_a_mask_lo_4 }; 
    wire dcache_atomics_legal_5 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_5_opcode =3'h2; 
    wire[3:0] dcache_atomics_a_5_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_5_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_219 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_5 = dcache__GEN_219 [1:0]; 
    wire[3:0] dcache__GEN_220 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_5 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_5 = dcache__GEN_220 [2:0]|3'h1; 
    wire dcache__GEN_221 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_15 = dcache_atomics_a_mask_sizeOH_5 [2]; 
    wire dcache_atomics_a_mask_bit_15 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_15 = dcache_atomics_a_mask_bit_15 ==1'h0; 
    wire dcache_atomics_a_mask_eq_70 = dcache_atomics_a_mask_nbit_15 &1'h1; 
    wire dcache_atomics_a_mask_acc_70 = dcache__GEN_221 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_70 ; 
    wire dcache_atomics_a_mask_eq_71 = dcache_atomics_a_mask_bit_15 &1'h1; 
    wire dcache_atomics_a_mask_acc_71 = dcache__GEN_221 | dcache_atomics_a_mask_size_15 & dcache_atomics_a_mask_eq_71 ; 
    wire dcache_atomics_a_mask_size_16 = dcache_atomics_a_mask_sizeOH_5 [1]; 
    wire dcache_atomics_a_mask_bit_16 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_16 = dcache_atomics_a_mask_bit_16 ==1'h0; 
    wire dcache_atomics_a_mask_eq_72 = dcache_atomics_a_mask_eq_70 & dcache_atomics_a_mask_nbit_16 ; 
    wire dcache_atomics_a_mask_acc_72 = dcache_atomics_a_mask_acc_70 | dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_72 ; 
    wire dcache_atomics_a_mask_eq_73 = dcache_atomics_a_mask_eq_70 & dcache_atomics_a_mask_bit_16 ; 
    wire dcache_atomics_a_mask_acc_73 = dcache_atomics_a_mask_acc_70 | dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_73 ; 
    wire dcache_atomics_a_mask_eq_74 = dcache_atomics_a_mask_eq_71 & dcache_atomics_a_mask_nbit_16 ; 
    wire dcache_atomics_a_mask_acc_74 = dcache_atomics_a_mask_acc_71 | dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_74 ; 
    wire dcache_atomics_a_mask_eq_75 = dcache_atomics_a_mask_eq_71 & dcache_atomics_a_mask_bit_16 ; 
    wire dcache_atomics_a_mask_acc_75 = dcache_atomics_a_mask_acc_71 | dcache_atomics_a_mask_size_16 & dcache_atomics_a_mask_eq_75 ; 
    wire dcache_atomics_a_mask_size_17 = dcache_atomics_a_mask_sizeOH_5 [0]; 
    wire dcache_atomics_a_mask_bit_17 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_17 = dcache_atomics_a_mask_bit_17 ==1'h0; 
    wire dcache_atomics_a_mask_eq_76 = dcache_atomics_a_mask_eq_72 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_76 = dcache_atomics_a_mask_acc_72 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_76 ; 
    wire dcache_atomics_a_mask_eq_77 = dcache_atomics_a_mask_eq_72 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_77 = dcache_atomics_a_mask_acc_72 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_77 ; 
    wire dcache_atomics_a_mask_eq_78 = dcache_atomics_a_mask_eq_73 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_78 = dcache_atomics_a_mask_acc_73 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_78 ; 
    wire dcache_atomics_a_mask_eq_79 = dcache_atomics_a_mask_eq_73 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_79 = dcache_atomics_a_mask_acc_73 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_79 ; 
    wire dcache_atomics_a_mask_eq_80 = dcache_atomics_a_mask_eq_74 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_80 = dcache_atomics_a_mask_acc_74 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_80 ; 
    wire dcache_atomics_a_mask_eq_81 = dcache_atomics_a_mask_eq_74 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_81 = dcache_atomics_a_mask_acc_74 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_81 ; 
    wire dcache_atomics_a_mask_eq_82 = dcache_atomics_a_mask_eq_75 & dcache_atomics_a_mask_nbit_17 ; 
    wire dcache_atomics_a_mask_acc_82 = dcache_atomics_a_mask_acc_75 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_82 ; 
    wire dcache_atomics_a_mask_eq_83 = dcache_atomics_a_mask_eq_75 & dcache_atomics_a_mask_bit_17 ; 
    wire dcache_atomics_a_mask_acc_83 = dcache_atomics_a_mask_acc_75 | dcache_atomics_a_mask_size_17 & dcache_atomics_a_mask_eq_83 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_5 ={ dcache_atomics_a_mask_acc_77 , dcache_atomics_a_mask_acc_76 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_5 ={ dcache_atomics_a_mask_acc_79 , dcache_atomics_a_mask_acc_78 }; 
    wire[3:0] dcache_atomics_a_mask_lo_5 ={ dcache_atomics_a_mask_lo_hi_5 , dcache_atomics_a_mask_lo_lo_5 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_5 ={ dcache_atomics_a_mask_acc_81 , dcache_atomics_a_mask_acc_80 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_5 ={ dcache_atomics_a_mask_acc_83 , dcache_atomics_a_mask_acc_82 }; 
    wire[3:0] dcache_atomics_a_mask_hi_5 ={ dcache_atomics_a_mask_hi_hi_5 , dcache_atomics_a_mask_hi_lo_5 }; 
    wire[7:0] dcache_atomics_a_5_mask ={ dcache_atomics_a_mask_hi_5 , dcache_atomics_a_mask_lo_5 }; 
    wire dcache_atomics_legal_6 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_6_opcode =3'h2; 
    wire[3:0] dcache_atomics_a_6_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_6_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_222 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_6 = dcache__GEN_222 [1:0]; 
    wire[3:0] dcache__GEN_223 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_6 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_6 = dcache__GEN_223 [2:0]|3'h1; 
    wire dcache__GEN_224 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_18 = dcache_atomics_a_mask_sizeOH_6 [2]; 
    wire dcache_atomics_a_mask_bit_18 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_18 = dcache_atomics_a_mask_bit_18 ==1'h0; 
    wire dcache_atomics_a_mask_eq_84 = dcache_atomics_a_mask_nbit_18 &1'h1; 
    wire dcache_atomics_a_mask_acc_84 = dcache__GEN_224 | dcache_atomics_a_mask_size_18 & dcache_atomics_a_mask_eq_84 ; 
    wire dcache_atomics_a_mask_eq_85 = dcache_atomics_a_mask_bit_18 &1'h1; 
    wire dcache_atomics_a_mask_acc_85 = dcache__GEN_224 | dcache_atomics_a_mask_size_18 & dcache_atomics_a_mask_eq_85 ; 
    wire dcache_atomics_a_mask_size_19 = dcache_atomics_a_mask_sizeOH_6 [1]; 
    wire dcache_atomics_a_mask_bit_19 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_19 = dcache_atomics_a_mask_bit_19 ==1'h0; 
    wire dcache_atomics_a_mask_eq_86 = dcache_atomics_a_mask_eq_84 & dcache_atomics_a_mask_nbit_19 ; 
    wire dcache_atomics_a_mask_acc_86 = dcache_atomics_a_mask_acc_84 | dcache_atomics_a_mask_size_19 & dcache_atomics_a_mask_eq_86 ; 
    wire dcache_atomics_a_mask_eq_87 = dcache_atomics_a_mask_eq_84 & dcache_atomics_a_mask_bit_19 ; 
    wire dcache_atomics_a_mask_acc_87 = dcache_atomics_a_mask_acc_84 | dcache_atomics_a_mask_size_19 & dcache_atomics_a_mask_eq_87 ; 
    wire dcache_atomics_a_mask_eq_88 = dcache_atomics_a_mask_eq_85 & dcache_atomics_a_mask_nbit_19 ; 
    wire dcache_atomics_a_mask_acc_88 = dcache_atomics_a_mask_acc_85 | dcache_atomics_a_mask_size_19 & dcache_atomics_a_mask_eq_88 ; 
    wire dcache_atomics_a_mask_eq_89 = dcache_atomics_a_mask_eq_85 & dcache_atomics_a_mask_bit_19 ; 
    wire dcache_atomics_a_mask_acc_89 = dcache_atomics_a_mask_acc_85 | dcache_atomics_a_mask_size_19 & dcache_atomics_a_mask_eq_89 ; 
    wire dcache_atomics_a_mask_size_20 = dcache_atomics_a_mask_sizeOH_6 [0]; 
    wire dcache_atomics_a_mask_bit_20 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_20 = dcache_atomics_a_mask_bit_20 ==1'h0; 
    wire dcache_atomics_a_mask_eq_90 = dcache_atomics_a_mask_eq_86 & dcache_atomics_a_mask_nbit_20 ; 
    wire dcache_atomics_a_mask_acc_90 = dcache_atomics_a_mask_acc_86 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_90 ; 
    wire dcache_atomics_a_mask_eq_91 = dcache_atomics_a_mask_eq_86 & dcache_atomics_a_mask_bit_20 ; 
    wire dcache_atomics_a_mask_acc_91 = dcache_atomics_a_mask_acc_86 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_91 ; 
    wire dcache_atomics_a_mask_eq_92 = dcache_atomics_a_mask_eq_87 & dcache_atomics_a_mask_nbit_20 ; 
    wire dcache_atomics_a_mask_acc_92 = dcache_atomics_a_mask_acc_87 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_92 ; 
    wire dcache_atomics_a_mask_eq_93 = dcache_atomics_a_mask_eq_87 & dcache_atomics_a_mask_bit_20 ; 
    wire dcache_atomics_a_mask_acc_93 = dcache_atomics_a_mask_acc_87 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_93 ; 
    wire dcache_atomics_a_mask_eq_94 = dcache_atomics_a_mask_eq_88 & dcache_atomics_a_mask_nbit_20 ; 
    wire dcache_atomics_a_mask_acc_94 = dcache_atomics_a_mask_acc_88 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_94 ; 
    wire dcache_atomics_a_mask_eq_95 = dcache_atomics_a_mask_eq_88 & dcache_atomics_a_mask_bit_20 ; 
    wire dcache_atomics_a_mask_acc_95 = dcache_atomics_a_mask_acc_88 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_95 ; 
    wire dcache_atomics_a_mask_eq_96 = dcache_atomics_a_mask_eq_89 & dcache_atomics_a_mask_nbit_20 ; 
    wire dcache_atomics_a_mask_acc_96 = dcache_atomics_a_mask_acc_89 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_96 ; 
    wire dcache_atomics_a_mask_eq_97 = dcache_atomics_a_mask_eq_89 & dcache_atomics_a_mask_bit_20 ; 
    wire dcache_atomics_a_mask_acc_97 = dcache_atomics_a_mask_acc_89 | dcache_atomics_a_mask_size_20 & dcache_atomics_a_mask_eq_97 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_6 ={ dcache_atomics_a_mask_acc_91 , dcache_atomics_a_mask_acc_90 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_6 ={ dcache_atomics_a_mask_acc_93 , dcache_atomics_a_mask_acc_92 }; 
    wire[3:0] dcache_atomics_a_mask_lo_6 ={ dcache_atomics_a_mask_lo_hi_6 , dcache_atomics_a_mask_lo_lo_6 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_6 ={ dcache_atomics_a_mask_acc_95 , dcache_atomics_a_mask_acc_94 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_6 ={ dcache_atomics_a_mask_acc_97 , dcache_atomics_a_mask_acc_96 }; 
    wire[3:0] dcache_atomics_a_mask_hi_6 ={ dcache_atomics_a_mask_hi_hi_6 , dcache_atomics_a_mask_hi_lo_6 }; 
    wire[7:0] dcache_atomics_a_6_mask ={ dcache_atomics_a_mask_hi_6 , dcache_atomics_a_mask_lo_6 }; 
    wire dcache_atomics_legal_7 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_7_opcode =3'h2; 
    wire[3:0] dcache_atomics_a_7_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_7_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_225 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_7 = dcache__GEN_225 [1:0]; 
    wire[3:0] dcache__GEN_226 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_7 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_7 = dcache__GEN_226 [2:0]|3'h1; 
    wire dcache__GEN_227 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_21 = dcache_atomics_a_mask_sizeOH_7 [2]; 
    wire dcache_atomics_a_mask_bit_21 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_21 = dcache_atomics_a_mask_bit_21 ==1'h0; 
    wire dcache_atomics_a_mask_eq_98 = dcache_atomics_a_mask_nbit_21 &1'h1; 
    wire dcache_atomics_a_mask_acc_98 = dcache__GEN_227 | dcache_atomics_a_mask_size_21 & dcache_atomics_a_mask_eq_98 ; 
    wire dcache_atomics_a_mask_eq_99 = dcache_atomics_a_mask_bit_21 &1'h1; 
    wire dcache_atomics_a_mask_acc_99 = dcache__GEN_227 | dcache_atomics_a_mask_size_21 & dcache_atomics_a_mask_eq_99 ; 
    wire dcache_atomics_a_mask_size_22 = dcache_atomics_a_mask_sizeOH_7 [1]; 
    wire dcache_atomics_a_mask_bit_22 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_22 = dcache_atomics_a_mask_bit_22 ==1'h0; 
    wire dcache_atomics_a_mask_eq_100 = dcache_atomics_a_mask_eq_98 & dcache_atomics_a_mask_nbit_22 ; 
    wire dcache_atomics_a_mask_acc_100 = dcache_atomics_a_mask_acc_98 | dcache_atomics_a_mask_size_22 & dcache_atomics_a_mask_eq_100 ; 
    wire dcache_atomics_a_mask_eq_101 = dcache_atomics_a_mask_eq_98 & dcache_atomics_a_mask_bit_22 ; 
    wire dcache_atomics_a_mask_acc_101 = dcache_atomics_a_mask_acc_98 | dcache_atomics_a_mask_size_22 & dcache_atomics_a_mask_eq_101 ; 
    wire dcache_atomics_a_mask_eq_102 = dcache_atomics_a_mask_eq_99 & dcache_atomics_a_mask_nbit_22 ; 
    wire dcache_atomics_a_mask_acc_102 = dcache_atomics_a_mask_acc_99 | dcache_atomics_a_mask_size_22 & dcache_atomics_a_mask_eq_102 ; 
    wire dcache_atomics_a_mask_eq_103 = dcache_atomics_a_mask_eq_99 & dcache_atomics_a_mask_bit_22 ; 
    wire dcache_atomics_a_mask_acc_103 = dcache_atomics_a_mask_acc_99 | dcache_atomics_a_mask_size_22 & dcache_atomics_a_mask_eq_103 ; 
    wire dcache_atomics_a_mask_size_23 = dcache_atomics_a_mask_sizeOH_7 [0]; 
    wire dcache_atomics_a_mask_bit_23 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_23 = dcache_atomics_a_mask_bit_23 ==1'h0; 
    wire dcache_atomics_a_mask_eq_104 = dcache_atomics_a_mask_eq_100 & dcache_atomics_a_mask_nbit_23 ; 
    wire dcache_atomics_a_mask_acc_104 = dcache_atomics_a_mask_acc_100 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_104 ; 
    wire dcache_atomics_a_mask_eq_105 = dcache_atomics_a_mask_eq_100 & dcache_atomics_a_mask_bit_23 ; 
    wire dcache_atomics_a_mask_acc_105 = dcache_atomics_a_mask_acc_100 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_105 ; 
    wire dcache_atomics_a_mask_eq_106 = dcache_atomics_a_mask_eq_101 & dcache_atomics_a_mask_nbit_23 ; 
    wire dcache_atomics_a_mask_acc_106 = dcache_atomics_a_mask_acc_101 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_106 ; 
    wire dcache_atomics_a_mask_eq_107 = dcache_atomics_a_mask_eq_101 & dcache_atomics_a_mask_bit_23 ; 
    wire dcache_atomics_a_mask_acc_107 = dcache_atomics_a_mask_acc_101 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_107 ; 
    wire dcache_atomics_a_mask_eq_108 = dcache_atomics_a_mask_eq_102 & dcache_atomics_a_mask_nbit_23 ; 
    wire dcache_atomics_a_mask_acc_108 = dcache_atomics_a_mask_acc_102 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_108 ; 
    wire dcache_atomics_a_mask_eq_109 = dcache_atomics_a_mask_eq_102 & dcache_atomics_a_mask_bit_23 ; 
    wire dcache_atomics_a_mask_acc_109 = dcache_atomics_a_mask_acc_102 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_109 ; 
    wire dcache_atomics_a_mask_eq_110 = dcache_atomics_a_mask_eq_103 & dcache_atomics_a_mask_nbit_23 ; 
    wire dcache_atomics_a_mask_acc_110 = dcache_atomics_a_mask_acc_103 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_110 ; 
    wire dcache_atomics_a_mask_eq_111 = dcache_atomics_a_mask_eq_103 & dcache_atomics_a_mask_bit_23 ; 
    wire dcache_atomics_a_mask_acc_111 = dcache_atomics_a_mask_acc_103 | dcache_atomics_a_mask_size_23 & dcache_atomics_a_mask_eq_111 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_7 ={ dcache_atomics_a_mask_acc_105 , dcache_atomics_a_mask_acc_104 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_7 ={ dcache_atomics_a_mask_acc_107 , dcache_atomics_a_mask_acc_106 }; 
    wire[3:0] dcache_atomics_a_mask_lo_7 ={ dcache_atomics_a_mask_lo_hi_7 , dcache_atomics_a_mask_lo_lo_7 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_7 ={ dcache_atomics_a_mask_acc_109 , dcache_atomics_a_mask_acc_108 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_7 ={ dcache_atomics_a_mask_acc_111 , dcache_atomics_a_mask_acc_110 }; 
    wire[3:0] dcache_atomics_a_mask_hi_7 ={ dcache_atomics_a_mask_hi_hi_7 , dcache_atomics_a_mask_hi_lo_7 }; 
    wire[7:0] dcache_atomics_a_7_mask ={ dcache_atomics_a_mask_hi_7 , dcache_atomics_a_mask_lo_7 }; 
    wire dcache_atomics_legal_8 =(2'h0<= dcache_s2_req_size & dcache_s2_req_size <=2'h3|1'h0)&(({1'h0, dcache_s2_req_addr }&35'hC8010000)==35'h0|({1'h0, dcache_s2_req_addr ^34'h8000000}&35'hC8000000)==35'h0)|1'h0; 
    wire[2:0] dcache_atomics_a_8_opcode =3'h2; 
    wire[3:0] dcache_atomics_a_8_size ={2'h0, dcache_s2_req_size }; 
    wire[31:0] dcache_atomics_a_8_address = dcache_s2_req_addr [31:0]; 
    wire[2:0] dcache__GEN_228 ={1'h0, dcache_s2_req_size }; 
    wire[1:0] dcache_atomics_a_mask_sizeOH_shiftAmount_8 = dcache__GEN_228 [1:0]; 
    wire[3:0] dcache__GEN_229 =4'h1<< dcache_atomics_a_mask_sizeOH_shiftAmount_8 ; 
    wire[2:0] dcache_atomics_a_mask_sizeOH_8 = dcache__GEN_229 [2:0]|3'h1; 
    wire dcache__GEN_230 = dcache_s2_req_size >=2'h3; 
    wire dcache_atomics_a_mask_size_24 = dcache_atomics_a_mask_sizeOH_8 [2]; 
    wire dcache_atomics_a_mask_bit_24 = dcache_s2_req_addr [2]; 
    wire dcache_atomics_a_mask_nbit_24 = dcache_atomics_a_mask_bit_24 ==1'h0; 
    wire dcache_atomics_a_mask_eq_112 = dcache_atomics_a_mask_nbit_24 &1'h1; 
    wire dcache_atomics_a_mask_acc_112 = dcache__GEN_230 | dcache_atomics_a_mask_size_24 & dcache_atomics_a_mask_eq_112 ; 
    wire dcache_atomics_a_mask_eq_113 = dcache_atomics_a_mask_bit_24 &1'h1; 
    wire dcache_atomics_a_mask_acc_113 = dcache__GEN_230 | dcache_atomics_a_mask_size_24 & dcache_atomics_a_mask_eq_113 ; 
    wire dcache_atomics_a_mask_size_25 = dcache_atomics_a_mask_sizeOH_8 [1]; 
    wire dcache_atomics_a_mask_bit_25 = dcache_s2_req_addr [1]; 
    wire dcache_atomics_a_mask_nbit_25 = dcache_atomics_a_mask_bit_25 ==1'h0; 
    wire dcache_atomics_a_mask_eq_114 = dcache_atomics_a_mask_eq_112 & dcache_atomics_a_mask_nbit_25 ; 
    wire dcache_atomics_a_mask_acc_114 = dcache_atomics_a_mask_acc_112 | dcache_atomics_a_mask_size_25 & dcache_atomics_a_mask_eq_114 ; 
    wire dcache_atomics_a_mask_eq_115 = dcache_atomics_a_mask_eq_112 & dcache_atomics_a_mask_bit_25 ; 
    wire dcache_atomics_a_mask_acc_115 = dcache_atomics_a_mask_acc_112 | dcache_atomics_a_mask_size_25 & dcache_atomics_a_mask_eq_115 ; 
    wire dcache_atomics_a_mask_eq_116 = dcache_atomics_a_mask_eq_113 & dcache_atomics_a_mask_nbit_25 ; 
    wire dcache_atomics_a_mask_acc_116 = dcache_atomics_a_mask_acc_113 | dcache_atomics_a_mask_size_25 & dcache_atomics_a_mask_eq_116 ; 
    wire dcache_atomics_a_mask_eq_117 = dcache_atomics_a_mask_eq_113 & dcache_atomics_a_mask_bit_25 ; 
    wire dcache_atomics_a_mask_acc_117 = dcache_atomics_a_mask_acc_113 | dcache_atomics_a_mask_size_25 & dcache_atomics_a_mask_eq_117 ; 
    wire dcache_atomics_a_mask_size_26 = dcache_atomics_a_mask_sizeOH_8 [0]; 
    wire dcache_atomics_a_mask_bit_26 = dcache_s2_req_addr [0]; 
    wire dcache_atomics_a_mask_nbit_26 = dcache_atomics_a_mask_bit_26 ==1'h0; 
    wire dcache_atomics_a_mask_eq_118 = dcache_atomics_a_mask_eq_114 & dcache_atomics_a_mask_nbit_26 ; 
    wire dcache_atomics_a_mask_acc_118 = dcache_atomics_a_mask_acc_114 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_118 ; 
    wire dcache_atomics_a_mask_eq_119 = dcache_atomics_a_mask_eq_114 & dcache_atomics_a_mask_bit_26 ; 
    wire dcache_atomics_a_mask_acc_119 = dcache_atomics_a_mask_acc_114 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_119 ; 
    wire dcache_atomics_a_mask_eq_120 = dcache_atomics_a_mask_eq_115 & dcache_atomics_a_mask_nbit_26 ; 
    wire dcache_atomics_a_mask_acc_120 = dcache_atomics_a_mask_acc_115 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_120 ; 
    wire dcache_atomics_a_mask_eq_121 = dcache_atomics_a_mask_eq_115 & dcache_atomics_a_mask_bit_26 ; 
    wire dcache_atomics_a_mask_acc_121 = dcache_atomics_a_mask_acc_115 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_121 ; 
    wire dcache_atomics_a_mask_eq_122 = dcache_atomics_a_mask_eq_116 & dcache_atomics_a_mask_nbit_26 ; 
    wire dcache_atomics_a_mask_acc_122 = dcache_atomics_a_mask_acc_116 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_122 ; 
    wire dcache_atomics_a_mask_eq_123 = dcache_atomics_a_mask_eq_116 & dcache_atomics_a_mask_bit_26 ; 
    wire dcache_atomics_a_mask_acc_123 = dcache_atomics_a_mask_acc_116 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_123 ; 
    wire dcache_atomics_a_mask_eq_124 = dcache_atomics_a_mask_eq_117 & dcache_atomics_a_mask_nbit_26 ; 
    wire dcache_atomics_a_mask_acc_124 = dcache_atomics_a_mask_acc_117 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_124 ; 
    wire dcache_atomics_a_mask_eq_125 = dcache_atomics_a_mask_eq_117 & dcache_atomics_a_mask_bit_26 ; 
    wire dcache_atomics_a_mask_acc_125 = dcache_atomics_a_mask_acc_117 | dcache_atomics_a_mask_size_26 & dcache_atomics_a_mask_eq_125 ; 
    wire[1:0] dcache_atomics_a_mask_lo_lo_8 ={ dcache_atomics_a_mask_acc_119 , dcache_atomics_a_mask_acc_118 }; 
    wire[1:0] dcache_atomics_a_mask_lo_hi_8 ={ dcache_atomics_a_mask_acc_121 , dcache_atomics_a_mask_acc_120 }; 
    wire[3:0] dcache_atomics_a_mask_lo_8 ={ dcache_atomics_a_mask_lo_hi_8 , dcache_atomics_a_mask_lo_lo_8 }; 
    wire[1:0] dcache_atomics_a_mask_hi_lo_8 ={ dcache_atomics_a_mask_acc_123 , dcache_atomics_a_mask_acc_122 }; 
    wire[1:0] dcache_atomics_a_mask_hi_hi_8 ={ dcache_atomics_a_mask_acc_125 , dcache_atomics_a_mask_acc_124 }; 
    wire[3:0] dcache_atomics_a_mask_hi_8 ={ dcache_atomics_a_mask_hi_hi_8 , dcache_atomics_a_mask_hi_lo_8 }; 
    wire[7:0] dcache_atomics_a_8_mask ={ dcache_atomics_a_mask_hi_8 , dcache_atomics_a_mask_lo_8 }; 
    wire dcache__GEN_231 =5'h4== dcache_s2_req_cmd ; 
    wire dcache__GEN_232 =5'h9== dcache_s2_req_cmd ; 
    wire dcache__GEN_233 =5'hA== dcache_s2_req_cmd ; 
    wire dcache__GEN_234 =5'hB== dcache_s2_req_cmd ; 
    wire dcache__GEN_235 =5'h8== dcache_s2_req_cmd ; 
    wire dcache__GEN_236 =5'hC== dcache_s2_req_cmd ; 
    wire dcache__GEN_237 =5'hD== dcache_s2_req_cmd ; 
    wire dcache__GEN_238 =5'hE== dcache_s2_req_cmd ; 
    wire dcache__GEN_239 =5'hF== dcache_s2_req_cmd ; 
    wire[2:0] dcache_atomics_opcode = dcache__GEN_239  ?  dcache_atomics_a_8_opcode : dcache__GEN_238  ?  dcache_atomics_a_7_opcode : dcache__GEN_237  ?  dcache_atomics_a_6_opcode : dcache__GEN_236  ?  dcache_atomics_a_5_opcode : dcache__GEN_235  ?  dcache_atomics_a_4_opcode : dcache__GEN_234  ?  dcache_atomics_a_3_opcode : dcache__GEN_233  ?  dcache_atomics_a_2_opcode : dcache__GEN_232  ?  dcache_atomics_a_1_opcode : dcache__GEN_231  ?  dcache_atomics_a_opcode : dcache__atomics_WIRE_1_opcode ; 
    wire[2:0] dcache_atomics_param = dcache__GEN_239  ?  dcache_atomics_a_8_param : dcache__GEN_238  ?  dcache_atomics_a_7_param : dcache__GEN_237  ?  dcache_atomics_a_6_param : dcache__GEN_236  ?  dcache_atomics_a_5_param : dcache__GEN_235  ?  dcache_atomics_a_4_param : dcache__GEN_234  ?  dcache_atomics_a_3_param : dcache__GEN_233  ?  dcache_atomics_a_2_param : dcache__GEN_232  ?  dcache_atomics_a_1_param : dcache__GEN_231  ?  dcache_atomics_a_param : dcache__atomics_WIRE_1_param ; 
    wire[3:0] dcache_atomics_size = dcache__GEN_239  ?  dcache_atomics_a_8_size : dcache__GEN_238  ?  dcache_atomics_a_7_size : dcache__GEN_237  ?  dcache_atomics_a_6_size : dcache__GEN_236  ?  dcache_atomics_a_5_size : dcache__GEN_235  ?  dcache_atomics_a_4_size : dcache__GEN_234  ?  dcache_atomics_a_3_size : dcache__GEN_233  ?  dcache_atomics_a_2_size : dcache__GEN_232  ?  dcache_atomics_a_1_size : dcache__GEN_231  ?  dcache_atomics_a_size : dcache__atomics_WIRE_1_size ; 
    wire dcache_atomics_source = dcache__GEN_239  ?  dcache_atomics_a_8_source : dcache__GEN_238  ?  dcache_atomics_a_7_source : dcache__GEN_237  ?  dcache_atomics_a_6_source : dcache__GEN_236  ?  dcache_atomics_a_5_source : dcache__GEN_235  ?  dcache_atomics_a_4_source : dcache__GEN_234  ?  dcache_atomics_a_3_source : dcache__GEN_233  ?  dcache_atomics_a_2_source : dcache__GEN_232  ?  dcache_atomics_a_1_source : dcache__GEN_231  ?  dcache_atomics_a_source : dcache__atomics_WIRE_1_source ; 
    wire[31:0] dcache_atomics_address = dcache__GEN_239  ?  dcache_atomics_a_8_address : dcache__GEN_238  ?  dcache_atomics_a_7_address : dcache__GEN_237  ?  dcache_atomics_a_6_address : dcache__GEN_236  ?  dcache_atomics_a_5_address : dcache__GEN_235  ?  dcache_atomics_a_4_address : dcache__GEN_234  ?  dcache_atomics_a_3_address : dcache__GEN_233  ?  dcache_atomics_a_2_address : dcache__GEN_232  ?  dcache_atomics_a_1_address : dcache__GEN_231  ?  dcache_atomics_a_address : dcache__atomics_WIRE_1_address ; 
    wire dcache_atomics_user_amba_prot_bufferable = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_bufferable : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_bufferable : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_bufferable : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_bufferable : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_bufferable : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_bufferable : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_bufferable : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_bufferable : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_bufferable : dcache__atomics_WIRE_1_user_amba_prot_bufferable ; 
    wire dcache_atomics_user_amba_prot_modifiable = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_modifiable : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_modifiable : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_modifiable : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_modifiable : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_modifiable : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_modifiable : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_modifiable : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_modifiable : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_modifiable : dcache__atomics_WIRE_1_user_amba_prot_modifiable ; 
    wire dcache_atomics_user_amba_prot_readalloc = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_readalloc : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_readalloc : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_readalloc : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_readalloc : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_readalloc : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_readalloc : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_readalloc : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_readalloc : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_readalloc : dcache__atomics_WIRE_1_user_amba_prot_readalloc ; 
    wire dcache_atomics_user_amba_prot_writealloc = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_writealloc : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_writealloc : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_writealloc : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_writealloc : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_writealloc : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_writealloc : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_writealloc : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_writealloc : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_writealloc : dcache__atomics_WIRE_1_user_amba_prot_writealloc ; 
    wire dcache_atomics_user_amba_prot_privileged = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_privileged : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_privileged : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_privileged : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_privileged : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_privileged : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_privileged : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_privileged : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_privileged : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_privileged : dcache__atomics_WIRE_1_user_amba_prot_privileged ; 
    wire dcache_atomics_user_amba_prot_secure = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_secure : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_secure : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_secure : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_secure : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_secure : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_secure : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_secure : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_secure : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_secure : dcache__atomics_WIRE_1_user_amba_prot_secure ; 
    wire dcache_atomics_user_amba_prot_fetch = dcache__GEN_239  ?  dcache_atomics_a_8_user_amba_prot_fetch : dcache__GEN_238  ?  dcache_atomics_a_7_user_amba_prot_fetch : dcache__GEN_237  ?  dcache_atomics_a_6_user_amba_prot_fetch : dcache__GEN_236  ?  dcache_atomics_a_5_user_amba_prot_fetch : dcache__GEN_235  ?  dcache_atomics_a_4_user_amba_prot_fetch : dcache__GEN_234  ?  dcache_atomics_a_3_user_amba_prot_fetch : dcache__GEN_233  ?  dcache_atomics_a_2_user_amba_prot_fetch : dcache__GEN_232  ?  dcache_atomics_a_1_user_amba_prot_fetch : dcache__GEN_231  ?  dcache_atomics_a_user_amba_prot_fetch : dcache__atomics_WIRE_1_user_amba_prot_fetch ; 
    wire[7:0] dcache_atomics_mask = dcache__GEN_239  ?  dcache_atomics_a_8_mask : dcache__GEN_238  ?  dcache_atomics_a_7_mask : dcache__GEN_237  ?  dcache_atomics_a_6_mask : dcache__GEN_236  ?  dcache_atomics_a_5_mask : dcache__GEN_235  ?  dcache_atomics_a_4_mask : dcache__GEN_234  ?  dcache_atomics_a_3_mask : dcache__GEN_233  ?  dcache_atomics_a_2_mask : dcache__GEN_232  ?  dcache_atomics_a_1_mask : dcache__GEN_231  ?  dcache_atomics_a_mask : dcache__atomics_WIRE_1_mask ; 
    wire[63:0] dcache_atomics_data = dcache__GEN_239  ?  dcache_atomics_a_8_data : dcache__GEN_238  ?  dcache_atomics_a_7_data : dcache__GEN_237  ?  dcache_atomics_a_6_data : dcache__GEN_236  ?  dcache_atomics_a_5_data : dcache__GEN_235  ?  dcache_atomics_a_4_data : dcache__GEN_234  ?  dcache_atomics_a_3_data : dcache__GEN_233  ?  dcache_atomics_a_2_data : dcache__GEN_232  ?  dcache_atomics_a_1_data : dcache__GEN_231  ?  dcache_atomics_a_data : dcache__atomics_WIRE_1_data ; 
    wire dcache_atomics_corrupt = dcache__GEN_239  ?  dcache_atomics_a_8_corrupt : dcache__GEN_238  ?  dcache_atomics_a_7_corrupt : dcache__GEN_237  ?  dcache_atomics_a_6_corrupt : dcache__GEN_236  ?  dcache_atomics_a_5_corrupt : dcache__GEN_235  ?  dcache_atomics_a_4_corrupt : dcache__GEN_234  ?  dcache_atomics_a_3_corrupt : dcache__GEN_233  ?  dcache_atomics_a_2_corrupt : dcache__GEN_232  ?  dcache_atomics_a_1_corrupt : dcache__GEN_231  ?  dcache_atomics_a_corrupt : dcache__atomics_WIRE_1_corrupt ; 
    wire[33:0] dcache__GEN_240 = dcache_s2_req_addr ^{2'h0, dcache_release_ack_addr }; 
  assign  dcache_tl_out_a_valid = dcache_io_cpu_s2_kill ==1'h0&( dcache_s2_valid_uncached_pending | dcache_s2_valid_cached_miss &( dcache_release_ack_wait & dcache__GEN_240 [20:6]==15'h0)==1'h0&( dcache_s2_victim_dirty ==1'h0|1'h0)); 
    wire dcache__GEN_241 = dcache_s2_uncached ==1'h0; 
    wire[33:0] dcache__GEN_242 ={ dcache_s2_req_addr [33:6],6'h0}; 
    wire dcache_tl_out_a_bits_legal =({1'h0, dcache__GEN_242 ^34'h80000000}&35'h80000000)==35'h0&1'h1|1'h0; 
    wire[2:0] dcache_tl_out_a_bits_a_param ={1'h0, dcache_s2_grow_param }; 
    wire[3:0] dcache_tl_out_a_bits_a_size =4'h6; 
    wire[31:0] dcache_tl_out_a_bits_a_address = dcache__GEN_242 [31:0]; 
    wire[3:0] dcache__GEN_243 =4'h1<< dcache_tl_out_a_bits_a_mask_sizeOH_shiftAmount ; 
    wire[2:0] dcache_tl_out_a_bits_a_mask_sizeOH = dcache__GEN_243 [2:0]|3'h1; 
    wire dcache_tl_out_a_bits_a_mask_size = dcache_tl_out_a_bits_a_mask_sizeOH [2]; 
    wire dcache_tl_out_a_bits_a_mask_bit = dcache__GEN_242 [2]; 
    wire dcache_tl_out_a_bits_a_mask_nbit = dcache_tl_out_a_bits_a_mask_bit ==1'h0; 
    wire dcache_tl_out_a_bits_a_mask_eq = dcache_tl_out_a_bits_a_mask_nbit &1'h1; 
    wire dcache_tl_out_a_bits_a_mask_eq_1 = dcache_tl_out_a_bits_a_mask_bit &1'h1; 
    wire dcache_tl_out_a_bits_a_mask_size_1 = dcache_tl_out_a_bits_a_mask_sizeOH [1]; 
    wire dcache_tl_out_a_bits_a_mask_bit_1 = dcache__GEN_242 [1]; 
    wire dcache_tl_out_a_bits_a_mask_nbit_1 = dcache_tl_out_a_bits_a_mask_bit_1 ==1'h0; 
    wire dcache_tl_out_a_bits_a_mask_eq_2 = dcache_tl_out_a_bits_a_mask_eq & dcache_tl_out_a_bits_a_mask_nbit_1 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_2 = dcache_tl_out_a_bits_a_mask_acc | dcache_tl_out_a_bits_a_mask_size_1 & dcache_tl_out_a_bits_a_mask_eq_2 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_3 = dcache_tl_out_a_bits_a_mask_eq & dcache_tl_out_a_bits_a_mask_bit_1 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_3 = dcache_tl_out_a_bits_a_mask_acc | dcache_tl_out_a_bits_a_mask_size_1 & dcache_tl_out_a_bits_a_mask_eq_3 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_4 = dcache_tl_out_a_bits_a_mask_eq_1 & dcache_tl_out_a_bits_a_mask_nbit_1 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_4 = dcache_tl_out_a_bits_a_mask_acc_1 | dcache_tl_out_a_bits_a_mask_size_1 & dcache_tl_out_a_bits_a_mask_eq_4 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_5 = dcache_tl_out_a_bits_a_mask_eq_1 & dcache_tl_out_a_bits_a_mask_bit_1 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_5 = dcache_tl_out_a_bits_a_mask_acc_1 | dcache_tl_out_a_bits_a_mask_size_1 & dcache_tl_out_a_bits_a_mask_eq_5 ; 
    wire dcache_tl_out_a_bits_a_mask_size_2 = dcache_tl_out_a_bits_a_mask_sizeOH [0]; 
    wire dcache_tl_out_a_bits_a_mask_bit_2 = dcache__GEN_242 [0]; 
    wire dcache_tl_out_a_bits_a_mask_nbit_2 = dcache_tl_out_a_bits_a_mask_bit_2 ==1'h0; 
    wire dcache_tl_out_a_bits_a_mask_eq_6 = dcache_tl_out_a_bits_a_mask_eq_2 & dcache_tl_out_a_bits_a_mask_nbit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_6 = dcache_tl_out_a_bits_a_mask_acc_2 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_6 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_7 = dcache_tl_out_a_bits_a_mask_eq_2 & dcache_tl_out_a_bits_a_mask_bit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_7 = dcache_tl_out_a_bits_a_mask_acc_2 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_7 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_8 = dcache_tl_out_a_bits_a_mask_eq_3 & dcache_tl_out_a_bits_a_mask_nbit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_8 = dcache_tl_out_a_bits_a_mask_acc_3 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_8 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_9 = dcache_tl_out_a_bits_a_mask_eq_3 & dcache_tl_out_a_bits_a_mask_bit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_9 = dcache_tl_out_a_bits_a_mask_acc_3 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_9 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_10 = dcache_tl_out_a_bits_a_mask_eq_4 & dcache_tl_out_a_bits_a_mask_nbit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_10 = dcache_tl_out_a_bits_a_mask_acc_4 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_10 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_11 = dcache_tl_out_a_bits_a_mask_eq_4 & dcache_tl_out_a_bits_a_mask_bit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_11 = dcache_tl_out_a_bits_a_mask_acc_4 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_11 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_12 = dcache_tl_out_a_bits_a_mask_eq_5 & dcache_tl_out_a_bits_a_mask_nbit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_12 = dcache_tl_out_a_bits_a_mask_acc_5 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_12 ; 
    wire dcache_tl_out_a_bits_a_mask_eq_13 = dcache_tl_out_a_bits_a_mask_eq_5 & dcache_tl_out_a_bits_a_mask_bit_2 ; 
    wire dcache_tl_out_a_bits_a_mask_acc_13 = dcache_tl_out_a_bits_a_mask_acc_5 | dcache_tl_out_a_bits_a_mask_size_2 & dcache_tl_out_a_bits_a_mask_eq_13 ; 
    wire[1:0] dcache_tl_out_a_bits_a_mask_lo_lo ={ dcache_tl_out_a_bits_a_mask_acc_7 , dcache_tl_out_a_bits_a_mask_acc_6 }; 
    wire[1:0] dcache_tl_out_a_bits_a_mask_lo_hi ={ dcache_tl_out_a_bits_a_mask_acc_9 , dcache_tl_out_a_bits_a_mask_acc_8 }; 
    wire[3:0] dcache_tl_out_a_bits_a_mask_lo ={ dcache_tl_out_a_bits_a_mask_lo_hi , dcache_tl_out_a_bits_a_mask_lo_lo }; 
    wire[1:0] dcache_tl_out_a_bits_a_mask_hi_lo ={ dcache_tl_out_a_bits_a_mask_acc_11 , dcache_tl_out_a_bits_a_mask_acc_10 }; 
    wire[1:0] dcache_tl_out_a_bits_a_mask_hi_hi ={ dcache_tl_out_a_bits_a_mask_acc_13 , dcache_tl_out_a_bits_a_mask_acc_12 }; 
    wire[3:0] dcache_tl_out_a_bits_a_mask_hi ={ dcache_tl_out_a_bits_a_mask_hi_hi , dcache_tl_out_a_bits_a_mask_hi_lo }; 
    wire[7:0] dcache_tl_out_a_bits_a_mask ={ dcache_tl_out_a_bits_a_mask_hi , dcache_tl_out_a_bits_a_mask_lo }; 
    wire[63:0] dcache_tl_out_a_bits_a_data =64'h0; 
    wire dcache__GEN_244 = dcache_s2_write ==1'h0; 
    wire dcache__GEN_245 = dcache_s2_req_cmd ==5'h11; 
    wire dcache__GEN_246 = dcache_s2_read ==1'h0; 
  assign  dcache_tl_out_a_bits_opcode = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_opcode : dcache__GEN_244  ?  dcache_get_opcode : dcache__GEN_245  ?  dcache_putpartial_opcode : dcache__GEN_246  ?  dcache_put_opcode : dcache_atomics_opcode ; 
  assign  dcache_tl_out_a_bits_param = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_param : dcache__GEN_244  ?  dcache_get_param : dcache__GEN_245  ?  dcache_putpartial_param : dcache__GEN_246  ?  dcache_put_param : dcache_atomics_param ; 
  assign  dcache_tl_out_a_bits_size = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_size : dcache__GEN_244  ?  dcache_get_size : dcache__GEN_245  ?  dcache_putpartial_size : dcache__GEN_246  ?  dcache_put_size : dcache_atomics_size ; 
  assign  dcache_tl_out_a_bits_source = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_source : dcache__GEN_244  ?  dcache_get_source : dcache__GEN_245  ?  dcache_putpartial_source : dcache__GEN_246  ?  dcache_put_source : dcache_atomics_source ; 
  assign  dcache_tl_out_a_bits_address = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_address : dcache__GEN_244  ?  dcache_get_address : dcache__GEN_245  ?  dcache_putpartial_address : dcache__GEN_246  ?  dcache_put_address : dcache_atomics_address ; 
  assign  dcache_tl_out_a_bits_mask = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_mask : dcache__GEN_244  ?  dcache_get_mask : dcache__GEN_245  ?  dcache_putpartial_mask : dcache__GEN_246  ?  dcache_put_mask : dcache_atomics_mask ; 
  assign  dcache_tl_out_a_bits_data = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_data : dcache__GEN_244  ?  dcache_get_data : dcache__GEN_245  ?  dcache_putpartial_data : dcache__GEN_246  ?  dcache_put_data : dcache_atomics_data ; 
  assign  dcache_tl_out_a_bits_corrupt = dcache__GEN_241  ?  dcache_tl_out_a_bits_a_corrupt : dcache__GEN_244  ?  dcache_get_corrupt : dcache__GEN_245  ?  dcache_putpartial_corrupt : dcache__GEN_246  ?  dcache_put_corrupt : dcache_atomics_corrupt ; 
  assign  dcache_tl_out_a_bits_user_amba_prot_privileged =(& dcache_s2_req_dprv )| dcache_s2_pma_cacheable ; 
    wire[1:0] dcache__GEN_247 =2'h1<< dcache_a_sel_shiftAmount ; 
    wire dcache_a_sel = dcache__GEN_247 [1]; 
    wire dcache__GEN_248 = dcache_tl_out_a_ready & dcache_tl_out_a_valid ; 
    wire dcache__GEN_249 = dcache__GEN_248  ? ( dcache_s2_uncached  ? ( dcache_a_sel  ? 1'h1: dcache_uncachedInFlight_0 ): dcache_uncachedInFlight_0 ): dcache_uncachedInFlight_0 ; 
    wire[4:0] dcache__GEN_250 = dcache_s2_write  ? ( dcache_s2_req_cmd ==5'h11 ? 5'h11:5'h1):5'h0; 
    wire dcache__GEN_251 = dcache__GEN_248  ? ( dcache_s2_uncached  ?  dcache_cached_grant_wait :1'h1): dcache_cached_grant_wait ; 
    wire dcache_nodeOut_d_ready ; 
    wire dcache__GEN_252 = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid ; 
    wire[26:0] dcache__GEN_253 =27'hFFF<< dcache_nodeOut_d_bits_size ; 
    wire[11:0] dcache__GEN_254 =~( dcache__GEN_253 [11:0]); 
    wire[8:0] dcache_beats1_decode = dcache__GEN_254 [11:3]; 
    wire dcache_beats1_opdata = dcache_nodeOut_d_bits_opcode [0]; 
    wire[8:0] dcache_beats1 = dcache_beats1_opdata  ?  dcache_beats1_decode :9'h0; reg[8:0] dcache_counter ; 
    wire[9:0] dcache__GEN_255 ={1'h0, dcache_counter }-10'h1; 
    wire[8:0] dcache_counter1 = dcache__GEN_255 [8:0]; 
    wire dcache_d_first = dcache_counter ==9'h0; 
    wire dcache_d_last = dcache_counter ==9'h1| dcache_beats1 ==9'h0; 
    wire dcache_d_done = dcache_d_last & dcache__GEN_252 ; 
    wire[8:0] dcache_count = dcache_beats1 &~ dcache_counter1 ; 
    wire[11:0] dcache_d_address_inc ={ dcache_count ,3'h0}; 
    wire dcache_grantIsUncached = dcache_nodeOut_d_bits_opcode ==3'h1| dcache_nodeOut_d_bits_opcode ==3'h0| dcache_nodeOut_d_bits_opcode ==3'h2; 
    wire dcache_grantIsUncachedData = dcache_nodeOut_d_bits_opcode ==3'h1; 
    wire[15:0] dcache_tl_d_data_encoded_lo_lo_1 ={ dcache_nodeOut_d_bits_data [15:8], dcache_nodeOut_d_bits_data [7:0]}; 
    wire[15:0] dcache_tl_d_data_encoded_lo_hi_1 ={ dcache_nodeOut_d_bits_data [31:24], dcache_nodeOut_d_bits_data [23:16]}; 
    wire[31:0] dcache_tl_d_data_encoded_lo_1 ={ dcache_tl_d_data_encoded_lo_hi_1 , dcache_tl_d_data_encoded_lo_lo_1 }; 
    wire[15:0] dcache_tl_d_data_encoded_hi_lo_1 ={ dcache_nodeOut_d_bits_data [47:40], dcache_nodeOut_d_bits_data [39:32]}; 
    wire[15:0] dcache_tl_d_data_encoded_hi_hi_1 ={ dcache_nodeOut_d_bits_data [63:56], dcache_nodeOut_d_bits_data [55:48]}; 
    wire[31:0] dcache_tl_d_data_encoded_hi_1 ={ dcache_tl_d_data_encoded_hi_hi_1 , dcache_tl_d_data_encoded_hi_lo_1 }; 
  assign  dcache_tl_d_data_encoded ={ dcache_tl_d_data_encoded_hi_1 , dcache_tl_d_data_encoded_lo_1 }; 
    wire dcache_grantIsCached = dcache_nodeOut_d_bits_opcode ==3'h4| dcache_nodeOut_d_bits_opcode ==3'h5; 
    wire dcache_grantIsVoluntary = dcache_nodeOut_d_bits_opcode ==3'h6; 
    wire dcache_grantIsRefill = dcache_nodeOut_d_bits_opcode ==3'h5; 
    reg dcache_grantInProgress ; reg[2:0] dcache_blockProbeAfterGrantCount ; 
    wire dcache__GEN_256 = dcache_blockProbeAfterGrantCount >3'h0; 
    wire[3:0] dcache__GEN_257 ={1'h0, dcache_blockProbeAfterGrantCount }-4'h1; 
    wire[2:0] dcache__GEN_258 = dcache__GEN_256  ?  dcache__GEN_257 [2:0]: dcache_blockProbeAfterGrantCount ; 
    wire dcache_canAcceptCachedGrant =( dcache_release_state ==4'h1| dcache_release_state ==4'h6| dcache_release_state ==4'h9)==1'h0; 
    wire[1:0] dcache__GEN_259 =2'h1<< dcache_uncachedRespIdxOH_shiftAmount ; 
    wire dcache_uncachedRespIdxOH = dcache__GEN_259 [1]; 
    wire dcache__GEN_260 = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid ; 
    wire dcache__GEN_261 = dcache__GEN_260 & dcache_grantIsCached ; 
    wire dcache__GEN_262 = dcache_cached_grant_wait ==1'h0; 
    wire dcache__GEN_263 = dcache_d_last  ? 1'h0:1'h1; 
  assign  dcache_replace = dcache__GEN_260  ? ( dcache_grantIsCached  ?  dcache_d_last :1'h0):1'h0; 
    wire dcache__GEN_264 = dcache__GEN_260 &~ dcache_grantIsCached ; 
    wire dcache__GEN_265 = dcache__GEN_264 & dcache_grantIsUncached ; 
    wire dcache__GEN_266 = dcache_uncachedRespIdxOH & dcache_d_last ; 
    wire dcache__GEN_267 = dcache_uncachedInFlight_0 ==1'h0; 
  assign  dcache_s1_data_way = dcache__GEN_260  ? ( dcache_grantIsCached  ? 2'h1: dcache_grantIsUncached  ? ( dcache_grantIsUncachedData  ? 2'h2:2'h1):2'h1):2'h1; 
    wire[31:0] dcache_s2_req_addr_dontCareBits ={ dcache_s1_paddr [31:3],3'h0}; 
    wire[33:0] dcache__GEN_268 ={2'h0, dcache_s2_req_addr_dontCareBits |{29'h0, dcache_uncachedResp_addr [2:0]}}; 
    wire dcache__GEN_269 = dcache_release_ack_wait ==1'h0; 
    wire dcache__GEN_270 = dcache__GEN_260  ? ( dcache_grantIsCached  ?  dcache_release_ack_wait : dcache_grantIsUncached  ?  dcache_release_ack_wait : dcache_grantIsVoluntary  ? 1'h0: dcache_release_ack_wait ): dcache_release_ack_wait ; 
    wire dcache_nodeOut_e_valid ; 
    wire[1:0] dcache_nodeOut_e_bits_sink = dcache_nodeOut_e_bits_e_sink ; 
    wire dcache__GEN_271 =( dcache_nodeOut_e_ready & dcache_nodeOut_e_valid )==( dcache_nodeOut_d_ready & dcache_nodeOut_d_valid & dcache_d_first & dcache_grantIsCached )==1'h0; 
    wire dcache__GEN_272 = dcache_nodeOut_d_valid & dcache_grantIsRefill & dcache_canAcceptCachedGrant ; 
    wire dcache__GEN_273 = dcache_grantIsRefill & dcache_dataArb_io_in_1_ready ==1'h0; 
  assign  dcache_nodeOut_e_valid = dcache__GEN_273  ? 1'h0: dcache_nodeOut_d_valid & dcache_d_first & dcache_grantIsCached & dcache_canAcceptCachedGrant ; 
    wire[33:0] dcache__GEN_274 ={ dcache_s2_vaddr [33:6],6'h0}|{22'h0, dcache_d_address_inc }; 
  assign  dcache_dataArb_io_in_1_bits_addr = dcache__GEN_274 [11:0]; 
  assign  dcache_dataArb_io_in_1_bits_way_en = dcache_refill_way [0]; 
  assign  dcache_metaArb_io_in_3_valid = dcache_grantIsCached & dcache_d_done & dcache_nodeOut_d_bits_denied ==1'h0; 
  assign  dcache_metaArb_io_in_3_bits_way_en = dcache_refill_way [0]; 
  assign  dcache_metaArb_io_in_3_bits_idx = dcache_s2_vaddr [11:6]; 
  assign  dcache_metaArb_io_in_3_bits_addr ={ dcache_io_cpu_req_bits_addr [33:12], dcache_s2_vaddr [11:0]}; 
    wire[21:0] dcache__s2_req_addr_33to12_0 = dcache_s2_req_addr [33:12]; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_c ={ dcache_s2_req_cmd ==5'h1| dcache_s2_req_cmd ==5'h11| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF, dcache_s2_req_cmd ==5'h1| dcache_s2_req_cmd ==5'h11| dcache_s2_req_cmd ==5'h7| dcache_s2_req_cmd ==5'h4| dcache_s2_req_cmd ==5'h9| dcache_s2_req_cmd ==5'hA| dcache_s2_req_cmd ==5'hB| dcache_s2_req_cmd ==5'h8| dcache_s2_req_cmd ==5'hC| dcache_s2_req_cmd ==5'hD| dcache_s2_req_cmd ==5'hE| dcache_s2_req_cmd ==5'hF| dcache_s2_req_cmd ==5'h3| dcache_s2_req_cmd ==5'h6}; 
    wire[3:0] dcache__GEN_275 ={ dcache_metaArb_io_in_3_bits_data_c , dcache_nodeOut_d_bits_param }; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_meta_state =4'hC== dcache__GEN_275  ? 2'h3:4'h4== dcache__GEN_275  ? 2'h2:4'h0== dcache__GEN_275  ? 2'h2:4'h1== dcache__GEN_275  ? 2'h1:2'h0; 
    wire[1:0] dcache_metaArb_io_in_3_bits_data_meta_1_coh_state = dcache_metaArb_io_in_3_bits_data_meta_state ; 
    wire[19:0] dcache_metaArb_io_in_3_bits_data_meta_1_tag = dcache__s2_req_addr_33to12_0 [19:0]; 
  assign  dcache_metaArb_io_in_3_bits_data ={ dcache_metaArb_io_in_3_bits_data_meta_1_coh_state , dcache_metaArb_io_in_3_bits_data_meta_1_tag }; 
    reg dcache_blockUncachedGrant ; 
    wire dcache__GEN_276 = dcache_grantIsUncachedData &( dcache_blockUncachedGrant | dcache_s1_valid ); 
  assign  dcache_nodeOut_d_ready = dcache__GEN_276  ? 1'h0: dcache__GEN_273  ? 1'h0: dcache_grantIsCached  ? ( dcache_d_first ==1'h0| dcache_nodeOut_e_ready )& dcache_canAcceptCachedGrant :1'h1; 
  assign  dcache__io_cpu_req_ready_output = dcache__GEN_276  ? ( dcache_nodeOut_d_valid  ? 1'h0: dcache__GEN_94 ): dcache__GEN_94 ; 
  assign  dcache_dataArb_io_in_1_valid = dcache__GEN_276  ? ( dcache_nodeOut_d_valid  ? 1'h1: dcache__GEN_272 ): dcache__GEN_272 ; 
  assign  dcache_dataArb_io_in_1_bits_write = dcache__GEN_276  ? ( dcache_nodeOut_d_valid  ? 1'h0:1'h1):1'h1; 
    wire dcache__GEN_277 = dcache_dataArb_io_in_1_ready ==1'h0; 
    wire dcache_block_probe_for_core_progress = dcache_blockProbeAfterGrantCount >3'h0| dcache_lrscValid ; 
    wire[31:0] dcache__GEN_278 = dcache_nodeOut_b_bits_address ^ dcache_release_ack_addr ; 
    wire dcache_block_probe_for_pending_release_ack = dcache_release_ack_wait & dcache__GEN_278 [20:6]==15'h0; 
    wire dcache_block_probe_for_ordering = dcache_releaseInFlight | dcache_block_probe_for_pending_release_ack | dcache_grantInProgress ; 
  assign  dcache_nodeOut_b_ready = dcache_metaArb_io_in_6_ready &( dcache_block_probe_for_core_progress | dcache_block_probe_for_ordering | dcache_s1_valid | dcache_s2_valid )==1'h0; 
    wire dcache_nodeOut_c_valid ; 
    wire dcache__GEN_279 = dcache_nodeOut_c_ready & dcache_nodeOut_c_valid ; 
    wire[3:0] dcache_nodeOut_c_bits_size ; 
    wire[26:0] dcache__GEN_280 =27'hFFF<< dcache_nodeOut_c_bits_size ; 
    wire[11:0] dcache__GEN_281 =~( dcache__GEN_280 [11:0]); 
    wire[8:0] dcache_beats1_decode_1 = dcache__GEN_281 [11:3]; 
    wire[2:0] dcache_nodeOut_c_bits_opcode ; 
    wire dcache_beats1_opdata_1 = dcache_nodeOut_c_bits_opcode [0]; 
    wire[8:0] dcache_beats1_1 = dcache_beats1_opdata_1  ?  dcache_beats1_decode_1 :9'h0; reg[8:0] dcache_counter_1 ; 
    wire[9:0] dcache__GEN_282 ={1'h0, dcache_counter_1 }-10'h1; 
    wire[8:0] dcache_counter1_1 = dcache__GEN_282 [8:0]; 
    wire dcache_c_first = dcache_counter_1 ==9'h0; 
    wire dcache_c_last = dcache_counter_1 ==9'h1| dcache_beats1_1 ==9'h0; 
    wire dcache_releaseDone = dcache_c_last & dcache__GEN_279 ; 
    wire[8:0] dcache_c_count = dcache_beats1_1 &~ dcache_counter1_1 ; 
    reg dcache_s1_release_data_valid ; 
    wire dcache_releaseRejected ; 
    reg dcache_s2_release_data_valid ; 
  assign  dcache_releaseRejected = dcache_s2_release_data_valid &( dcache_nodeOut_c_ready & dcache_nodeOut_c_valid )==1'h0; 
    wire[2:0] dcache__GEN_283 ={2'h0, dcache_s1_release_data_valid }+{1'h0,{1'h0, dcache_s2_release_data_valid }}; 
    wire[10:0] dcache__GEN_284 ={1'h0,{1'h0, dcache_c_count }}+{9'h0, dcache_releaseRejected  ? 2'h0: dcache__GEN_283 [1:0]}; 
    wire[9:0] dcache_releaseDataBeat = dcache__GEN_284 [9:0]; 
    wire[63:0] dcache_nackResponseMessage_data =64'h0; 
    wire[63:0] dcache_cleanReleaseMessage_data =64'h0; 
    wire[63:0] dcache_dirtyReleaseMessage_data =64'h0; 
    wire dcache__GEN_285 = dcache_s2_release_data_valid &( dcache_c_first & dcache_release_ack_wait )==1'h0; 
    wire[1:0] dcache_metaArb_io_in_4_bits_data_meta_coh_state = dcache_newCoh_state ; 
    wire dcache__GEN_286 =( dcache_s2_valid_flush_line | dcache_s2_flush_valid | dcache__io_cpu_s2_nack_output )==1'h0; 
    wire dcache_discard_line = dcache_s2_valid_flush_line & dcache_s2_req_size [1]| dcache_s2_flush_valid & dcache_flushing_req_size [1]; 
    wire[3:0] dcache__GEN_287 = dcache_s2_victim_dirty & dcache_discard_line ==1'h0 ? 4'h1:4'h6; 
    wire[31:0] dcache_probe_bits_res_address ={{ dcache_s2_victim_tag , dcache_s2_req_addr [11:6]},6'h0}; 
    wire dcache__GEN_288 = dcache_s2_probe &~ dcache_s2_meta_error ; 
    wire dcache__GEN_289 = dcache__GEN_288 &~ dcache_s2_prb_ack_data ; 
    wire dcache__GEN_290 = dcache_s2_probe_state_state >2'h0; 
    wire dcache_probeNack = dcache_s2_meta_error  ? 1'h1: dcache_s2_prb_ack_data  ? 1'h1: dcache__GEN_290  ? 1'h1: dcache_releaseDone ==1'h0; 
    wire[3:0] dcache__GEN_291 = dcache_s2_probe  ? ( dcache_s2_meta_error  ? 4'h4: dcache_s2_prb_ack_data  ? 4'h2: dcache__GEN_290  ? ( dcache_releaseDone  ? 4'h7:4'h3): dcache_releaseDone  ? 4'h0:4'h5): dcache_s2_victimize  ?  dcache__GEN_287 : dcache_release_state ; 
  assign  dcache_s1_nack = dcache_s2_probe  ? ( dcache_probeNack  ? 1'h1: dcache__GEN_196 ): dcache__GEN_196 ; 
    wire dcache__GEN_292 = dcache_release_state ==4'h4; 
  assign  dcache_metaArb_io_in_6_valid = dcache__GEN_292  ? 1'h1: dcache_nodeOut_b_valid &( dcache_block_probe_for_core_progress ==1'h0| dcache_lrscBackingOff ); 
  assign  dcache_metaArb_io_in_6_bits_idx = dcache__GEN_292  ?  dcache_probe_bits_address [11:6]: dcache_nodeOut_b_bits_address [11:6]; 
  assign  dcache_metaArb_io_in_6_bits_addr = dcache__GEN_292  ? { dcache_io_cpu_req_bits_addr [33:32], dcache_probe_bits_address }:{ dcache_io_cpu_req_bits_addr [33:32], dcache_nodeOut_b_bits_address }; 
    wire[3:0] dcache__GEN_293 = dcache__GEN_292  ? ( dcache_metaArb_io_in_6_ready  ? 4'h0: dcache__GEN_291 ): dcache__GEN_291 ; 
    wire dcache__GEN_294 = dcache_release_state ==4'h5; 
    wire[3:0] dcache__GEN_295 = dcache__GEN_294  ? ( dcache_releaseDone  ? 4'h0: dcache__GEN_293 ): dcache__GEN_293 ; 
    wire dcache__GEN_296 = dcache_release_state ==4'h3; 
  assign  dcache_nodeOut_c_valid = dcache__GEN_296  ? 1'h1: dcache__GEN_294  ? 1'h1: dcache_s2_probe  ? ( dcache_s2_meta_error  ?  dcache__GEN_285 : dcache_s2_prb_ack_data  ?  dcache__GEN_285 :1'h1): dcache__GEN_285 ; 
    wire[3:0] dcache__GEN_297 = dcache__GEN_296  ? ( dcache_releaseDone  ? 4'h7: dcache__GEN_295 ): dcache__GEN_295 ; 
    wire dcache__GEN_298 = dcache_release_state ==4'h2; 
    wire[3:0] dcache__GEN_299 = dcache__GEN_298  ? ( dcache_releaseDone  ? 4'h7: dcache__GEN_297 ): dcache__GEN_297 ; 
    wire dcache__GEN_300 = dcache_release_state ==4'h1| dcache_release_state ==4'h6| dcache_release_state ==4'h9; 
    wire dcache__GEN_301 = dcache_release_state ==4'h9; 
    wire[3:0] dcache_nodeOut_c_bits_c_size =4'h6; 
    wire[31:0] dcache_nodeOut_c_bits_c_address =32'h0; 
    wire[63:0] dcache_nodeOut_c_bits_c_data =64'h0; 
    wire[3:0] dcache_nodeOut_c_bits_c_1_size =4'h6; 
    wire[31:0] dcache_nodeOut_c_bits_c_1_address =32'h0; 
    wire[63:0] dcache_nodeOut_c_bits_c_1_data =64'h0; 
  assign  dcache_nodeOut_c_bits_opcode = dcache__GEN_300  ? ( dcache__GEN_301  ?  dcache_nodeOut_c_bits_c_opcode : dcache_nodeOut_c_bits_c_1_opcode ): dcache__GEN_298  ?  dcache_dirtyReleaseMessage_opcode : dcache__GEN_296  ?  dcache_cleanReleaseMessage_opcode : dcache_s2_probe  ? ( dcache_s2_meta_error  ?  dcache_nackResponseMessage_opcode : dcache_s2_prb_ack_data  ?  dcache_nackResponseMessage_opcode : dcache__GEN_290  ?  dcache_cleanReleaseMessage_opcode : dcache_nackResponseMessage_opcode ): dcache_nackResponseMessage_opcode ; 
    wire[2:0] dcache_nodeOut_c_bits_param = dcache__GEN_300  ? ( dcache__GEN_301  ?  dcache_nodeOut_c_bits_c_param : dcache_nodeOut_c_bits_c_1_param ): dcache__GEN_298  ?  dcache_dirtyReleaseMessage_param : dcache__GEN_296  ?  dcache_cleanReleaseMessage_param : dcache_s2_probe  ? ( dcache_s2_meta_error  ?  dcache_nackResponseMessage_param : dcache_s2_prb_ack_data  ?  dcache_nackResponseMessage_param : dcache__GEN_290  ?  dcache_cleanReleaseMessage_param : dcache_nackResponseMessage_param ): dcache_nackResponseMessage_param ; 
  assign  dcache_nodeOut_c_bits_size = dcache__GEN_300  ? ( dcache__GEN_301  ?  dcache_nodeOut_c_bits_c_size : dcache_nodeOut_c_bits_c_1_size ): dcache__GEN_298  ?  dcache_dirtyReleaseMessage_size : dcache__GEN_296  ?  dcache_cleanReleaseMessage_size : dcache_s2_probe  ? ( dcache_s2_meta_error  ?  dcache_nackResponseMessage_size : dcache_s2_prb_ack_data  ?  dcache_nackResponseMessage_size : dcache__GEN_290  ?  dcache_cleanReleaseMessage_size : dcache_nackResponseMessage_size ): dcache_nackResponseMessage_size ; 
  assign  dcache_newCoh_state = dcache__GEN_300  ?  dcache_voluntaryNewCoh_state : dcache_probeNewCoh_state ; 
    wire[1:0] dcache_releaseWay = dcache__GEN_300  ?  dcache_s2_victim_or_hit_way :{1'h0, dcache_s2_probe_way }; 
    wire dcache__GEN_302 = dcache_nodeOut_c_ready & dcache_nodeOut_c_valid & dcache_c_first ; 
    wire dcache_nodeOut_c_bits_corrupt = dcache_inWriteback & dcache_s2_data_error_uncorrectable ; 
  assign  dcache_dataArb_io_in_2_valid = dcache_inWriteback & dcache_releaseDataBeat <10'h8; 
  assign  dcache_dataArb_io_in_2_bits_addr ={ dcache_probe_bits_address [11:6],6'h0}|{6'h0,{ dcache_releaseDataBeat [2:0],3'h0}}; 
  assign  dcache_metaArb_io_in_4_valid = dcache_release_state ==4'h6| dcache_release_state ==4'h7; 
  assign  dcache_metaArb_io_in_4_bits_way_en = dcache_releaseWay [0]; 
  assign  dcache_metaArb_io_in_4_bits_idx = dcache_probe_bits_address [11:6]; 
  assign  dcache_metaArb_io_in_4_bits_addr ={ dcache_io_cpu_req_bits_addr [33:12], dcache_probe_bits_address [11:0]}; 
    wire[19:0] dcache_metaArb_io_in_4_bits_data_meta_tag = dcache_nodeOut_c_bits_address [31:12]; 
  assign  dcache_metaArb_io_in_4_bits_data ={ dcache_metaArb_io_in_4_bits_data_meta_coh_state , dcache_metaArb_io_in_4_bits_data_meta_tag }; 
    wire dcache__GEN_303 = dcache_metaArb_io_in_4_ready & dcache_metaArb_io_in_4_valid ; 
    wire dcache_s1_xcpt_valid = dcache_tlb_io_req_valid & dcache_s1_req_no_xcpt ==1'h0& dcache_s1_nack ==1'h0; 
    reg dcache_io_cpu_s2_xcpt_REG ; 
  assign  dcache__io_cpu_s2_xcpt_pf_ld_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_pf_ld : dcache__io_cpu_s2_xcpt_WIRE_pf_ld ; 
  assign  dcache__io_cpu_s2_xcpt_pf_st_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_pf_st : dcache__io_cpu_s2_xcpt_WIRE_pf_st ; 
  assign  dcache__io_cpu_s2_xcpt_gf_ld_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_gf_ld : dcache__io_cpu_s2_xcpt_WIRE_gf_ld ; 
  assign  dcache__io_cpu_s2_xcpt_gf_st_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_gf_st : dcache__io_cpu_s2_xcpt_WIRE_gf_st ; 
  assign  dcache__io_cpu_s2_xcpt_ae_ld_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_ae_ld : dcache__io_cpu_s2_xcpt_WIRE_ae_ld ; 
  assign  dcache__io_cpu_s2_xcpt_ae_st_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_ae_st : dcache__io_cpu_s2_xcpt_WIRE_ae_st ; 
  assign  dcache__io_cpu_s2_xcpt_ma_ld_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_ma_ld : dcache__io_cpu_s2_xcpt_WIRE_ma_ld ; 
  assign  dcache__io_cpu_s2_xcpt_ma_st_output = dcache_io_cpu_s2_xcpt_REG  ?  dcache_s2_tlb_xcpt_ma_st : dcache__io_cpu_s2_xcpt_WIRE_ma_st ; reg[63:0] dcache_s2_uncached_data_word ; 
    reg dcache_doUncachedResp ; 
  assign  dcache__io_cpu_replay_next_output = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid & dcache_grantIsUncachedData ; 
    wire dcache__GEN_304 = dcache_s2_valid_hit ==1'h0==1'h0; 
  always @( posedge  dcache_clock )
         begin 
             if ( dcache_reset ==1'h0& dcache__GEN_91 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
                     if (1)$fatal;
                 end 
             if ( dcache_reset ==1'h0& dcache__GEN_97 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:306 assert(!(s1_valid_masked && s1_req.cmd === M_PWR) || (s1_mask_xwr | ~io.cpu.s1_data.mask).andR)\n");
                     if (1)$fatal;
                 end 
             if ( dcache_reset ==1'h0& dcache__GEN_174 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:1162 assert(!needsRead(req) || res)\n");
                     if (1)$fatal;
                 end 
             if ( dcache_reset ==1'h0& dcache__GEN_175 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:487 assert(pstore1_rmw || pstore1_valid_not_rmw(io.cpu.s2_kill) === pstore1_valid)\n");
                     if (1)$fatal;
                 end 
             if ( dcache__GEN_261 & dcache_reset ==1'h0& dcache__GEN_262 )
                 begin 
                     if (1)$error("Assertion failed: A GrantData was unexpected by the dcache.\n    at DCache.scala:654 assert(cached_grant_wait, \"A GrantData was unexpected by the dcache.\")\n");
                     if (1)$fatal;
                 end 
             if ( dcache__GEN_265 & dcache__GEN_266 & dcache_reset ==1'h0& dcache__GEN_267 )
                 begin 
                     if (1)$error("Assertion failed: An AccessAck was unexpected by the dcache.\n    at DCache.scala:664 assert(f, \"An AccessAck was unexpected by the dcache.\") // TODO must handle Ack coming back on same cycle!\n");
                     if (1)$fatal;
                 end 
             if ( dcache__GEN_264 &~ dcache_grantIsUncached & dcache_grantIsVoluntary & dcache_reset ==1'h0& dcache__GEN_269 )
                 begin 
                     if (1)$error("Assertion failed: A ReleaseAck was unexpected by the dcache.\n    at DCache.scala:685 assert(release_ack_wait, \"A ReleaseAck was unexpected by the dcache.\") // TODO should handle Ack coming back on same cycle!\n");
                     if (1)$fatal;
                 end 
             if ( dcache_reset ==1'h0& dcache__GEN_271 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:693 assert(tl_out.e.fire === (tl_out.d.fire && d_first && grantIsCached))\n");
                     if (1)$fatal;
                 end 
             if ( dcache_s2_victimize & dcache_reset ==1'h0& dcache__GEN_286 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:794 assert(s2_valid_flush_line || s2_flush_valid || io.cpu.s2_nack)\n");
                     if (1)$fatal;
                 end 
             if ( dcache_doUncachedResp & dcache_reset ==1'h0& dcache__GEN_304 )
                 begin 
                     if (1)$error("Assertion failed\n    at DCache.scala:928 assert(!s2_valid_hit)\n");
                     if (1)$fatal;
                 end 
         end
    wire[63:0] dcache_s2_data_word_possibly_uncached = dcache_s2_data_word |64'h0; 
    wire[31:0] dcache_io_cpu_resp_bits_data_shifted = dcache_s2_req_addr [2] ?  dcache_s2_data_word_possibly_uncached [63:32]: dcache_s2_data_word_possibly_uncached [31:0]; 
    wire[31:0] dcache_io_cpu_resp_bits_data_zeroed = dcache_io_cpu_resp_bits_data_doZero  ? 32'h0: dcache_io_cpu_resp_bits_data_shifted ; 
    wire[63:0] dcache__GEN_305 ={ dcache_size ==2'h2| dcache_io_cpu_resp_bits_data_doZero  ? ( dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_zeroed [31] ? 32'hFFFFFFFF:32'h0): dcache_s2_data_word_possibly_uncached [63:32], dcache_io_cpu_resp_bits_data_zeroed }; 
    wire[15:0] dcache_io_cpu_resp_bits_data_shifted_1 = dcache_s2_req_addr [1] ?  dcache__GEN_305 [31:16]: dcache__GEN_305 [15:0]; 
    wire[15:0] dcache_io_cpu_resp_bits_data_zeroed_1 = dcache_io_cpu_resp_bits_data_doZero_1  ? 16'h0: dcache_io_cpu_resp_bits_data_shifted_1 ; 
    wire[63:0] dcache__GEN_306 ={ dcache_size ==2'h1| dcache_io_cpu_resp_bits_data_doZero_1  ? ( dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_zeroed_1 [15] ? 48'hFFFFFFFFFFFF:48'h0): dcache__GEN_305 [63:16], dcache_io_cpu_resp_bits_data_zeroed_1 }; 
    wire[7:0] dcache_io_cpu_resp_bits_data_shifted_2 = dcache_s2_req_addr [0] ?  dcache__GEN_306 [15:8]: dcache__GEN_306 [7:0]; 
    wire dcache_io_cpu_resp_bits_data_doZero_2 = dcache_s2_sc &1'h1; 
    wire[7:0] dcache_io_cpu_resp_bits_data_zeroed_2 = dcache_io_cpu_resp_bits_data_doZero_2  ? 8'h0: dcache_io_cpu_resp_bits_data_shifted_2 ; 
    wire[31:0] dcache_io_cpu_resp_bits_data_word_bypass_shifted = dcache_s2_req_addr [2] ?  dcache_s2_data_word_possibly_uncached [63:32]: dcache_s2_data_word_possibly_uncached [31:0]; 
    wire[31:0] dcache_io_cpu_resp_bits_data_word_bypass_zeroed = dcache_io_cpu_resp_bits_data_word_bypass_doZero  ? 32'h0: dcache_io_cpu_resp_bits_data_word_bypass_shifted ;  
    wire dcache_amoalus_0_clock;
    wire dcache_amoalus_0_reset;
    wire[7:0] dcache_amoalus_0_io_mask;
    wire[4:0] dcache_amoalus_0_io_cmd;
    wire[63:0] dcache_amoalus_0_io_lhs;
    wire[63:0] dcache_amoalus_0_io_rhs;
    wire[63:0] dcache_amoalus_0_io_out;
    wire[63:0] dcache_amoalus_0_io_out_unmasked;

    wire[3:0] dcache_amoalus_0_less_signed_mask =4'h2; 
    wire[3:0] dcache_amoalus_0_less_signed_mask_1 =4'h2; 
    wire dcache_amoalus_0_max = dcache_amoalus_0_io_cmd ==5'hD| dcache_amoalus_0_io_cmd ==5'hF; 
    wire dcache_amoalus_0_min = dcache_amoalus_0_io_cmd ==5'hC| dcache_amoalus_0_io_cmd ==5'hE; 
    wire dcache_amoalus_0_add = dcache_amoalus_0_io_cmd ==5'h8; 
    wire dcache_amoalus_0_logic_and = dcache_amoalus_0_io_cmd ==5'hA| dcache_amoalus_0_io_cmd ==5'hB; 
    wire dcache_amoalus_0_logic_xor = dcache_amoalus_0_io_cmd ==5'h9| dcache_amoalus_0_io_cmd ==5'hA; 
    wire[63:0] dcache_amoalus_0_adder_out_mask =~({32'h0,{ dcache_amoalus_0_io_mask [3]==1'h0,31'h0}}|64'h0); 
    wire[64:0] dcache_amoalus_0__GEN ={1'h0, dcache_amoalus_0_io_lhs & dcache_amoalus_0_adder_out_mask }+{1'h0, dcache_amoalus_0_io_rhs & dcache_amoalus_0_adder_out_mask }; 
    wire[63:0] dcache_amoalus_0_adder_out = dcache_amoalus_0__GEN [63:0]; 
    wire dcache_amoalus_0_less_signed =( dcache_amoalus_0_io_cmd &{1'h0, dcache_amoalus_0_less_signed_mask })=={1'h0, dcache_amoalus_0_less_signed_mask &4'hC}; 
    wire dcache_amoalus_0_less_signed_1 =( dcache_amoalus_0_io_cmd &{1'h0, dcache_amoalus_0_less_signed_mask_1 })=={1'h0, dcache_amoalus_0_less_signed_mask_1 &4'hC}; 
    wire dcache_amoalus_0_less = dcache_amoalus_0_io_mask [4] ? ( dcache_amoalus_0_io_lhs [63]== dcache_amoalus_0_io_rhs [63] ?  dcache_amoalus_0_io_lhs [63:32]< dcache_amoalus_0_io_rhs [63:32]| dcache_amoalus_0_io_lhs [63:32]== dcache_amoalus_0_io_rhs [63:32]& dcache_amoalus_0_io_lhs [31:0]< dcache_amoalus_0_io_rhs [31:0]: dcache_amoalus_0_less_signed  ?  dcache_amoalus_0_io_lhs [63]: dcache_amoalus_0_io_rhs [63]): dcache_amoalus_0_io_lhs [31]== dcache_amoalus_0_io_rhs [31] ?  dcache_amoalus_0_io_lhs [31:0]< dcache_amoalus_0_io_rhs [31:0]: dcache_amoalus_0_less_signed_1  ?  dcache_amoalus_0_io_lhs [31]: dcache_amoalus_0_io_rhs [31]; 
    wire[63:0] dcache_amoalus_0_minmax =( dcache_amoalus_0_less  ?  dcache_amoalus_0_min : dcache_amoalus_0_max ) ?  dcache_amoalus_0_io_lhs : dcache_amoalus_0_io_rhs ; 
    wire[63:0] dcache_amoalus_0_logic_0 =( dcache_amoalus_0_logic_and  ?  dcache_amoalus_0_io_lhs & dcache_amoalus_0_io_rhs :64'h0)|( dcache_amoalus_0_logic_xor  ?  dcache_amoalus_0_io_lhs ^ dcache_amoalus_0_io_rhs :64'h0); 
    wire[63:0] dcache_amoalus_0_out = dcache_amoalus_0_add  ?  dcache_amoalus_0_adder_out : dcache_amoalus_0_logic_and | dcache_amoalus_0_logic_xor  ?  dcache_amoalus_0_logic_0 : dcache_amoalus_0_minmax ; 
    wire[15:0] dcache_amoalus_0_wmask_lo_lo ={ dcache_amoalus_0_io_mask [1] ? 8'hFF:8'h0, dcache_amoalus_0_io_mask [0] ? 8'hFF:8'h0}; 
    wire[15:0] dcache_amoalus_0_wmask_lo_hi ={ dcache_amoalus_0_io_mask [3] ? 8'hFF:8'h0, dcache_amoalus_0_io_mask [2] ? 8'hFF:8'h0}; 
    wire[31:0] dcache_amoalus_0_wmask_lo ={ dcache_amoalus_0_wmask_lo_hi , dcache_amoalus_0_wmask_lo_lo }; 
    wire[15:0] dcache_amoalus_0_wmask_hi_lo ={ dcache_amoalus_0_io_mask [5] ? 8'hFF:8'h0, dcache_amoalus_0_io_mask [4] ? 8'hFF:8'h0}; 
    wire[15:0] dcache_amoalus_0_wmask_hi_hi ={ dcache_amoalus_0_io_mask [7] ? 8'hFF:8'h0, dcache_amoalus_0_io_mask [6] ? 8'hFF:8'h0}; 
    wire[31:0] dcache_amoalus_0_wmask_hi ={ dcache_amoalus_0_wmask_hi_hi , dcache_amoalus_0_wmask_hi_lo }; 
    wire[63:0] dcache_amoalus_0_wmask ={ dcache_amoalus_0_wmask_hi , dcache_amoalus_0_wmask_lo }; 
  assign  dcache_amoalus_0_io_out = dcache_amoalus_0_wmask & dcache_amoalus_0_out |~ dcache_amoalus_0_wmask & dcache_amoalus_0_io_lhs ; 
  assign  dcache_amoalus_0_io_out_unmasked = dcache_amoalus_0_out ;
    assign dcache_amoalus_0_clock = dcache_clock;
    assign dcache_amoalus_0_reset = dcache_reset;
    assign dcache_amoalus_0_io_mask = dcache_pstore1_mask;
    assign dcache_amoalus_0_io_cmd = dcache_pstore1_cmd;
    assign dcache_amoalus_0_io_lhs = dcache_s2_data_word;
    assign dcache_amoalus_0_io_rhs = dcache_pstore1_data;
    assign dcache_pstore1_storegen_data = dcache_amoalus_0_io_out;
     
    reg dcache_REG ; 
    wire dcache__GEN_307 = dcache_REG  ? 1'h1: dcache_resetting ; 
    wire[6:0] dcache_flushCounterNext ={1'h0, dcache_flushCounter }+7'h1; 
    wire dcache_flushDone =&( dcache_flushCounterNext [6]); 
    wire[5:0] dcache_flushCounterWrap = dcache_flushCounterNext [5:0]; 
  assign  dcache_metaArb_io_in_5_valid = dcache_flushing & dcache_flushed ==1'h0; 
  assign  dcache_metaArb_io_in_5_bits_addr ={ dcache_io_cpu_req_bits_addr [33:12],{ dcache_metaArb_io_in_5_bits_idx ,6'h0}}; 
    wire[1:0] dcache_metaArb_io_in_0_bits_data_meta_1_coh_state = dcache_metaArb_io_in_0_bits_data_meta_state ; 
    wire[19:0] dcache_metaArb_io_in_0_bits_data_meta_1_tag =20'h0; 
  assign  dcache_metaArb_io_in_0_bits_data ={ dcache_metaArb_io_in_0_bits_data_meta_1_coh_state , dcache_metaArb_io_in_0_bits_data_meta_1_tag }; 
    wire dcache__GEN_308 = dcache_tl_out_a_ready & dcache_tl_out_a_valid ; 
    wire[26:0] dcache__GEN_309 =27'hFFF<< dcache_tl_out_a_bits_size ; 
    wire[11:0] dcache__GEN_310 =~( dcache__GEN_309 [11:0]); 
    wire[8:0] dcache_io_cpu_perf_acquire_beats1_decode = dcache__GEN_310 [11:3]; 
    wire dcache_io_cpu_perf_acquire_beats1_opdata = dcache_tl_out_a_bits_opcode [2]==1'h0; 
    wire[8:0] dcache_io_cpu_perf_acquire_beats1 = dcache_io_cpu_perf_acquire_beats1_opdata  ?  dcache_io_cpu_perf_acquire_beats1_decode :9'h0; reg[8:0] dcache_io_cpu_perf_acquire_counter ; 
    wire[9:0] dcache__GEN_311 ={1'h0, dcache_io_cpu_perf_acquire_counter }-10'h1; 
    wire[8:0] dcache_io_cpu_perf_acquire_counter1 = dcache__GEN_311 [8:0]; 
    wire dcache_io_cpu_perf_acquire_first = dcache_io_cpu_perf_acquire_counter ==9'h0; 
    wire dcache_io_cpu_perf_acquire_last = dcache_io_cpu_perf_acquire_counter ==9'h1| dcache_io_cpu_perf_acquire_beats1 ==9'h0; 
    wire dcache_io_cpu_perf_acquire_done = dcache_io_cpu_perf_acquire_last & dcache__GEN_308 ; 
    wire[8:0] dcache_io_cpu_perf_acquire_count = dcache_io_cpu_perf_acquire_beats1 &~ dcache_io_cpu_perf_acquire_counter1 ; 
    wire dcache__GEN_312 = dcache_nodeOut_c_ready & dcache_nodeOut_c_valid ; 
    wire[26:0] dcache__GEN_313 =27'hFFF<< dcache_nodeOut_c_bits_size ; 
    wire[11:0] dcache__GEN_314 =~( dcache__GEN_313 [11:0]); 
    wire[8:0] dcache_io_cpu_perf_release_beats1_decode = dcache__GEN_314 [11:3]; 
    wire dcache_io_cpu_perf_release_beats1_opdata = dcache_nodeOut_c_bits_opcode [0]; 
    wire[8:0] dcache_io_cpu_perf_release_beats1 = dcache_io_cpu_perf_release_beats1_opdata  ?  dcache_io_cpu_perf_release_beats1_decode :9'h0; reg[8:0] dcache_io_cpu_perf_release_counter ; 
    wire[9:0] dcache__GEN_315 ={1'h0, dcache_io_cpu_perf_release_counter }-10'h1; 
    wire[8:0] dcache_io_cpu_perf_release_counter1 = dcache__GEN_315 [8:0]; 
    wire dcache_io_cpu_perf_release_first = dcache_io_cpu_perf_release_counter ==9'h0; 
    wire dcache_io_cpu_perf_release_last = dcache_io_cpu_perf_release_counter ==9'h1| dcache_io_cpu_perf_release_beats1 ==9'h0; 
    wire dcache_io_cpu_perf_release_done = dcache_io_cpu_perf_release_last & dcache__GEN_312 ; 
    wire[8:0] dcache_io_cpu_perf_release_count = dcache_io_cpu_perf_release_beats1 &~ dcache_io_cpu_perf_release_counter1 ; 
    wire dcache__io_cpu_perf_canAcceptStoreThenLoad_output =( dcache_s2_valid & dcache_s2_write & dcache_pstore1_rmw & dcache_s1_valid & dcache_s1_write & dcache_s1_waw_hazard ==1'h0| dcache_pstore2_valid & dcache_pstore1_valid_likely & dcache_s1_valid & dcache_s1_write )==1'h0; reg[2:0] dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count ; 
    wire dcache__GEN_316 = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid & dcache_grantIsRefill ; 
    wire[3:0] dcache__GEN_317 ={1'h0, dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count }+4'h1; 
    wire dcache_io_cpu_perf_blocked_near_end_of_refill = dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count >=3'h6; 
    reg dcache_data_error ; 
    reg dcache_data_error_uncorrectable ; 
    wire[31:0] dcache_error_addr ={ dcache_metaArb_io_in_1_valid  ? { dcache_s2_meta_corrected_0_tag , dcache_metaArb_io_in_1_bits_addr [11:6]}: dcache_probe_bits_address [31:6],6'h0}; 
    wire dcache__io_errors_bus_valid_output = dcache_nodeOut_d_ready & dcache_nodeOut_d_valid &( dcache_nodeOut_d_bits_denied | dcache_nodeOut_d_bits_corrupt ); 
    wire[33:0] dcache__GEN_318 = dcache_grantIsCached  ? { dcache_s2_req_addr [33:6],6'h0}:34'h0; 
    wire dcache__GEN_319 = dcache_s2_valid_data_error ==1'h0; 
    wire dcache__GEN_320 = dcache_s2_valid_data_error & dcache_s2_data_error_uncorrectable ==1'h0; 
    wire dcache__GEN_321 = dcache_s2_valid_data_error & dcache_s2_data_error_uncorrectable ; 
    wire dcache__GEN_322 = dcache_s2_victim_dirty ==1'h0; 
    wire dcache__GEN_323 = dcache_s2_meta_error ==1'h0; 
    wire dcache__GEN_324 = dcache_s2_meta_error & dcache_s2_meta_error_uncorrectable ==1'h0; 
    wire dcache__GEN_325 = dcache_s2_meta_error & dcache_s2_meta_error_uncorrectable ; 
  always @( posedge  dcache_clock )
         begin  
             dcache_clock_en_reg  <=1'h1;
             if ( dcache_s2_victimize )
                 begin  
                     dcache_probe_bits_opcode  <= dcache_probe_bits_res_opcode ; 
                     dcache_probe_bits_param  <= dcache_probe_bits_res_param ; 
                     dcache_probe_bits_size  <= dcache_probe_bits_res_size ; 
                     dcache_probe_bits_source  <= dcache_probe_bits_res_source ; 
                     dcache_probe_bits_address  <= dcache_probe_bits_res_address ; 
                     dcache_probe_bits_mask  <= dcache_probe_bits_res_mask ; 
                     dcache_probe_bits_data  <= dcache_probe_bits_res_data ; 
                     dcache_probe_bits_corrupt  <= dcache_probe_bits_res_corrupt ;
                 end 
              else 
                 if ( dcache__GEN_88 )
                     begin  
                         dcache_probe_bits_opcode  <= dcache_nodeOut_b_bits_opcode ; 
                         dcache_probe_bits_param  <= dcache_nodeOut_b_bits_param ; 
                         dcache_probe_bits_size  <= dcache_nodeOut_b_bits_size ; 
                         dcache_probe_bits_source  <= dcache_nodeOut_b_bits_source ; 
                         dcache_probe_bits_address  <= dcache_nodeOut_b_bits_address ; 
                         dcache_probe_bits_mask  <= dcache_nodeOut_b_bits_mask ; 
                         dcache_probe_bits_data  <= dcache_nodeOut_b_bits_data ; 
                         dcache_probe_bits_corrupt  <= dcache_nodeOut_b_bits_corrupt ;
                     end 
                  else 
                     begin 
                     end 
             if ( dcache_s0_clk_en )
                 begin  
                     dcache_s1_req_addr  <= dcache_s0_req_addr ; 
                     dcache_s1_req_tag  <= dcache_s0_req_tag ; 
                     dcache_s1_req_cmd  <= dcache_s0_req_cmd ; 
                     dcache_s1_req_size  <= dcache_s0_req_size ; 
                     dcache_s1_req_signed  <= dcache_s0_req_signed ; 
                     dcache_s1_req_dprv  <= dcache_s0_req_dprv ; 
                     dcache_s1_req_dv  <= dcache_s0_req_dv ; 
                     dcache_s1_req_phys  <= dcache_s0_req_phys ; 
                     dcache_s1_req_no_alloc  <= dcache_s0_req_no_alloc ; 
                     dcache_s1_req_no_xcpt  <= dcache_s0_req_no_xcpt ; 
                     dcache_s1_req_data  <= dcache_s0_req_data ; 
                     dcache_s1_req_mask  <= dcache_s0_req_mask ; 
                     dcache_s1_did_read  <= dcache__GEN_93 ; 
                     dcache_s1_read_mask  <= dcache_dataArb_io_in_3_bits_wordMask ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache__GEN_90 )
                 begin  
                     dcache_s1_tlb_req_vaddr  <= dcache_s0_tlb_req_vaddr ; 
                     dcache_s1_tlb_req_passthrough  <= dcache_s0_tlb_req_passthrough ; 
                     dcache_s1_tlb_req_size  <= dcache_s0_tlb_req_size ; 
                     dcache_s1_tlb_req_cmd  <= dcache_s0_tlb_req_cmd ; 
                     dcache_s1_tlb_req_prv  <= dcache_s0_tlb_req_prv ; 
                     dcache_s1_tlb_req_v  <= dcache_s0_tlb_req_v ;
                 end 
              else 
                 begin 
                 end  
             dcache_s1_flush_valid  <= dcache_metaArb_io_in_5_ready & dcache_metaArb_io_in_5_valid & dcache_s1_flush_valid ==1'h0& dcache_s2_flush_valid_pre_tag_ecc ==1'h0& dcache_release_state ==4'h0& dcache_release_ack_wait ==1'h0;
             if ( dcache__GEN_300 )
                 begin 
                     if ( dcache__GEN_302 ) 
                         dcache_release_ack_addr  <= dcache_probe_bits_address ;
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end 
             if ( dcache__GEN_248 )
                 begin 
                     if ( dcache_s2_uncached )
                         begin 
                             if ( dcache_a_sel )
                                 begin  
                                     dcache_uncachedReqs_0_addr  <= dcache_s2_req_addr ; 
                                     dcache_uncachedReqs_0_tag  <= dcache_s2_req_tag ; 
                                     dcache_uncachedReqs_0_cmd  <= dcache__GEN_250 ; 
                                     dcache_uncachedReqs_0_size  <= dcache_s2_req_size ; 
                                     dcache_uncachedReqs_0_signed  <= dcache_s2_req_signed ; 
                                     dcache_uncachedReqs_0_dprv  <= dcache_s2_req_dprv ; 
                                     dcache_uncachedReqs_0_dv  <= dcache_s2_req_dv ; 
                                     dcache_uncachedReqs_0_phys  <= dcache_s2_req_phys ; 
                                     dcache_uncachedReqs_0_no_alloc  <= dcache_s2_req_no_alloc ; 
                                     dcache_uncachedReqs_0_no_xcpt  <= dcache_s2_req_no_xcpt ; 
                                     dcache_uncachedReqs_0_data  <= dcache_s2_req_data ; 
                                     dcache_uncachedReqs_0_mask  <= dcache_s2_req_mask ;
                                 end 
                              else 
                                 begin 
                                 end 
                         end 
                      else  
                         dcache_refill_way  <= dcache_s2_victim_or_hit_way ;
                 end 
              else 
                 begin 
                 end  
             dcache_s2_not_nacked_in_s1  <= dcache_s1_nack ==1'h0;
             if ( dcache__GEN_260 )
                 begin 
                     if ( dcache_grantIsCached )
                         begin 
                             if ( dcache__GEN_98 )
                                 begin  
                                     dcache_s2_req_addr  <= dcache__GEN_103 ; 
                                     dcache_s2_req_tag  <= dcache_s1_req_tag ; 
                                     dcache_s2_req_cmd  <= dcache_s1_req_cmd ; 
                                     dcache_s2_req_size  <= dcache_s1_req_size ; 
                                     dcache_s2_req_signed  <= dcache_s1_req_signed ;
                                 end 
                              else 
                                 begin 
                                 end 
                         end 
                      else 
                         if ( dcache_grantIsUncached )
                             begin 
                                 if ( dcache_grantIsUncachedData )
                                     begin  
                                         dcache_s2_req_addr  <= dcache__GEN_268 ; 
                                         dcache_s2_req_tag  <= dcache_uncachedResp_tag ; 
                                         dcache_s2_req_cmd  <=5'h0; 
                                         dcache_s2_req_size  <= dcache_uncachedResp_size ; 
                                         dcache_s2_req_signed  <= dcache_uncachedResp_signed ; 
                                         dcache_s2_uncached_resp_addr  <= dcache_uncachedResp_addr ;
                                     end 
                                  else 
                                     if ( dcache__GEN_98 )
                                         begin  
                                             dcache_s2_req_addr  <= dcache__GEN_103 ; 
                                             dcache_s2_req_tag  <= dcache_s1_req_tag ; 
                                             dcache_s2_req_cmd  <= dcache_s1_req_cmd ; 
                                             dcache_s2_req_size  <= dcache_s1_req_size ; 
                                             dcache_s2_req_signed  <= dcache_s1_req_signed ;
                                         end 
                                      else 
                                         begin 
                                         end 
                             end 
                          else 
                             if ( dcache__GEN_98 )
                                 begin  
                                     dcache_s2_req_addr  <= dcache__GEN_103 ; 
                                     dcache_s2_req_tag  <= dcache_s1_req_tag ; 
                                     dcache_s2_req_cmd  <= dcache_s1_req_cmd ; 
                                     dcache_s2_req_size  <= dcache_s1_req_size ; 
                                     dcache_s2_req_signed  <= dcache_s1_req_signed ;
                                 end 
                              else 
                                 begin 
                                 end 
                 end 
              else 
                 if ( dcache__GEN_98 )
                     begin  
                         dcache_s2_req_addr  <= dcache__GEN_103 ; 
                         dcache_s2_req_tag  <= dcache_s1_req_tag ; 
                         dcache_s2_req_cmd  <= dcache_s1_req_cmd ; 
                         dcache_s2_req_size  <= dcache_s1_req_size ; 
                         dcache_s2_req_signed  <= dcache_s1_req_signed ;
                     end 
                  else 
                     begin 
                     end 
             if ( dcache__GEN_98 )
                 begin  
                     dcache_s2_req_dprv  <= dcache_s1_req_dprv ; 
                     dcache_s2_req_dv  <= dcache_s1_req_dv ; 
                     dcache_s2_req_phys  <= dcache_s1_req_phys ; 
                     dcache_s2_req_no_alloc  <= dcache_s1_req_no_alloc ; 
                     dcache_s2_req_no_xcpt  <= dcache_s1_req_no_xcpt ; 
                     dcache_s2_req_data  <= dcache_s1_req_data ; 
                     dcache_s2_req_mask  <= dcache_s1_req_mask ; 
                     dcache_s2_tlb_xcpt_miss  <= dcache_tlb_io_resp_miss ; 
                     dcache_s2_tlb_xcpt_paddr  <= dcache_tlb_io_resp_paddr ; 
                     dcache_s2_tlb_xcpt_gpa  <= dcache_tlb_io_resp_gpa ; 
                     dcache_s2_tlb_xcpt_gpa_is_pte  <= dcache_tlb_io_resp_gpa_is_pte ; 
                     dcache_s2_tlb_xcpt_pf_ld  <= dcache_tlb_io_resp_pf_ld ; 
                     dcache_s2_tlb_xcpt_pf_st  <= dcache_tlb_io_resp_pf_st ; 
                     dcache_s2_tlb_xcpt_pf_inst  <= dcache_tlb_io_resp_pf_inst ; 
                     dcache_s2_tlb_xcpt_gf_ld  <= dcache_tlb_io_resp_gf_ld ; 
                     dcache_s2_tlb_xcpt_gf_st  <= dcache_tlb_io_resp_gf_st ; 
                     dcache_s2_tlb_xcpt_gf_inst  <= dcache_tlb_io_resp_gf_inst ; 
                     dcache_s2_tlb_xcpt_ae_ld  <= dcache_tlb_io_resp_ae_ld ; 
                     dcache_s2_tlb_xcpt_ae_st  <= dcache_tlb_io_resp_ae_st ; 
                     dcache_s2_tlb_xcpt_ae_inst  <= dcache_tlb_io_resp_ae_inst ; 
                     dcache_s2_tlb_xcpt_ma_ld  <= dcache_tlb_io_resp_ma_ld ; 
                     dcache_s2_tlb_xcpt_ma_st  <= dcache_tlb_io_resp_ma_st ; 
                     dcache_s2_tlb_xcpt_ma_inst  <= dcache_tlb_io_resp_ma_inst ; 
                     dcache_s2_tlb_xcpt_cacheable  <= dcache_tlb_io_resp_cacheable ; 
                     dcache_s2_tlb_xcpt_must_alloc  <= dcache_tlb_io_resp_must_alloc ; 
                     dcache_s2_tlb_xcpt_prefetchable  <= dcache_tlb_io_resp_prefetchable ; 
                     dcache_s2_pma_miss  <= dcache__GEN_105 ; 
                     dcache_s2_pma_paddr  <= dcache__GEN_106 ; 
                     dcache_s2_pma_gpa  <= dcache__GEN_107 ; 
                     dcache_s2_pma_gpa_is_pte  <= dcache__GEN_108 ; 
                     dcache_s2_pma_pf_ld  <= dcache__GEN_109 ; 
                     dcache_s2_pma_pf_st  <= dcache__GEN_110 ; 
                     dcache_s2_pma_pf_inst  <= dcache__GEN_111 ; 
                     dcache_s2_pma_gf_ld  <= dcache__GEN_112 ; 
                     dcache_s2_pma_gf_st  <= dcache__GEN_113 ; 
                     dcache_s2_pma_gf_inst  <= dcache__GEN_114 ; 
                     dcache_s2_pma_ae_ld  <= dcache__GEN_115 ; 
                     dcache_s2_pma_ae_st  <= dcache__GEN_116 ; 
                     dcache_s2_pma_ae_inst  <= dcache__GEN_117 ; 
                     dcache_s2_pma_ma_ld  <= dcache__GEN_118 ; 
                     dcache_s2_pma_ma_st  <= dcache__GEN_119 ; 
                     dcache_s2_pma_ma_inst  <= dcache__GEN_120 ; 
                     dcache_s2_pma_cacheable  <= dcache__GEN_121 ; 
                     dcache_s2_pma_must_alloc  <= dcache__GEN_122 ; 
                     dcache_s2_pma_prefetchable  <= dcache__GEN_123 ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache__GEN_124 ) 
                 dcache_s2_vaddr_r  <= dcache_s1_vaddr ;
              else 
                 begin 
                 end  
             dcache_s2_flush_valid_pre_tag_ecc  <= dcache_s1_flush_valid ;
             if ( dcache_s1_meta_clk_en )
                 begin  
                     dcache_s2_meta_correctable_errors  <=1'h0; 
                     dcache_s2_meta_uncorrectable_errors  <=1'h0; 
                     dcache_s2_meta_corrected_r  <= dcache_tag_array_s1_meta_data_0 ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache_s2_data_en ) 
                 dcache_s2_data  <= dcache__s2_data_WIRE ;
              else 
                 begin 
                 end 
             if ( dcache_s1_probe )
                 begin  
                     dcache_s2_probe_way  <= dcache_s1_hit_way ; 
                     dcache_s2_probe_state_state  <= dcache_s1_hit_state_state ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache_s1_valid_not_nacked )
                 begin  
                     dcache_s2_hit_way  <= dcache_s1_hit_way ; 
                     dcache_s2_waw_hazard  <= dcache_s1_waw_hazard ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache__GEN_126 ) 
                 dcache_s2_hit_state_state  <= dcache_s1_hit_state_state ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_135 ) 
                 dcache_s2_victim_way_r  <= dcache_s1_victim_way ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_162 ) 
                 dcache_lrscAddr  <= dcache_s2_req_addr [33:6];
              else 
                 begin 
                 end  
             dcache_s2_correct_REG  <= dcache_any_pstore_valid | dcache_s2_valid ;
             if ( dcache__GEN_167 ) 
                 dcache_pstore1_cmd  <= dcache_s1_req_cmd ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_168 ) 
                 dcache_pstore1_addr  <= dcache_s1_vaddr ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_169 ) 
                 dcache_pstore1_data  <= dcache_io_cpu_s1_data_data ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_170 ) 
                 dcache_pstore1_way  <= dcache_s1_hit_way ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_171 ) 
                 dcache_pstore1_mask  <= dcache_s1_mask ;
              else 
                 begin 
                 end 
             if ( dcache__GEN_173 ) 
                 dcache_pstore1_rmw_r  <= dcache__GEN_172 ;
              else 
                 begin 
                 end  
             dcache_pstore_drain_on_miss_REG  <= dcache__io_cpu_s2_nack_output ;
             if ( dcache_advance_pstore1 )
                 begin  
                     dcache_pstore2_addr  <= dcache__GEN_176 ; 
                     dcache_pstore2_way  <= dcache__GEN_177 ;
                 end 
              else 
                 begin 
                 end 
             if ( dcache__GEN_178 ) 
                 dcache_pstore2_storegen_data_r  <= dcache_pstore1_storegen_data [7:0];
              else 
                 begin 
                 end 
             if ( dcache__GEN_179 ) 
                 dcache_pstore2_storegen_data_r_1  <= dcache_pstore1_storegen_data [15:8];
              else 
                 begin 
                 end 
             if ( dcache__GEN_180 ) 
                 dcache_pstore2_storegen_data_r_2  <= dcache_pstore1_storegen_data [23:16];
              else 
                 begin 
                 end 
             if ( dcache__GEN_181 ) 
                 dcache_pstore2_storegen_data_r_3  <= dcache_pstore1_storegen_data [31:24];
              else 
                 begin 
                 end 
             if ( dcache__GEN_182 ) 
                 dcache_pstore2_storegen_data_r_4  <= dcache_pstore1_storegen_data [39:32];
              else 
                 begin 
                 end 
             if ( dcache__GEN_183 ) 
                 dcache_pstore2_storegen_data_r_5  <= dcache_pstore1_storegen_data [47:40];
              else 
                 begin 
                 end 
             if ( dcache__GEN_184 ) 
                 dcache_pstore2_storegen_data_r_6  <= dcache_pstore1_storegen_data [55:48];
              else 
                 begin 
                 end 
             if ( dcache__GEN_185 ) 
                 dcache_pstore2_storegen_data_r_7  <= dcache_pstore1_storegen_data [63:56];
              else 
                 begin 
                 end 
             if ( dcache__GEN_186 ) 
                 dcache_pstore2_storegen_mask  <= dcache__GEN_187 ;
              else 
                 begin 
                 end  
             dcache_io_cpu_s2_nack_cause_raw_REG  <= dcache_s1_raw_hazard ;
             if ( dcache__GEN_276 )
                 begin 
                     if ( dcache_nodeOut_d_valid ) 
                         dcache_blockUncachedGrant  <= dcache__GEN_277 ;
                      else  
                         dcache_blockUncachedGrant  <= dcache_dataArb_io_out_valid ;
                 end 
              else  
                 dcache_blockUncachedGrant  <= dcache_dataArb_io_out_valid ; 
             dcache_s1_release_data_valid  <= dcache_dataArb_io_in_2_ready & dcache_dataArb_io_in_2_valid ; 
             dcache_s2_release_data_valid  <= dcache_s1_release_data_valid & dcache_releaseRejected ==1'h0; 
             dcache_io_cpu_s2_xcpt_REG  <= dcache_s1_xcpt_valid ;
             if ( dcache__io_cpu_replay_next_output ) 
                 dcache_s2_uncached_data_word  <= dcache_s1_uncached_data_word ;
              else 
                 begin 
                 end  
             dcache_doUncachedResp  <= dcache__io_cpu_replay_next_output ; 
             dcache_REG  <= dcache_reset ; 
             dcache_data_error  <= dcache_nodeOut_c_ready & dcache_nodeOut_c_valid & dcache_inWriteback & dcache_s2_data_error ; 
             dcache_data_error_uncorrectable  <= dcache_s2_data_error_uncorrectable ;
         end
  always @( posedge  dcache_tlb_clock )
         begin 
             if ( dcache_tlb_do_refill )
                 begin 
                     if ( dcache__GEN_2 )
                         begin  
                             dcache_tlb_special_entry_level  <= dcache_tlb_io_ptw_resp_bits_level ; 
                             dcache_tlb_special_entry_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                             dcache_tlb_special_entry_tag_v  <= dcache_tlb_refill_v ; 
                             dcache_tlb_special_entry_data_0  <= dcache__GEN_3 ; 
                             dcache_tlb_special_entry_valid_0  <=1'h1;
                         end 
                      else 
                         if ( dcache__GEN_5 )
                             begin 
                                 if ( dcache__GEN_7 )
                                     begin  
                                         dcache_tlb_superpage_entries_0_level  <= dcache__GEN_8 ; 
                                         dcache_tlb_superpage_entries_0_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                                         dcache_tlb_superpage_entries_0_tag_v  <= dcache_tlb_refill_v ; 
                                         dcache_tlb_superpage_entries_0_data_0  <= dcache__GEN_9 ; 
                                         dcache_tlb_superpage_entries_0_valid_0  <= dcache__GEN_10 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_11 )
                                     begin  
                                         dcache_tlb_superpage_entries_1_level  <= dcache__GEN_12 ; 
                                         dcache_tlb_superpage_entries_1_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                                         dcache_tlb_superpage_entries_1_tag_v  <= dcache_tlb_refill_v ; 
                                         dcache_tlb_superpage_entries_1_data_0  <= dcache__GEN_13 ; 
                                         dcache_tlb_superpage_entries_1_valid_0  <= dcache__GEN_14 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_15 )
                                     begin  
                                         dcache_tlb_superpage_entries_2_level  <= dcache__GEN_16 ; 
                                         dcache_tlb_superpage_entries_2_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                                         dcache_tlb_superpage_entries_2_tag_v  <= dcache_tlb_refill_v ; 
                                         dcache_tlb_superpage_entries_2_data_0  <= dcache__GEN_17 ; 
                                         dcache_tlb_superpage_entries_2_valid_0  <= dcache__GEN_18 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_19 )
                                     begin  
                                         dcache_tlb_superpage_entries_3_level  <= dcache__GEN_20 ; 
                                         dcache_tlb_superpage_entries_3_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                                         dcache_tlb_superpage_entries_3_tag_v  <= dcache_tlb_refill_v ; 
                                         dcache_tlb_superpage_entries_3_data_0  <= dcache__GEN_21 ; 
                                         dcache_tlb_superpage_entries_3_valid_0  <= dcache__GEN_22 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin  
                                 dcache_tlb_sectored_entries_0_0_level  <=2'h0; 
                                 dcache_tlb_sectored_entries_0_0_tag_vpn  <= dcache_tlb_r_refill_tag ; 
                                 dcache_tlb_sectored_entries_0_0_tag_v  <= dcache_tlb_refill_v ;
                                 if ( dcache__GEN_30 ) 
                                     dcache_tlb_sectored_entries_0_0_data_0  <= dcache__GEN_29 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_31 ) 
                                     dcache_tlb_sectored_entries_0_0_data_1  <= dcache__GEN_29 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_32 ) 
                                     dcache_tlb_sectored_entries_0_0_data_2  <= dcache__GEN_29 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_33 ) 
                                     dcache_tlb_sectored_entries_0_0_data_3  <= dcache__GEN_29 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache_tlb_invalidate_refill )
                                     begin  
                                         dcache_tlb_sectored_entries_0_0_valid_0  <=1'h0; 
                                         dcache_tlb_sectored_entries_0_0_valid_1  <=1'h0; 
                                         dcache_tlb_sectored_entries_0_0_valid_2  <=1'h0; 
                                         dcache_tlb_sectored_entries_0_0_valid_3  <=1'h0;
                                     end 
                                  else 
                                     begin 
                                         if ( dcache__GEN_25 ) 
                                             dcache_tlb_sectored_entries_0_0_valid_0  <=1'h1;
                                          else 
                                             if ( dcache__GEN_24 ) 
                                                 dcache_tlb_sectored_entries_0_0_valid_0  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_26 ) 
                                             dcache_tlb_sectored_entries_0_0_valid_1  <=1'h1;
                                          else 
                                             if ( dcache__GEN_24 ) 
                                                 dcache_tlb_sectored_entries_0_0_valid_1  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_27 ) 
                                             dcache_tlb_sectored_entries_0_0_valid_2  <=1'h1;
                                          else 
                                             if ( dcache__GEN_24 ) 
                                                 dcache_tlb_sectored_entries_0_0_valid_2  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_28 ) 
                                             dcache_tlb_sectored_entries_0_0_valid_3  <=1'h1;
                                          else 
                                             if ( dcache__GEN_24 ) 
                                                 dcache_tlb_sectored_entries_0_0_valid_3  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                     end 
                             end  
                     dcache_tlb_r_gpa_valid  <= dcache_tlb_io_ptw_resp_bits_gpa_valid ; 
                     dcache_tlb_r_gpa  <= dcache_tlb_io_ptw_resp_bits_gpa_bits ; 
                     dcache_tlb_r_gpa_is_pte  <= dcache_tlb_io_ptw_resp_bits_gpa_is_pte ;
                 end 
              else 
                 begin 
                 end 
         end
  always @( posedge  dcache_tlb_clock )
         begin 
             if ( dcache_tlb_reset )
                 begin  
                     dcache_tlb_state  <=2'h0; 
                     dcache_tlb_v_entries_use_stage1  <=1'h0; 
                     dcache_tlb_state_reg_1  <=3'h0;
                 end 
              else 
                 if ( dcache__GEN_35 )
                     begin 
                         if ( dcache__GEN_36 ) 
                             dcache_tlb_state_reg_1  <= dcache__GEN_39 ;
                          else 
                             begin 
                             end 
                     end 
                  else 
                     begin 
                     end 
         end
  always @( posedge  dcache_pma_checker_clock )
         begin 
             if ( dcache_pma_checker_do_refill )
                 begin 
                     if ( dcache__GEN_42 )
                         begin  
                             dcache_pma_checker_special_entry_level  <= dcache_pma_checker_io_ptw_resp_bits_level ; 
                             dcache_pma_checker_special_entry_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                             dcache_pma_checker_special_entry_tag_v  <= dcache_pma_checker_refill_v ; 
                             dcache_pma_checker_special_entry_data_0  <= dcache__GEN_43 ; 
                             dcache_pma_checker_special_entry_valid_0  <=1'h1;
                         end 
                      else 
                         if ( dcache__GEN_45 )
                             begin 
                                 if ( dcache__GEN_47 )
                                     begin  
                                         dcache_pma_checker_superpage_entries_0_level  <= dcache__GEN_48 ; 
                                         dcache_pma_checker_superpage_entries_0_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                                         dcache_pma_checker_superpage_entries_0_tag_v  <= dcache_pma_checker_refill_v ; 
                                         dcache_pma_checker_superpage_entries_0_data_0  <= dcache__GEN_49 ; 
                                         dcache_pma_checker_superpage_entries_0_valid_0  <= dcache__GEN_50 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_51 )
                                     begin  
                                         dcache_pma_checker_superpage_entries_1_level  <= dcache__GEN_52 ; 
                                         dcache_pma_checker_superpage_entries_1_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                                         dcache_pma_checker_superpage_entries_1_tag_v  <= dcache_pma_checker_refill_v ; 
                                         dcache_pma_checker_superpage_entries_1_data_0  <= dcache__GEN_53 ; 
                                         dcache_pma_checker_superpage_entries_1_valid_0  <= dcache__GEN_54 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_55 )
                                     begin  
                                         dcache_pma_checker_superpage_entries_2_level  <= dcache__GEN_56 ; 
                                         dcache_pma_checker_superpage_entries_2_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                                         dcache_pma_checker_superpage_entries_2_tag_v  <= dcache_pma_checker_refill_v ; 
                                         dcache_pma_checker_superpage_entries_2_data_0  <= dcache__GEN_57 ; 
                                         dcache_pma_checker_superpage_entries_2_valid_0  <= dcache__GEN_58 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_59 )
                                     begin  
                                         dcache_pma_checker_superpage_entries_3_level  <= dcache__GEN_60 ; 
                                         dcache_pma_checker_superpage_entries_3_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                                         dcache_pma_checker_superpage_entries_3_tag_v  <= dcache_pma_checker_refill_v ; 
                                         dcache_pma_checker_superpage_entries_3_data_0  <= dcache__GEN_61 ; 
                                         dcache_pma_checker_superpage_entries_3_valid_0  <= dcache__GEN_62 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin  
                                 dcache_pma_checker_sectored_entries_0_0_level  <=2'h0; 
                                 dcache_pma_checker_sectored_entries_0_0_tag_vpn  <= dcache_pma_checker_r_refill_tag ; 
                                 dcache_pma_checker_sectored_entries_0_0_tag_v  <= dcache_pma_checker_refill_v ;
                                 if ( dcache__GEN_70 ) 
                                     dcache_pma_checker_sectored_entries_0_0_data_0  <= dcache__GEN_69 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_71 ) 
                                     dcache_pma_checker_sectored_entries_0_0_data_1  <= dcache__GEN_69 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_72 ) 
                                     dcache_pma_checker_sectored_entries_0_0_data_2  <= dcache__GEN_69 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache__GEN_73 ) 
                                     dcache_pma_checker_sectored_entries_0_0_data_3  <= dcache__GEN_69 ;
                                  else 
                                     begin 
                                     end 
                                 if ( dcache_pma_checker_invalidate_refill )
                                     begin  
                                         dcache_pma_checker_sectored_entries_0_0_valid_0  <=1'h0; 
                                         dcache_pma_checker_sectored_entries_0_0_valid_1  <=1'h0; 
                                         dcache_pma_checker_sectored_entries_0_0_valid_2  <=1'h0; 
                                         dcache_pma_checker_sectored_entries_0_0_valid_3  <=1'h0;
                                     end 
                                  else 
                                     begin 
                                         if ( dcache__GEN_65 ) 
                                             dcache_pma_checker_sectored_entries_0_0_valid_0  <=1'h1;
                                          else 
                                             if ( dcache__GEN_64 ) 
                                                 dcache_pma_checker_sectored_entries_0_0_valid_0  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_66 ) 
                                             dcache_pma_checker_sectored_entries_0_0_valid_1  <=1'h1;
                                          else 
                                             if ( dcache__GEN_64 ) 
                                                 dcache_pma_checker_sectored_entries_0_0_valid_1  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_67 ) 
                                             dcache_pma_checker_sectored_entries_0_0_valid_2  <=1'h1;
                                          else 
                                             if ( dcache__GEN_64 ) 
                                                 dcache_pma_checker_sectored_entries_0_0_valid_2  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( dcache__GEN_68 ) 
                                             dcache_pma_checker_sectored_entries_0_0_valid_3  <=1'h1;
                                          else 
                                             if ( dcache__GEN_64 ) 
                                                 dcache_pma_checker_sectored_entries_0_0_valid_3  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                     end 
                             end  
                     dcache_pma_checker_r_gpa_valid  <= dcache_pma_checker_io_ptw_resp_bits_gpa_valid ; 
                     dcache_pma_checker_r_gpa  <= dcache_pma_checker_io_ptw_resp_bits_gpa_bits ; 
                     dcache_pma_checker_r_gpa_is_pte  <= dcache_pma_checker_io_ptw_resp_bits_gpa_is_pte ;
                 end 
              else 
                 begin 
                 end 
         end
  always @( posedge  dcache_pma_checker_clock )
         begin 
             if ( dcache_pma_checker_reset )
                 begin  
                     dcache_pma_checker_state  <=2'h0; 
                     dcache_pma_checker_v_entries_use_stage1  <=1'h0; 
                     dcache_pma_checker_state_reg_1  <=3'h0;
                 end 
              else 
                 if ( dcache__GEN_75 )
                     begin 
                         if ( dcache__GEN_76 ) 
                             dcache_pma_checker_state_reg_1  <= dcache__GEN_79 ;
                          else 
                             begin 
                             end 
                     end 
                  else 
                     begin 
                     end 
         end
  always @( posedge  dcache_clock )
         begin 
             if ( dcache_reset )
                 begin  
                     dcache_s1_valid  <=1'h0; 
                     dcache_s1_probe  <=1'h0; 
                     dcache_s1_tlb_req_valid  <=1'h0; 
                     dcache_s2_tlb_req_valid  <=1'h0; 
                     dcache_flushed  <=1'h1; 
                     dcache_flushing  <=1'h0; 
                     dcache_cached_grant_wait  <=1'h0; 
                     dcache_resetting  <=1'h0; 
                     dcache_flushCounter  <=6'h0; 
                     dcache_release_ack_wait  <=1'h0; 
                     dcache_release_state  <=4'h0; 
                     dcache_uncachedInFlight_0  <= dcache__uncachedInFlight_WIRE_0 ; 
                     dcache_s2_valid  <=1'h0; 
                     dcache_s2_probe  <=1'h0; 
                     dcache_lrscCount  <=7'h0; 
                     dcache_pstore2_valid  <=1'h0; 
                     dcache_pstore1_held  <=1'h0; 
                     dcache_counter  <=9'h0; 
                     dcache_grantInProgress  <=1'h0; 
                     dcache_blockProbeAfterGrantCount  <=3'h0; 
                     dcache_counter_1  <=9'h0; 
                     dcache_io_cpu_perf_acquire_counter  <=9'h0; 
                     dcache_io_cpu_perf_release_counter  <=9'h0; 
                     dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count  <=3'h0;
                 end 
              else 
                 begin  
                     dcache_s1_valid  <= dcache__io_cpu_req_ready_output & dcache_io_cpu_req_valid ;
                     if ( dcache__GEN_292 )
                         begin 
                             if ( dcache_metaArb_io_in_6_ready ) 
                                 dcache_s1_probe  <=1'h1;
                              else  
                                 dcache_s1_probe  <= dcache__GEN_87 ;
                         end 
                      else  
                         dcache_s1_probe  <= dcache__GEN_87 ; 
                     dcache_s1_tlb_req_valid  <= dcache__tlb_port_req_ready_output & dcache_tlb_port_req_valid ; 
                     dcache_s2_tlb_req_valid  <= dcache_s1_tlb_req_valid ;
                     if ( dcache__GEN_260 )
                         begin 
                             if ( dcache_grantIsCached )
                                 begin 
                                     if ( dcache_d_last )
                                         begin  
                                             dcache_cached_grant_wait  <=1'h0; 
                                             dcache_blockProbeAfterGrantCount  <=3'h7;
                                         end 
                                      else 
                                         begin 
                                             if ( dcache__GEN_248 )
                                                 begin 
                                                     if ( dcache_s2_uncached )
                                                         begin 
                                                         end 
                                                      else  
                                                         dcache_cached_grant_wait  <=1'h1;
                                                 end 
                                              else 
                                                 begin 
                                                 end 
                                             if ( dcache__GEN_256 ) 
                                                 dcache_blockProbeAfterGrantCount  <= dcache__GEN_257 [2:0];
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                     if ( dcache__GEN_248 )
                                         begin 
                                             if ( dcache_s2_uncached )
                                                 begin 
                                                     if ( dcache_a_sel ) 
                                                         dcache_uncachedInFlight_0  <=1'h1;
                                                      else 
                                                         begin 
                                                         end 
                                                 end 
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else 
                                         begin 
                                         end  
                                     dcache_grantInProgress  <= dcache__GEN_263 ;
                                 end 
                              else 
                                 begin 
                                     if ( dcache__GEN_248 )
                                         begin 
                                             if ( dcache_s2_uncached )
                                                 begin 
                                                 end 
                                              else  
                                                 dcache_cached_grant_wait  <=1'h1;
                                         end 
                                      else 
                                         begin 
                                         end 
                                     if ( dcache_grantIsUncached )
                                         begin 
                                             if ( dcache__GEN_266 ) 
                                                 dcache_uncachedInFlight_0  <=1'h0;
                                              else 
                                                 if ( dcache__GEN_248 )
                                                     begin 
                                                         if ( dcache_s2_uncached )
                                                             begin 
                                                                 if ( dcache_a_sel ) 
                                                                     dcache_uncachedInFlight_0  <=1'h1;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                             end 
                                                          else 
                                                             begin 
                                                             end 
                                                     end 
                                                  else 
                                                     begin 
                                                     end 
                                         end 
                                      else 
                                         if ( dcache__GEN_248 )
                                             begin 
                                                 if ( dcache_s2_uncached )
                                                     begin 
                                                         if ( dcache_a_sel ) 
                                                             dcache_uncachedInFlight_0  <=1'h1;
                                                          else 
                                                             begin 
                                                             end 
                                                     end 
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin 
                                             end 
                                     if ( dcache__GEN_256 ) 
                                         dcache_blockProbeAfterGrantCount  <= dcache__GEN_257 [2:0];
                                      else 
                                         begin 
                                         end 
                                 end 
                         end 
                      else 
                         begin 
                             if ( dcache__GEN_248 )
                                 begin 
                                     if ( dcache_s2_uncached )
                                         begin 
                                             if ( dcache_a_sel ) 
                                                 dcache_uncachedInFlight_0  <=1'h1;
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else  
                                         dcache_cached_grant_wait  <=1'h1;
                                 end 
                              else 
                                 begin 
                                 end 
                             if ( dcache__GEN_256 ) 
                                 dcache_blockProbeAfterGrantCount  <= dcache__GEN_257 [2:0];
                              else 
                                 begin 
                                 end 
                         end 
                     if ( dcache_resetting )
                         begin 
                             if ( dcache_flushDone ) 
                                 dcache_resetting  <=1'h0;
                              else 
                                 if ( dcache_REG ) 
                                     dcache_resetting  <=1'h1;
                                  else 
                                     begin 
                                     end 
                         end 
                      else 
                         if ( dcache_REG ) 
                             dcache_resetting  <=1'h1;
                          else 
                             begin 
                             end 
                     if ( dcache_resetting ) 
                         dcache_flushCounter  <= dcache_flushCounterNext [5:0];
                      else 
                         begin 
                         end 
                     if ( dcache__GEN_300 )
                         begin 
                             if ( dcache__GEN_302 ) 
                                 dcache_release_ack_wait  <=1'h1;
                              else 
                                 if ( dcache__GEN_260 )
                                     begin 
                                         if ( dcache_grantIsCached )
                                             begin 
                                             end 
                                          else 
                                             if ( dcache_grantIsUncached )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( dcache_grantIsVoluntary ) 
                                                     dcache_release_ack_wait  <=1'h0;
                                                  else 
                                                     begin 
                                                     end 
                                     end 
                                  else 
                                     begin 
                                     end 
                         end 
                      else 
                         if ( dcache__GEN_260 )
                             begin 
                                 if ( dcache_grantIsCached )
                                     begin 
                                     end 
                                  else 
                                     if ( dcache_grantIsUncached )
                                         begin 
                                         end 
                                      else 
                                         if ( dcache_grantIsVoluntary ) 
                                             dcache_release_ack_wait  <=1'h0;
                                          else 
                                             begin 
                                             end 
                             end 
                          else 
                             begin 
                             end 
                     if ( dcache__GEN_303 ) 
                         dcache_release_state  <=4'h0;
                      else 
                         if ( dcache__GEN_300 )
                             begin 
                                 if ( dcache_releaseDone ) 
                                     dcache_release_state  <=4'h6;
                                  else 
                                     if ( dcache__GEN_298 )
                                         begin 
                                             if ( dcache_releaseDone ) 
                                                 dcache_release_state  <=4'h7;
                                              else 
                                                 if ( dcache__GEN_296 )
                                                     begin 
                                                         if ( dcache_releaseDone ) 
                                                             dcache_release_state  <=4'h7;
                                                          else 
                                                             if ( dcache__GEN_294 )
                                                                 begin 
                                                                     if ( dcache_releaseDone ) 
                                                                         dcache_release_state  <=4'h0;
                                                                      else 
                                                                         if ( dcache__GEN_292 )
                                                                             begin 
                                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else 
                                                                                     if ( dcache_s2_probe )
                                                                                         begin 
                                                                                             if ( dcache_s2_meta_error ) 
                                                                                                 dcache_release_state  <=4'h4;
                                                                                              else 
                                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                                     dcache_release_state  <=4'h2;
                                                                                                  else 
                                                                                                     if ( dcache__GEN_290 )
                                                                                                         begin 
                                                                                                             if ( dcache_releaseDone ) 
                                                                                                                 dcache_release_state  <=4'h7;
                                                                                                              else  
                                                                                                                 dcache_release_state  <=4'h3;
                                                                                                         end 
                                                                                                      else 
                                                                                                         if ( dcache_releaseDone ) 
                                                                                                             dcache_release_state  <=4'h0;
                                                                                                          else  
                                                                                                             dcache_release_state  <=4'h5;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_s2_victimize ) 
                                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                                          else 
                                                                                             begin 
                                                                                             end 
                                                                             end 
                                                                          else 
                                                                             if ( dcache_s2_probe )
                                                                                 begin 
                                                                                     if ( dcache_s2_meta_error ) 
                                                                                         dcache_release_state  <=4'h4;
                                                                                      else 
                                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                                             dcache_release_state  <=4'h2;
                                                                                          else 
                                                                                             if ( dcache__GEN_290 )
                                                                                                 begin 
                                                                                                     if ( dcache_releaseDone ) 
                                                                                                         dcache_release_state  <=4'h7;
                                                                                                      else  
                                                                                                         dcache_release_state  <=4'h3;
                                                                                                 end 
                                                                                              else 
                                                                                                 if ( dcache_releaseDone ) 
                                                                                                     dcache_release_state  <=4'h0;
                                                                                                  else  
                                                                                                     dcache_release_state  <=4'h5;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_s2_victimize ) 
                                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                                  else 
                                                                                     begin 
                                                                                     end 
                                                                 end 
                                                              else 
                                                                 if ( dcache__GEN_292 )
                                                                     begin 
                                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else 
                                                                             if ( dcache_s2_probe )
                                                                                 begin 
                                                                                     if ( dcache_s2_meta_error ) 
                                                                                         dcache_release_state  <=4'h4;
                                                                                      else 
                                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                                             dcache_release_state  <=4'h2;
                                                                                          else 
                                                                                             if ( dcache__GEN_290 )
                                                                                                 begin 
                                                                                                     if ( dcache_releaseDone ) 
                                                                                                         dcache_release_state  <=4'h7;
                                                                                                      else  
                                                                                                         dcache_release_state  <=4'h3;
                                                                                                 end 
                                                                                              else 
                                                                                                 if ( dcache_releaseDone ) 
                                                                                                     dcache_release_state  <=4'h0;
                                                                                                  else  
                                                                                                     dcache_release_state  <=4'h5;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_s2_victimize ) 
                                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                                  else 
                                                                                     begin 
                                                                                     end 
                                                                     end 
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                     end 
                                                  else 
                                                     if ( dcache__GEN_294 )
                                                         begin 
                                                             if ( dcache_releaseDone ) 
                                                                 dcache_release_state  <=4'h0;
                                                              else 
                                                                 if ( dcache__GEN_292 )
                                                                     begin 
                                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else 
                                                                             if ( dcache_s2_probe )
                                                                                 begin 
                                                                                     if ( dcache_s2_meta_error ) 
                                                                                         dcache_release_state  <=4'h4;
                                                                                      else 
                                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                                             dcache_release_state  <=4'h2;
                                                                                          else 
                                                                                             if ( dcache__GEN_290 )
                                                                                                 begin 
                                                                                                     if ( dcache_releaseDone ) 
                                                                                                         dcache_release_state  <=4'h7;
                                                                                                      else  
                                                                                                         dcache_release_state  <=4'h3;
                                                                                                 end 
                                                                                              else 
                                                                                                 if ( dcache_releaseDone ) 
                                                                                                     dcache_release_state  <=4'h0;
                                                                                                  else  
                                                                                                     dcache_release_state  <=4'h5;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_s2_victimize ) 
                                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                                  else 
                                                                                     begin 
                                                                                     end 
                                                                     end 
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                         end 
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                         end 
                                      else 
                                         if ( dcache__GEN_296 )
                                             begin 
                                                 if ( dcache_releaseDone ) 
                                                     dcache_release_state  <=4'h7;
                                                  else 
                                                     if ( dcache__GEN_294 )
                                                         begin 
                                                             if ( dcache_releaseDone ) 
                                                                 dcache_release_state  <=4'h0;
                                                              else 
                                                                 if ( dcache__GEN_292 )
                                                                     begin 
                                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else 
                                                                             if ( dcache_s2_probe )
                                                                                 begin 
                                                                                     if ( dcache_s2_meta_error ) 
                                                                                         dcache_release_state  <=4'h4;
                                                                                      else 
                                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                                             dcache_release_state  <=4'h2;
                                                                                          else 
                                                                                             if ( dcache__GEN_290 )
                                                                                                 begin 
                                                                                                     if ( dcache_releaseDone ) 
                                                                                                         dcache_release_state  <=4'h7;
                                                                                                      else  
                                                                                                         dcache_release_state  <=4'h3;
                                                                                                 end 
                                                                                              else 
                                                                                                 if ( dcache_releaseDone ) 
                                                                                                     dcache_release_state  <=4'h0;
                                                                                                  else  
                                                                                                     dcache_release_state  <=4'h5;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_s2_victimize ) 
                                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                                  else 
                                                                                     begin 
                                                                                     end 
                                                                     end 
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                         end 
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                             end 
                                          else 
                                             if ( dcache__GEN_294 )
                                                 begin 
                                                     if ( dcache_releaseDone ) 
                                                         dcache_release_state  <=4'h0;
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                 end 
                                              else 
                                                 if ( dcache__GEN_292 )
                                                     begin 
                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                             dcache_release_state  <=4'h0;
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                     end 
                                                  else 
                                                     if ( dcache_s2_probe )
                                                         begin 
                                                             if ( dcache_s2_meta_error ) 
                                                                 dcache_release_state  <=4'h4;
                                                              else 
                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                     dcache_release_state  <=4'h2;
                                                                  else 
                                                                     if ( dcache__GEN_290 )
                                                                         begin 
                                                                             if ( dcache_releaseDone ) 
                                                                                 dcache_release_state  <=4'h7;
                                                                              else  
                                                                                 dcache_release_state  <=4'h3;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_releaseDone ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else  
                                                                             dcache_release_state  <=4'h5;
                                                         end 
                                                      else 
                                                         if ( dcache_s2_victimize ) 
                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                          else 
                                                             begin 
                                                             end 
                             end 
                          else 
                             if ( dcache__GEN_298 )
                                 begin 
                                     if ( dcache_releaseDone ) 
                                         dcache_release_state  <=4'h7;
                                      else 
                                         if ( dcache__GEN_296 )
                                             begin 
                                                 if ( dcache_releaseDone ) 
                                                     dcache_release_state  <=4'h7;
                                                  else 
                                                     if ( dcache__GEN_294 )
                                                         begin 
                                                             if ( dcache_releaseDone ) 
                                                                 dcache_release_state  <=4'h0;
                                                              else 
                                                                 if ( dcache__GEN_292 )
                                                                     begin 
                                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else 
                                                                             if ( dcache_s2_probe )
                                                                                 begin 
                                                                                     if ( dcache_s2_meta_error ) 
                                                                                         dcache_release_state  <=4'h4;
                                                                                      else 
                                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                                             dcache_release_state  <=4'h2;
                                                                                          else 
                                                                                             if ( dcache__GEN_290 )
                                                                                                 begin 
                                                                                                     if ( dcache_releaseDone ) 
                                                                                                         dcache_release_state  <=4'h7;
                                                                                                      else  
                                                                                                         dcache_release_state  <=4'h3;
                                                                                                 end 
                                                                                              else 
                                                                                                 if ( dcache_releaseDone ) 
                                                                                                     dcache_release_state  <=4'h0;
                                                                                                  else  
                                                                                                     dcache_release_state  <=4'h5;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_s2_victimize ) 
                                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                                  else 
                                                                                     begin 
                                                                                     end 
                                                                     end 
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                         end 
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                             end 
                                          else 
                                             if ( dcache__GEN_294 )
                                                 begin 
                                                     if ( dcache_releaseDone ) 
                                                         dcache_release_state  <=4'h0;
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                 end 
                                              else 
                                                 if ( dcache__GEN_292 )
                                                     begin 
                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                             dcache_release_state  <=4'h0;
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                     end 
                                                  else 
                                                     if ( dcache_s2_probe )
                                                         begin 
                                                             if ( dcache_s2_meta_error ) 
                                                                 dcache_release_state  <=4'h4;
                                                              else 
                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                     dcache_release_state  <=4'h2;
                                                                  else 
                                                                     if ( dcache__GEN_290 )
                                                                         begin 
                                                                             if ( dcache_releaseDone ) 
                                                                                 dcache_release_state  <=4'h7;
                                                                              else  
                                                                                 dcache_release_state  <=4'h3;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_releaseDone ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else  
                                                                             dcache_release_state  <=4'h5;
                                                         end 
                                                      else 
                                                         if ( dcache_s2_victimize ) 
                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                          else 
                                                             begin 
                                                             end 
                                 end 
                              else 
                                 if ( dcache__GEN_296 )
                                     begin 
                                         if ( dcache_releaseDone ) 
                                             dcache_release_state  <=4'h7;
                                          else 
                                             if ( dcache__GEN_294 )
                                                 begin 
                                                     if ( dcache_releaseDone ) 
                                                         dcache_release_state  <=4'h0;
                                                      else 
                                                         if ( dcache__GEN_292 )
                                                             begin 
                                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else 
                                                                     if ( dcache_s2_probe )
                                                                         begin 
                                                                             if ( dcache_s2_meta_error ) 
                                                                                 dcache_release_state  <=4'h4;
                                                                              else 
                                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                                     dcache_release_state  <=4'h2;
                                                                                  else 
                                                                                     if ( dcache__GEN_290 )
                                                                                         begin 
                                                                                             if ( dcache_releaseDone ) 
                                                                                                 dcache_release_state  <=4'h7;
                                                                                              else  
                                                                                                 dcache_release_state  <=4'h3;
                                                                                         end 
                                                                                      else 
                                                                                         if ( dcache_releaseDone ) 
                                                                                             dcache_release_state  <=4'h0;
                                                                                          else  
                                                                                             dcache_release_state  <=4'h5;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_s2_victimize ) 
                                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                                          else 
                                                                             begin 
                                                                             end 
                                                             end 
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                 end 
                                              else 
                                                 if ( dcache__GEN_292 )
                                                     begin 
                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                             dcache_release_state  <=4'h0;
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                     end 
                                                  else 
                                                     if ( dcache_s2_probe )
                                                         begin 
                                                             if ( dcache_s2_meta_error ) 
                                                                 dcache_release_state  <=4'h4;
                                                              else 
                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                     dcache_release_state  <=4'h2;
                                                                  else 
                                                                     if ( dcache__GEN_290 )
                                                                         begin 
                                                                             if ( dcache_releaseDone ) 
                                                                                 dcache_release_state  <=4'h7;
                                                                              else  
                                                                                 dcache_release_state  <=4'h3;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_releaseDone ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else  
                                                                             dcache_release_state  <=4'h5;
                                                         end 
                                                      else 
                                                         if ( dcache_s2_victimize ) 
                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                          else 
                                                             begin 
                                                             end 
                                     end 
                                  else 
                                     if ( dcache__GEN_294 )
                                         begin 
                                             if ( dcache_releaseDone ) 
                                                 dcache_release_state  <=4'h0;
                                              else 
                                                 if ( dcache__GEN_292 )
                                                     begin 
                                                         if ( dcache_metaArb_io_in_6_ready ) 
                                                             dcache_release_state  <=4'h0;
                                                          else 
                                                             if ( dcache_s2_probe )
                                                                 begin 
                                                                     if ( dcache_s2_meta_error ) 
                                                                         dcache_release_state  <=4'h4;
                                                                      else 
                                                                         if ( dcache_s2_prb_ack_data ) 
                                                                             dcache_release_state  <=4'h2;
                                                                          else 
                                                                             if ( dcache__GEN_290 )
                                                                                 begin 
                                                                                     if ( dcache_releaseDone ) 
                                                                                         dcache_release_state  <=4'h7;
                                                                                      else  
                                                                                         dcache_release_state  <=4'h3;
                                                                                 end 
                                                                              else 
                                                                                 if ( dcache_releaseDone ) 
                                                                                     dcache_release_state  <=4'h0;
                                                                                  else  
                                                                                     dcache_release_state  <=4'h5;
                                                                 end 
                                                              else 
                                                                 if ( dcache_s2_victimize ) 
                                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                                  else 
                                                                     begin 
                                                                     end 
                                                     end 
                                                  else 
                                                     if ( dcache_s2_probe )
                                                         begin 
                                                             if ( dcache_s2_meta_error ) 
                                                                 dcache_release_state  <=4'h4;
                                                              else 
                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                     dcache_release_state  <=4'h2;
                                                                  else 
                                                                     if ( dcache__GEN_290 )
                                                                         begin 
                                                                             if ( dcache_releaseDone ) 
                                                                                 dcache_release_state  <=4'h7;
                                                                              else  
                                                                                 dcache_release_state  <=4'h3;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_releaseDone ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else  
                                                                             dcache_release_state  <=4'h5;
                                                         end 
                                                      else 
                                                         if ( dcache_s2_victimize ) 
                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                          else 
                                                             begin 
                                                             end 
                                         end 
                                      else 
                                         if ( dcache__GEN_292 )
                                             begin 
                                                 if ( dcache_metaArb_io_in_6_ready ) 
                                                     dcache_release_state  <=4'h0;
                                                  else 
                                                     if ( dcache_s2_probe )
                                                         begin 
                                                             if ( dcache_s2_meta_error ) 
                                                                 dcache_release_state  <=4'h4;
                                                              else 
                                                                 if ( dcache_s2_prb_ack_data ) 
                                                                     dcache_release_state  <=4'h2;
                                                                  else 
                                                                     if ( dcache__GEN_290 )
                                                                         begin 
                                                                             if ( dcache_releaseDone ) 
                                                                                 dcache_release_state  <=4'h7;
                                                                              else  
                                                                                 dcache_release_state  <=4'h3;
                                                                         end 
                                                                      else 
                                                                         if ( dcache_releaseDone ) 
                                                                             dcache_release_state  <=4'h0;
                                                                          else  
                                                                             dcache_release_state  <=4'h5;
                                                         end 
                                                      else 
                                                         if ( dcache_s2_victimize ) 
                                                             dcache_release_state  <= dcache__GEN_287 ;
                                                          else 
                                                             begin 
                                                             end 
                                             end 
                                          else 
                                             if ( dcache_s2_probe )
                                                 begin 
                                                     if ( dcache_s2_meta_error ) 
                                                         dcache_release_state  <=4'h4;
                                                      else 
                                                         if ( dcache_s2_prb_ack_data ) 
                                                             dcache_release_state  <=4'h2;
                                                          else 
                                                             if ( dcache__GEN_290 )
                                                                 begin 
                                                                     if ( dcache_releaseDone ) 
                                                                         dcache_release_state  <=4'h7;
                                                                      else  
                                                                         dcache_release_state  <=4'h3;
                                                                 end 
                                                              else 
                                                                 if ( dcache_releaseDone ) 
                                                                     dcache_release_state  <=4'h0;
                                                                  else  
                                                                     dcache_release_state  <=4'h5;
                                                 end 
                                              else 
                                                 if ( dcache_s2_victimize ) 
                                                     dcache_release_state  <= dcache__GEN_287 ;
                                                  else 
                                                     begin 
                                                     end  
                     dcache_s2_valid  <= dcache_s1_valid_masked & dcache_s1_sfence ==1'h0; 
                     dcache_s2_probe  <= dcache_s1_probe ;
                     if ( dcache_s1_probe ) 
                         dcache_lrscCount  <=7'h0;
                      else 
                         if ( dcache__GEN_166 ) 
                             dcache_lrscCount  <=7'h3;
                          else 
                             if ( dcache__GEN_164 ) 
                                 dcache_lrscCount  <= dcache__GEN_165 [6:0];
                              else 
                                 if ( dcache__GEN_162 ) 
                                     dcache_lrscCount  <= dcache__GEN_163 ;
                                  else 
                                     begin 
                                     end  
                     dcache_pstore2_valid  <= dcache_pstore2_valid & dcache_pstore_drain ==1'h0| dcache_advance_pstore1 ; 
                     dcache_pstore1_held  <=( dcache_s2_valid_hit & dcache_s2_write & dcache_s2_sc_fail ==1'h0& dcache_io_cpu_s2_kill ==1'h0& dcache_s2_store_merge ==1'h0| dcache_pstore1_held )& dcache_pstore2_valid & dcache_pstore_drain ==1'h0;
                     if ( dcache__GEN_252 )
                         begin 
                             if ( dcache_d_first ) 
                                 dcache_counter  <= dcache_beats1 ;
                              else  
                                 dcache_counter  <= dcache_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( dcache__GEN_279 )
                         begin 
                             if ( dcache_c_first ) 
                                 dcache_counter_1  <= dcache_beats1_1 ;
                              else  
                                 dcache_counter_1  <= dcache_counter1_1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( dcache__GEN_308 )
                         begin 
                             if ( dcache_io_cpu_perf_acquire_first ) 
                                 dcache_io_cpu_perf_acquire_counter  <= dcache_io_cpu_perf_acquire_beats1 ;
                              else  
                                 dcache_io_cpu_perf_acquire_counter  <= dcache_io_cpu_perf_acquire_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( dcache__GEN_312 )
                         begin 
                             if ( dcache_io_cpu_perf_release_first ) 
                                 dcache_io_cpu_perf_release_counter  <= dcache_io_cpu_perf_release_beats1 ;
                              else  
                                 dcache_io_cpu_perf_release_counter  <= dcache_io_cpu_perf_release_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( dcache__GEN_316 ) 
                         dcache_io_cpu_perf_blocked_near_end_of_refill_refill_count  <= dcache__GEN_317 [2:0];
                      else 
                         begin 
                         end 
                 end 
         end
  assign  dcache_auto_out_a_valid = dcache_nodeOut_a_valid ; 
  assign  dcache_auto_out_a_bits_opcode = dcache_nodeOut_a_bits_opcode ; 
  assign  dcache_auto_out_a_bits_param = dcache_nodeOut_a_bits_param ; 
  assign  dcache_auto_out_a_bits_size = dcache_nodeOut_a_bits_size ; 
  assign  dcache_auto_out_a_bits_source = dcache_nodeOut_a_bits_source ; 
  assign  dcache_auto_out_a_bits_address = dcache_nodeOut_a_bits_address ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_bufferable = dcache_nodeOut_a_bits_user_amba_prot_bufferable ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_modifiable = dcache_nodeOut_a_bits_user_amba_prot_modifiable ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_readalloc = dcache_nodeOut_a_bits_user_amba_prot_readalloc ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_writealloc = dcache_nodeOut_a_bits_user_amba_prot_writealloc ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_privileged = dcache_nodeOut_a_bits_user_amba_prot_privileged ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_secure = dcache_nodeOut_a_bits_user_amba_prot_secure ; 
  assign  dcache_auto_out_a_bits_user_amba_prot_fetch = dcache_nodeOut_a_bits_user_amba_prot_fetch ; 
  assign  dcache_auto_out_a_bits_mask = dcache_nodeOut_a_bits_mask ; 
  assign  dcache_auto_out_a_bits_data = dcache_nodeOut_a_bits_data ; 
  assign  dcache_auto_out_a_bits_corrupt = dcache_nodeOut_a_bits_corrupt ; 
  assign  dcache_auto_out_b_ready = dcache_nodeOut_b_ready ; 
  assign  dcache_auto_out_c_valid = dcache_nodeOut_c_valid ; 
  assign  dcache_auto_out_c_bits_opcode = dcache_nodeOut_c_bits_opcode ; 
  assign  dcache_auto_out_c_bits_param = dcache_nodeOut_c_bits_param ; 
  assign  dcache_auto_out_c_bits_size = dcache_nodeOut_c_bits_size ; 
  assign  dcache_auto_out_c_bits_source = dcache_nodeOut_c_bits_source ; 
  assign  dcache_auto_out_c_bits_address = dcache_nodeOut_c_bits_address ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_bufferable = dcache_nodeOut_c_bits_user_amba_prot_bufferable ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_modifiable = dcache_nodeOut_c_bits_user_amba_prot_modifiable ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_readalloc = dcache_nodeOut_c_bits_user_amba_prot_readalloc ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_writealloc = dcache_nodeOut_c_bits_user_amba_prot_writealloc ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_privileged = dcache_nodeOut_c_bits_user_amba_prot_privileged ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_secure = dcache_nodeOut_c_bits_user_amba_prot_secure ; 
  assign  dcache_auto_out_c_bits_user_amba_prot_fetch = dcache_nodeOut_c_bits_user_amba_prot_fetch ; 
  assign  dcache_auto_out_c_bits_data = dcache_nodeOut_c_bits_data ; 
  assign  dcache_auto_out_c_bits_corrupt = dcache_nodeOut_c_bits_corrupt ; 
  assign  dcache_auto_out_d_ready = dcache_nodeOut_d_ready ; 
  assign  dcache_auto_out_e_valid = dcache_nodeOut_e_valid ; 
  assign  dcache_auto_out_e_bits_sink = dcache_nodeOut_e_bits_sink ; 
  assign  dcache_io_cpu_req_ready = dcache__io_cpu_req_ready_output ; 
  assign  dcache_io_cpu_s2_nack = dcache__io_cpu_s2_nack_output ; 
  assign  dcache_io_cpu_s2_nack_cause_raw = dcache_io_cpu_s2_nack_cause_raw_REG |( dcache_s2_waw_hazard ==1'h0| dcache_s2_store_merge )==1'h0; 
  assign  dcache_io_cpu_s2_uncached = dcache_s2_uncached & dcache_s2_hit ==1'h0; 
  assign  dcache_io_cpu_s2_paddr = dcache_s2_req_addr [31:0]; 
  assign  dcache_io_cpu_resp_valid =( dcache_s2_valid_hit_pre_data_ecc | dcache_doUncachedResp )& dcache_s2_data_error ==1'h0; 
  assign  dcache_io_cpu_resp_bits_addr = dcache_doUncachedResp  ?  dcache_s2_uncached_resp_addr : dcache_s2_req_addr ; 
  assign  dcache_io_cpu_resp_bits_tag = dcache_s2_req_tag ; 
  assign  dcache_io_cpu_resp_bits_cmd = dcache_s2_req_cmd ; 
  assign  dcache_io_cpu_resp_bits_size = dcache_s2_req_size ; 
  assign  dcache_io_cpu_resp_bits_signed = dcache_s2_req_signed ; 
  assign  dcache_io_cpu_resp_bits_dprv = dcache_s2_req_dprv ; 
  assign  dcache_io_cpu_resp_bits_dv = dcache_s2_req_dv ; 
  assign  dcache_io_cpu_resp_bits_data ={ dcache_size ==2'h0| dcache_io_cpu_resp_bits_data_doZero_2  ? ( dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_zeroed_2 [7] ? 56'hFFFFFFFFFFFFFF:56'h0): dcache__GEN_306 [63:8], dcache_io_cpu_resp_bits_data_zeroed_2 }|{63'h0, dcache_s2_sc_fail }; 
  assign  dcache_io_cpu_resp_bits_mask = dcache_s2_req_mask ; 
  assign  dcache_io_cpu_resp_bits_replay = dcache_doUncachedResp ; 
  assign  dcache_io_cpu_resp_bits_has_data = dcache_s2_read ; 
  assign  dcache_io_cpu_resp_bits_data_word_bypass ={ dcache_size ==2'h2| dcache_io_cpu_resp_bits_data_word_bypass_doZero  ? ( dcache_s2_req_signed & dcache_io_cpu_resp_bits_data_word_bypass_zeroed [31] ? 32'hFFFFFFFF:32'h0): dcache_s2_data_word_possibly_uncached [63:32], dcache_io_cpu_resp_bits_data_word_bypass_zeroed }; 
  assign  dcache_io_cpu_resp_bits_data_raw = dcache_s2_data_word ; 
  assign  dcache_io_cpu_resp_bits_store_data = dcache_pstore1_data ; 
  assign  dcache_io_cpu_replay_next = dcache__io_cpu_replay_next_output ; 
  assign  dcache_io_cpu_s2_xcpt_ma_ld = dcache__io_cpu_s2_xcpt_ma_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_ma_st = dcache__io_cpu_s2_xcpt_ma_st_output ; 
  assign  dcache_io_cpu_s2_xcpt_pf_ld = dcache__io_cpu_s2_xcpt_pf_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_pf_st = dcache__io_cpu_s2_xcpt_pf_st_output ; 
  assign  dcache_io_cpu_s2_xcpt_gf_ld = dcache__io_cpu_s2_xcpt_gf_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_gf_st = dcache__io_cpu_s2_xcpt_gf_st_output ; 
  assign  dcache_io_cpu_s2_xcpt_ae_ld = dcache__io_cpu_s2_xcpt_ae_ld_output ; 
  assign  dcache_io_cpu_s2_xcpt_ae_st = dcache__io_cpu_s2_xcpt_ae_st_output ; 
  assign  dcache_io_cpu_s2_gpa = dcache_s2_tlb_xcpt_gpa ; 
  assign  dcache_io_cpu_s2_gpa_is_pte = dcache_s2_tlb_xcpt_gpa_is_pte ; 
  assign  dcache_io_cpu_ordered =( dcache_s1_valid & dcache_s1_req_no_xcpt ==1'h0| dcache_s2_valid & dcache_s2_req_no_xcpt ==1'h0| dcache_cached_grant_wait |(| dcache_uncachedInFlight_0 ))==1'h0; 
  assign  dcache_io_cpu_perf_acquire = dcache_io_cpu_perf_acquire_done ; 
  assign  dcache_io_cpu_perf_release = dcache_io_cpu_perf_release_done ; 
  assign  dcache_io_cpu_perf_grant = dcache_nodeOut_d_valid & dcache_d_last ; 
  assign  dcache_io_cpu_perf_tlbMiss = dcache_io_ptw_req_ready & dcache__io_ptw_req_valid_output ; 
  assign  dcache_io_cpu_perf_blocked = dcache_cached_grant_wait & dcache_io_cpu_perf_blocked_near_end_of_refill ==1'h0; 
  assign  dcache_io_cpu_perf_canAcceptStoreThenLoad = dcache__io_cpu_perf_canAcceptStoreThenLoad_output ; 
  assign  dcache_io_cpu_perf_canAcceptStoreThenRMW = dcache__io_cpu_perf_canAcceptStoreThenLoad_output & dcache_pstore2_valid ==1'h0; 
  assign  dcache_io_cpu_perf_canAcceptLoadThenLoad =( dcache_s1_valid & dcache_s1_write &( dcache_s1_req_cmd ==5'h0| dcache_s1_req_cmd ==5'h10| dcache_s1_req_cmd ==5'h6| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF|( dcache_s1_req_cmd ==5'h1| dcache_s1_req_cmd ==5'h11| dcache_s1_req_cmd ==5'h7| dcache_s1_req_cmd ==5'h4| dcache_s1_req_cmd ==5'h9| dcache_s1_req_cmd ==5'hA| dcache_s1_req_cmd ==5'hB| dcache_s1_req_cmd ==5'h8| dcache_s1_req_cmd ==5'hC| dcache_s1_req_cmd ==5'hD| dcache_s1_req_cmd ==5'hE| dcache_s1_req_cmd ==5'hF)&( dcache_s1_req_cmd ==5'h11| dcache_s1_req_size <2'h0))&( dcache_s2_valid & dcache_s2_write & dcache_s2_waw_hazard ==1'h0| dcache_pstore1_held | dcache_pstore2_valid ))==1'h0; 
  assign  dcache_io_cpu_perf_storeBufferEmptyAfterLoad =( dcache_s1_valid & dcache_s1_write | dcache_s2_valid & dcache_s2_write & dcache_s2_waw_hazard ==1'h0| dcache_pstore1_held | dcache_pstore2_valid )==1'h0; 
  assign  dcache_io_cpu_perf_storeBufferEmptyAfterStore =( dcache_s1_valid & dcache_s1_write | dcache_s2_valid & dcache_s2_write & dcache_pstore1_rmw |( dcache_s2_valid & dcache_s2_write & dcache_s2_waw_hazard ==1'h0| dcache_pstore1_held )& dcache_pstore2_valid )==1'h0; 
  assign  dcache_io_cpu_clock_enabled = dcache_clock_en_reg ; 
  assign  dcache_io_ptw_req_valid = dcache__io_ptw_req_valid_output ; 
  assign  dcache_io_ptw_req_bits_valid = dcache_tlb_io_ptw_req_bits_valid ; 
  assign  dcache_io_ptw_req_bits_bits_addr = dcache_tlb_io_ptw_req_bits_bits_addr ; 
  assign  dcache_io_ptw_req_bits_bits_need_gpa = dcache_tlb_io_ptw_req_bits_bits_need_gpa ; 
  assign  dcache_io_ptw_req_bits_bits_vstage1 = dcache_tlb_io_ptw_req_bits_bits_vstage1 ; 
  assign  dcache_io_ptw_req_bits_bits_stage2 = dcache_tlb_io_ptw_req_bits_bits_stage2 ; 
  assign  dcache_io_ptw_customCSRs_csrs_0_stall = dcache_tlb_io_ptw_customCSRs_csrs_0_stall ; 
  assign  dcache_io_ptw_customCSRs_csrs_0_set = dcache_tlb_io_ptw_customCSRs_csrs_0_set ; 
  assign  dcache_io_ptw_customCSRs_csrs_0_sdata = dcache_tlb_io_ptw_customCSRs_csrs_0_sdata ; 
  assign  dcache_io_ptw_customCSRs_csrs_1_stall = dcache_tlb_io_ptw_customCSRs_csrs_1_stall ; 
  assign  dcache_io_ptw_customCSRs_csrs_1_set = dcache_tlb_io_ptw_customCSRs_csrs_1_set ; 
  assign  dcache_io_ptw_customCSRs_csrs_1_sdata = dcache_tlb_io_ptw_customCSRs_csrs_1_sdata ; 
  assign  dcache_io_ptw_customCSRs_csrs_2_stall = dcache_tlb_io_ptw_customCSRs_csrs_2_stall ; 
  assign  dcache_io_ptw_customCSRs_csrs_2_set = dcache_tlb_io_ptw_customCSRs_csrs_2_set ; 
  assign  dcache_io_ptw_customCSRs_csrs_2_sdata = dcache_tlb_io_ptw_customCSRs_csrs_2_sdata ; 
  assign  dcache_io_ptw_customCSRs_csrs_3_stall = dcache_tlb_io_ptw_customCSRs_csrs_3_stall ; 
  assign  dcache_io_ptw_customCSRs_csrs_3_set = dcache_tlb_io_ptw_customCSRs_csrs_3_set ; 
  assign  dcache_io_ptw_customCSRs_csrs_3_sdata = dcache_tlb_io_ptw_customCSRs_csrs_3_sdata ; 
  assign  dcache_io_errors_bus_valid = dcache__io_errors_bus_valid_output ; 
  assign  dcache_io_errors_bus_bits = dcache__GEN_318 [31:0]; 
  assign  dcache_tlb_port_req_ready = dcache__tlb_port_req_ready_output ; 
  assign  dcache_tlb_port_s1_resp_miss = dcache_tlb_io_resp_miss ; 
  assign  dcache_tlb_port_s1_resp_paddr = dcache_tlb_io_resp_paddr ; 
  assign  dcache_tlb_port_s1_resp_gpa = dcache_tlb_io_resp_gpa ; 
  assign  dcache_tlb_port_s1_resp_gpa_is_pte = dcache_tlb_io_resp_gpa_is_pte ; 
  assign  dcache_tlb_port_s1_resp_pf_ld = dcache_tlb_io_resp_pf_ld ; 
  assign  dcache_tlb_port_s1_resp_pf_st = dcache_tlb_io_resp_pf_st ; 
  assign  dcache_tlb_port_s1_resp_pf_inst = dcache_tlb_io_resp_pf_inst ; 
  assign  dcache_tlb_port_s1_resp_gf_ld = dcache_tlb_io_resp_gf_ld ; 
  assign  dcache_tlb_port_s1_resp_gf_st = dcache_tlb_io_resp_gf_st ; 
  assign  dcache_tlb_port_s1_resp_gf_inst = dcache_tlb_io_resp_gf_inst ; 
  assign  dcache_tlb_port_s1_resp_ae_ld = dcache_tlb_io_resp_ae_ld ; 
  assign  dcache_tlb_port_s1_resp_ae_st = dcache_tlb_io_resp_ae_st ; 
  assign  dcache_tlb_port_s1_resp_ae_inst = dcache_tlb_io_resp_ae_inst ; 
  assign  dcache_tlb_port_s1_resp_ma_ld = dcache_tlb_io_resp_ma_ld ; 
  assign  dcache_tlb_port_s1_resp_ma_st = dcache_tlb_io_resp_ma_st ; 
  assign  dcache_tlb_port_s1_resp_ma_inst = dcache_tlb_io_resp_ma_inst ; 
  assign  dcache_tlb_port_s1_resp_cacheable = dcache_tlb_io_resp_cacheable ; 
  assign  dcache_tlb_port_s1_resp_must_alloc = dcache_tlb_io_resp_must_alloc ; 
  assign  dcache_tlb_port_s1_resp_prefetchable = dcache_tlb_io_resp_prefetchable ;
    assign dcache_clock = clock;
    assign dcache_reset = reset;
    assign dcache_auto_out_a_ready = widget_auto_in_a_ready;
    assign widget_auto_in_a_valid = dcache_auto_out_a_valid;
    assign widget_auto_in_a_bits_opcode = dcache_auto_out_a_bits_opcode;
    assign widget_auto_in_a_bits_param = dcache_auto_out_a_bits_param;
    assign widget_auto_in_a_bits_size = dcache_auto_out_a_bits_size;
    assign widget_auto_in_a_bits_source = dcache_auto_out_a_bits_source;
    assign widget_auto_in_a_bits_address = dcache_auto_out_a_bits_address;
    assign widget_auto_in_a_bits_user_amba_prot_bufferable = dcache_auto_out_a_bits_user_amba_prot_bufferable;
    assign widget_auto_in_a_bits_user_amba_prot_modifiable = dcache_auto_out_a_bits_user_amba_prot_modifiable;
    assign widget_auto_in_a_bits_user_amba_prot_readalloc = dcache_auto_out_a_bits_user_amba_prot_readalloc;
    assign widget_auto_in_a_bits_user_amba_prot_writealloc = dcache_auto_out_a_bits_user_amba_prot_writealloc;
    assign widget_auto_in_a_bits_user_amba_prot_privileged = dcache_auto_out_a_bits_user_amba_prot_privileged;
    assign widget_auto_in_a_bits_user_amba_prot_secure = dcache_auto_out_a_bits_user_amba_prot_secure;
    assign widget_auto_in_a_bits_user_amba_prot_fetch = dcache_auto_out_a_bits_user_amba_prot_fetch;
    assign widget_auto_in_a_bits_mask = dcache_auto_out_a_bits_mask;
    assign widget_auto_in_a_bits_data = dcache_auto_out_a_bits_data;
    assign widget_auto_in_a_bits_corrupt = dcache_auto_out_a_bits_corrupt;
    assign widget_auto_in_b_ready = dcache_auto_out_b_ready;
    assign dcache_auto_out_b_valid = widget_auto_in_b_valid;
    assign dcache_auto_out_b_bits_opcode = widget_auto_in_b_bits_opcode;
    assign dcache_auto_out_b_bits_param = widget_auto_in_b_bits_param;
    assign dcache_auto_out_b_bits_size = widget_auto_in_b_bits_size;
    assign dcache_auto_out_b_bits_source = widget_auto_in_b_bits_source;
    assign dcache_auto_out_b_bits_address = widget_auto_in_b_bits_address;
    assign dcache_auto_out_b_bits_mask = widget_auto_in_b_bits_mask;
    assign dcache_auto_out_b_bits_data = widget_auto_in_b_bits_data;
    assign dcache_auto_out_b_bits_corrupt = widget_auto_in_b_bits_corrupt;
    assign dcache_auto_out_c_ready = widget_auto_in_c_ready;
    assign widget_auto_in_c_valid = dcache_auto_out_c_valid;
    assign widget_auto_in_c_bits_opcode = dcache_auto_out_c_bits_opcode;
    assign widget_auto_in_c_bits_param = dcache_auto_out_c_bits_param;
    assign widget_auto_in_c_bits_size = dcache_auto_out_c_bits_size;
    assign widget_auto_in_c_bits_source = dcache_auto_out_c_bits_source;
    assign widget_auto_in_c_bits_address = dcache_auto_out_c_bits_address;
    assign widget_auto_in_c_bits_user_amba_prot_bufferable = dcache_auto_out_c_bits_user_amba_prot_bufferable;
    assign widget_auto_in_c_bits_user_amba_prot_modifiable = dcache_auto_out_c_bits_user_amba_prot_modifiable;
    assign widget_auto_in_c_bits_user_amba_prot_readalloc = dcache_auto_out_c_bits_user_amba_prot_readalloc;
    assign widget_auto_in_c_bits_user_amba_prot_writealloc = dcache_auto_out_c_bits_user_amba_prot_writealloc;
    assign widget_auto_in_c_bits_user_amba_prot_privileged = dcache_auto_out_c_bits_user_amba_prot_privileged;
    assign widget_auto_in_c_bits_user_amba_prot_secure = dcache_auto_out_c_bits_user_amba_prot_secure;
    assign widget_auto_in_c_bits_user_amba_prot_fetch = dcache_auto_out_c_bits_user_amba_prot_fetch;
    assign widget_auto_in_c_bits_data = dcache_auto_out_c_bits_data;
    assign widget_auto_in_c_bits_corrupt = dcache_auto_out_c_bits_corrupt;
    assign widget_auto_in_d_ready = dcache_auto_out_d_ready;
    assign dcache_auto_out_d_valid = widget_auto_in_d_valid;
    assign dcache_auto_out_d_bits_opcode = widget_auto_in_d_bits_opcode;
    assign dcache_auto_out_d_bits_param = widget_auto_in_d_bits_param;
    assign dcache_auto_out_d_bits_size = widget_auto_in_d_bits_size;
    assign dcache_auto_out_d_bits_source = widget_auto_in_d_bits_source;
    assign dcache_auto_out_d_bits_sink = widget_auto_in_d_bits_sink;
    assign dcache_auto_out_d_bits_denied = widget_auto_in_d_bits_denied;
    assign dcache_auto_out_d_bits_data = widget_auto_in_d_bits_data;
    assign dcache_auto_out_d_bits_corrupt = widget_auto_in_d_bits_corrupt;
    assign dcache_auto_out_e_ready = widget_auto_in_e_ready;
    assign widget_auto_in_e_valid = dcache_auto_out_e_valid;
    assign widget_auto_in_e_bits_sink = dcache_auto_out_e_bits_sink;
    assign _dcache_io_cpu_req_ready = dcache_io_cpu_req_ready;
    assign dcache_io_cpu_req_valid = _dcacheArb_io_mem_req_valid;
    assign dcache_io_cpu_req_bits_addr = _dcacheArb_io_mem_req_bits_addr;
    assign dcache_io_cpu_req_bits_tag = _dcacheArb_io_mem_req_bits_tag;
    assign dcache_io_cpu_req_bits_cmd = _dcacheArb_io_mem_req_bits_cmd;
    assign dcache_io_cpu_req_bits_size = _dcacheArb_io_mem_req_bits_size;
    assign dcache_io_cpu_req_bits_signed = _dcacheArb_io_mem_req_bits_signed;
    assign dcache_io_cpu_req_bits_dprv = _dcacheArb_io_mem_req_bits_dprv;
    assign dcache_io_cpu_req_bits_dv = _dcacheArb_io_mem_req_bits_dv;
    assign dcache_io_cpu_req_bits_phys = _dcacheArb_io_mem_req_bits_phys;
    assign dcache_io_cpu_req_bits_no_alloc = _dcacheArb_io_mem_req_bits_no_alloc;
    assign dcache_io_cpu_req_bits_no_xcpt = _dcacheArb_io_mem_req_bits_no_xcpt;
    assign dcache_io_cpu_req_bits_data = _dcacheArb_io_mem_req_bits_data;
    assign dcache_io_cpu_req_bits_mask = _dcacheArb_io_mem_req_bits_mask;
    assign dcache_io_cpu_s1_kill = _dcacheArb_io_mem_s1_kill;
    assign dcache_io_cpu_s1_data_data = _dcacheArb_io_mem_s1_data_data;
    assign dcache_io_cpu_s1_data_mask = _dcacheArb_io_mem_s1_data_mask;
    assign _dcache_io_cpu_s2_nack = dcache_io_cpu_s2_nack;
    assign _dcache_io_cpu_s2_nack_cause_raw = dcache_io_cpu_s2_nack_cause_raw;
    assign dcache_io_cpu_s2_kill = _dcacheArb_io_mem_s2_kill;
    assign _dcache_io_cpu_s2_uncached = dcache_io_cpu_s2_uncached;
    assign _dcache_io_cpu_s2_paddr = dcache_io_cpu_s2_paddr;
    assign _dcache_io_cpu_resp_valid = dcache_io_cpu_resp_valid;
    assign _dcache_io_cpu_resp_bits_addr = dcache_io_cpu_resp_bits_addr;
    assign _dcache_io_cpu_resp_bits_tag = dcache_io_cpu_resp_bits_tag;
    assign _dcache_io_cpu_resp_bits_cmd = dcache_io_cpu_resp_bits_cmd;
    assign _dcache_io_cpu_resp_bits_size = dcache_io_cpu_resp_bits_size;
    assign _dcache_io_cpu_resp_bits_signed = dcache_io_cpu_resp_bits_signed;
    assign _dcache_io_cpu_resp_bits_dprv = dcache_io_cpu_resp_bits_dprv;
    assign _dcache_io_cpu_resp_bits_dv = dcache_io_cpu_resp_bits_dv;
    assign _dcache_io_cpu_resp_bits_data = dcache_io_cpu_resp_bits_data;
    assign _dcache_io_cpu_resp_bits_mask = dcache_io_cpu_resp_bits_mask;
    assign _dcache_io_cpu_resp_bits_replay = dcache_io_cpu_resp_bits_replay;
    assign _dcache_io_cpu_resp_bits_has_data = dcache_io_cpu_resp_bits_has_data;
    assign _dcache_io_cpu_resp_bits_data_word_bypass = dcache_io_cpu_resp_bits_data_word_bypass;
    assign _dcache_io_cpu_resp_bits_data_raw = dcache_io_cpu_resp_bits_data_raw;
    assign _dcache_io_cpu_resp_bits_store_data = dcache_io_cpu_resp_bits_store_data;
    assign _dcache_io_cpu_replay_next = dcache_io_cpu_replay_next;
    assign _dcache_io_cpu_s2_xcpt_ma_ld = dcache_io_cpu_s2_xcpt_ma_ld;
    assign _dcache_io_cpu_s2_xcpt_ma_st = dcache_io_cpu_s2_xcpt_ma_st;
    assign _dcache_io_cpu_s2_xcpt_pf_ld = dcache_io_cpu_s2_xcpt_pf_ld;
    assign _dcache_io_cpu_s2_xcpt_pf_st = dcache_io_cpu_s2_xcpt_pf_st;
    assign _dcache_io_cpu_s2_xcpt_gf_ld = dcache_io_cpu_s2_xcpt_gf_ld;
    assign _dcache_io_cpu_s2_xcpt_gf_st = dcache_io_cpu_s2_xcpt_gf_st;
    assign _dcache_io_cpu_s2_xcpt_ae_ld = dcache_io_cpu_s2_xcpt_ae_ld;
    assign _dcache_io_cpu_s2_xcpt_ae_st = dcache_io_cpu_s2_xcpt_ae_st;
    assign _dcache_io_cpu_s2_gpa = dcache_io_cpu_s2_gpa;
    assign _dcache_io_cpu_s2_gpa_is_pte = dcache_io_cpu_s2_gpa_is_pte;
    assign _dcache_io_cpu_ordered = dcache_io_cpu_ordered;
    assign _dcache_io_cpu_perf_acquire = dcache_io_cpu_perf_acquire;
    assign _dcache_io_cpu_perf_release = dcache_io_cpu_perf_release;
    assign _dcache_io_cpu_perf_grant = dcache_io_cpu_perf_grant;
    assign _dcache_io_cpu_perf_tlbMiss = dcache_io_cpu_perf_tlbMiss;
    assign _dcache_io_cpu_perf_blocked = dcache_io_cpu_perf_blocked;
    assign _dcache_io_cpu_perf_canAcceptStoreThenLoad = dcache_io_cpu_perf_canAcceptStoreThenLoad;
    assign _dcache_io_cpu_perf_canAcceptStoreThenRMW = dcache_io_cpu_perf_canAcceptStoreThenRMW;
    assign _dcache_io_cpu_perf_canAcceptLoadThenLoad = dcache_io_cpu_perf_canAcceptLoadThenLoad;
    assign _dcache_io_cpu_perf_storeBufferEmptyAfterLoad = dcache_io_cpu_perf_storeBufferEmptyAfterLoad;
    assign _dcache_io_cpu_perf_storeBufferEmptyAfterStore = dcache_io_cpu_perf_storeBufferEmptyAfterStore;
    assign dcache_io_cpu_keep_clock_enabled = _dcacheArb_io_mem_keep_clock_enabled;
    assign _dcache_io_cpu_clock_enabled = dcache_io_cpu_clock_enabled;
    assign dcache_io_ptw_req_ready = _ptw_io_requestor_0_req_ready;
    assign _dcache_io_ptw_req_valid = dcache_io_ptw_req_valid;
    assign _dcache_io_ptw_req_bits_valid = dcache_io_ptw_req_bits_valid;
    assign _dcache_io_ptw_req_bits_bits_addr = dcache_io_ptw_req_bits_bits_addr;
    assign _dcache_io_ptw_req_bits_bits_need_gpa = dcache_io_ptw_req_bits_bits_need_gpa;
    assign _dcache_io_ptw_req_bits_bits_vstage1 = dcache_io_ptw_req_bits_bits_vstage1;
    assign _dcache_io_ptw_req_bits_bits_stage2 = dcache_io_ptw_req_bits_bits_stage2;
    assign dcache_io_ptw_resp_valid = _ptw_io_requestor_0_resp_valid;
    assign dcache_io_ptw_resp_bits_ae_ptw = _ptw_io_requestor_0_resp_bits_ae_ptw;
    assign dcache_io_ptw_resp_bits_ae_final = _ptw_io_requestor_0_resp_bits_ae_final;
    assign dcache_io_ptw_resp_bits_pf = _ptw_io_requestor_0_resp_bits_pf;
    assign dcache_io_ptw_resp_bits_gf = _ptw_io_requestor_0_resp_bits_gf;
    assign dcache_io_ptw_resp_bits_hr = _ptw_io_requestor_0_resp_bits_hr;
    assign dcache_io_ptw_resp_bits_hw = _ptw_io_requestor_0_resp_bits_hw;
    assign dcache_io_ptw_resp_bits_hx = _ptw_io_requestor_0_resp_bits_hx;
    assign dcache_io_ptw_resp_bits_pte_reserved_for_future = _ptw_io_requestor_0_resp_bits_pte_reserved_for_future;
    assign dcache_io_ptw_resp_bits_pte_ppn = _ptw_io_requestor_0_resp_bits_pte_ppn;
    assign dcache_io_ptw_resp_bits_pte_reserved_for_software = _ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
    assign dcache_io_ptw_resp_bits_pte_d = _ptw_io_requestor_0_resp_bits_pte_d;
    assign dcache_io_ptw_resp_bits_pte_a = _ptw_io_requestor_0_resp_bits_pte_a;
    assign dcache_io_ptw_resp_bits_pte_g = _ptw_io_requestor_0_resp_bits_pte_g;
    assign dcache_io_ptw_resp_bits_pte_u = _ptw_io_requestor_0_resp_bits_pte_u;
    assign dcache_io_ptw_resp_bits_pte_x = _ptw_io_requestor_0_resp_bits_pte_x;
    assign dcache_io_ptw_resp_bits_pte_w = _ptw_io_requestor_0_resp_bits_pte_w;
    assign dcache_io_ptw_resp_bits_pte_r = _ptw_io_requestor_0_resp_bits_pte_r;
    assign dcache_io_ptw_resp_bits_pte_v = _ptw_io_requestor_0_resp_bits_pte_v;
    assign dcache_io_ptw_resp_bits_level = _ptw_io_requestor_0_resp_bits_level;
    assign dcache_io_ptw_resp_bits_fragmented_superpage = _ptw_io_requestor_0_resp_bits_fragmented_superpage;
    assign dcache_io_ptw_resp_bits_homogeneous = _ptw_io_requestor_0_resp_bits_homogeneous;
    assign dcache_io_ptw_resp_bits_gpa_valid = _ptw_io_requestor_0_resp_bits_gpa_valid;
    assign dcache_io_ptw_resp_bits_gpa_bits = _ptw_io_requestor_0_resp_bits_gpa_bits;
    assign dcache_io_ptw_resp_bits_gpa_is_pte = _ptw_io_requestor_0_resp_bits_gpa_is_pte;
    assign dcache_io_ptw_ptbr_mode = _ptw_io_requestor_0_ptbr_mode;
    assign dcache_io_ptw_ptbr_asid = _ptw_io_requestor_0_ptbr_asid;
    assign dcache_io_ptw_ptbr_ppn = _ptw_io_requestor_0_ptbr_ppn;
    assign dcache_io_ptw_hgatp_mode = _ptw_io_requestor_0_hgatp_mode;
    assign dcache_io_ptw_hgatp_asid = _ptw_io_requestor_0_hgatp_asid;
    assign dcache_io_ptw_hgatp_ppn = _ptw_io_requestor_0_hgatp_ppn;
    assign dcache_io_ptw_vsatp_mode = _ptw_io_requestor_0_vsatp_mode;
    assign dcache_io_ptw_vsatp_asid = _ptw_io_requestor_0_vsatp_asid;
    assign dcache_io_ptw_vsatp_ppn = _ptw_io_requestor_0_vsatp_ppn;
    assign dcache_io_ptw_status_debug = _ptw_io_requestor_0_status_debug;
    assign dcache_io_ptw_status_cease = _ptw_io_requestor_0_status_cease;
    assign dcache_io_ptw_status_wfi = _ptw_io_requestor_0_status_wfi;
    assign dcache_io_ptw_status_isa = _ptw_io_requestor_0_status_isa;
    assign dcache_io_ptw_status_dprv = _ptw_io_requestor_0_status_dprv;
    assign dcache_io_ptw_status_dv = _ptw_io_requestor_0_status_dv;
    assign dcache_io_ptw_status_prv = _ptw_io_requestor_0_status_prv;
    assign dcache_io_ptw_status_v = _ptw_io_requestor_0_status_v;
    assign dcache_io_ptw_status_sd = _ptw_io_requestor_0_status_sd;
    assign dcache_io_ptw_status_zero2 = _ptw_io_requestor_0_status_zero2;
    assign dcache_io_ptw_status_mpv = _ptw_io_requestor_0_status_mpv;
    assign dcache_io_ptw_status_gva = _ptw_io_requestor_0_status_gva;
    assign dcache_io_ptw_status_mbe = _ptw_io_requestor_0_status_mbe;
    assign dcache_io_ptw_status_sbe = _ptw_io_requestor_0_status_sbe;
    assign dcache_io_ptw_status_sxl = _ptw_io_requestor_0_status_sxl;
    assign dcache_io_ptw_status_uxl = _ptw_io_requestor_0_status_uxl;
    assign dcache_io_ptw_status_sd_rv32 = _ptw_io_requestor_0_status_sd_rv32;
    assign dcache_io_ptw_status_zero1 = _ptw_io_requestor_0_status_zero1;
    assign dcache_io_ptw_status_tsr = _ptw_io_requestor_0_status_tsr;
    assign dcache_io_ptw_status_tw = _ptw_io_requestor_0_status_tw;
    assign dcache_io_ptw_status_tvm = _ptw_io_requestor_0_status_tvm;
    assign dcache_io_ptw_status_mxr = _ptw_io_requestor_0_status_mxr;
    assign dcache_io_ptw_status_sum = _ptw_io_requestor_0_status_sum;
    assign dcache_io_ptw_status_mprv = _ptw_io_requestor_0_status_mprv;
    assign dcache_io_ptw_status_xs = _ptw_io_requestor_0_status_xs;
    assign dcache_io_ptw_status_fs = _ptw_io_requestor_0_status_fs;
    assign dcache_io_ptw_status_mpp = _ptw_io_requestor_0_status_mpp;
    assign dcache_io_ptw_status_vs = _ptw_io_requestor_0_status_vs;
    assign dcache_io_ptw_status_spp = _ptw_io_requestor_0_status_spp;
    assign dcache_io_ptw_status_mpie = _ptw_io_requestor_0_status_mpie;
    assign dcache_io_ptw_status_ube = _ptw_io_requestor_0_status_ube;
    assign dcache_io_ptw_status_spie = _ptw_io_requestor_0_status_spie;
    assign dcache_io_ptw_status_upie = _ptw_io_requestor_0_status_upie;
    assign dcache_io_ptw_status_mie = _ptw_io_requestor_0_status_mie;
    assign dcache_io_ptw_status_hie = _ptw_io_requestor_0_status_hie;
    assign dcache_io_ptw_status_sie = _ptw_io_requestor_0_status_sie;
    assign dcache_io_ptw_status_uie = _ptw_io_requestor_0_status_uie;
    assign dcache_io_ptw_hstatus_zero6 = _ptw_io_requestor_0_hstatus_zero6;
    assign dcache_io_ptw_hstatus_vsxl = _ptw_io_requestor_0_hstatus_vsxl;
    assign dcache_io_ptw_hstatus_zero5 = _ptw_io_requestor_0_hstatus_zero5;
    assign dcache_io_ptw_hstatus_vtsr = _ptw_io_requestor_0_hstatus_vtsr;
    assign dcache_io_ptw_hstatus_vtw = _ptw_io_requestor_0_hstatus_vtw;
    assign dcache_io_ptw_hstatus_vtvm = _ptw_io_requestor_0_hstatus_vtvm;
    assign dcache_io_ptw_hstatus_zero3 = _ptw_io_requestor_0_hstatus_zero3;
    assign dcache_io_ptw_hstatus_vgein = _ptw_io_requestor_0_hstatus_vgein;
    assign dcache_io_ptw_hstatus_zero2 = _ptw_io_requestor_0_hstatus_zero2;
    assign dcache_io_ptw_hstatus_hu = _ptw_io_requestor_0_hstatus_hu;
    assign dcache_io_ptw_hstatus_spvp = _ptw_io_requestor_0_hstatus_spvp;
    assign dcache_io_ptw_hstatus_spv = _ptw_io_requestor_0_hstatus_spv;
    assign dcache_io_ptw_hstatus_gva = _ptw_io_requestor_0_hstatus_gva;
    assign dcache_io_ptw_hstatus_vsbe = _ptw_io_requestor_0_hstatus_vsbe;
    assign dcache_io_ptw_hstatus_zero1 = _ptw_io_requestor_0_hstatus_zero1;
    assign dcache_io_ptw_gstatus_debug = _ptw_io_requestor_0_gstatus_debug;
    assign dcache_io_ptw_gstatus_cease = _ptw_io_requestor_0_gstatus_cease;
    assign dcache_io_ptw_gstatus_wfi = _ptw_io_requestor_0_gstatus_wfi;
    assign dcache_io_ptw_gstatus_isa = _ptw_io_requestor_0_gstatus_isa;
    assign dcache_io_ptw_gstatus_dprv = _ptw_io_requestor_0_gstatus_dprv;
    assign dcache_io_ptw_gstatus_dv = _ptw_io_requestor_0_gstatus_dv;
    assign dcache_io_ptw_gstatus_prv = _ptw_io_requestor_0_gstatus_prv;
    assign dcache_io_ptw_gstatus_v = _ptw_io_requestor_0_gstatus_v;
    assign dcache_io_ptw_gstatus_sd = _ptw_io_requestor_0_gstatus_sd;
    assign dcache_io_ptw_gstatus_zero2 = _ptw_io_requestor_0_gstatus_zero2;
    assign dcache_io_ptw_gstatus_mpv = _ptw_io_requestor_0_gstatus_mpv;
    assign dcache_io_ptw_gstatus_gva = _ptw_io_requestor_0_gstatus_gva;
    assign dcache_io_ptw_gstatus_mbe = _ptw_io_requestor_0_gstatus_mbe;
    assign dcache_io_ptw_gstatus_sbe = _ptw_io_requestor_0_gstatus_sbe;
    assign dcache_io_ptw_gstatus_sxl = _ptw_io_requestor_0_gstatus_sxl;
    assign dcache_io_ptw_gstatus_uxl = _ptw_io_requestor_0_gstatus_uxl;
    assign dcache_io_ptw_gstatus_sd_rv32 = _ptw_io_requestor_0_gstatus_sd_rv32;
    assign dcache_io_ptw_gstatus_zero1 = _ptw_io_requestor_0_gstatus_zero1;
    assign dcache_io_ptw_gstatus_tsr = _ptw_io_requestor_0_gstatus_tsr;
    assign dcache_io_ptw_gstatus_tw = _ptw_io_requestor_0_gstatus_tw;
    assign dcache_io_ptw_gstatus_tvm = _ptw_io_requestor_0_gstatus_tvm;
    assign dcache_io_ptw_gstatus_mxr = _ptw_io_requestor_0_gstatus_mxr;
    assign dcache_io_ptw_gstatus_sum = _ptw_io_requestor_0_gstatus_sum;
    assign dcache_io_ptw_gstatus_mprv = _ptw_io_requestor_0_gstatus_mprv;
    assign dcache_io_ptw_gstatus_xs = _ptw_io_requestor_0_gstatus_xs;
    assign dcache_io_ptw_gstatus_fs = _ptw_io_requestor_0_gstatus_fs;
    assign dcache_io_ptw_gstatus_mpp = _ptw_io_requestor_0_gstatus_mpp;
    assign dcache_io_ptw_gstatus_vs = _ptw_io_requestor_0_gstatus_vs;
    assign dcache_io_ptw_gstatus_spp = _ptw_io_requestor_0_gstatus_spp;
    assign dcache_io_ptw_gstatus_mpie = _ptw_io_requestor_0_gstatus_mpie;
    assign dcache_io_ptw_gstatus_ube = _ptw_io_requestor_0_gstatus_ube;
    assign dcache_io_ptw_gstatus_spie = _ptw_io_requestor_0_gstatus_spie;
    assign dcache_io_ptw_gstatus_upie = _ptw_io_requestor_0_gstatus_upie;
    assign dcache_io_ptw_gstatus_mie = _ptw_io_requestor_0_gstatus_mie;
    assign dcache_io_ptw_gstatus_hie = _ptw_io_requestor_0_gstatus_hie;
    assign dcache_io_ptw_gstatus_sie = _ptw_io_requestor_0_gstatus_sie;
    assign dcache_io_ptw_gstatus_uie = _ptw_io_requestor_0_gstatus_uie;
    assign dcache_io_ptw_pmp_0_cfg_l = _ptw_io_requestor_0_pmp_0_cfg_l;
    assign dcache_io_ptw_pmp_0_cfg_res = _ptw_io_requestor_0_pmp_0_cfg_res;
    assign dcache_io_ptw_pmp_0_cfg_a = _ptw_io_requestor_0_pmp_0_cfg_a;
    assign dcache_io_ptw_pmp_0_cfg_x = _ptw_io_requestor_0_pmp_0_cfg_x;
    assign dcache_io_ptw_pmp_0_cfg_w = _ptw_io_requestor_0_pmp_0_cfg_w;
    assign dcache_io_ptw_pmp_0_cfg_r = _ptw_io_requestor_0_pmp_0_cfg_r;
    assign dcache_io_ptw_pmp_0_addr = _ptw_io_requestor_0_pmp_0_addr;
    assign dcache_io_ptw_pmp_0_mask = _ptw_io_requestor_0_pmp_0_mask;
    assign dcache_io_ptw_pmp_1_cfg_l = _ptw_io_requestor_0_pmp_1_cfg_l;
    assign dcache_io_ptw_pmp_1_cfg_res = _ptw_io_requestor_0_pmp_1_cfg_res;
    assign dcache_io_ptw_pmp_1_cfg_a = _ptw_io_requestor_0_pmp_1_cfg_a;
    assign dcache_io_ptw_pmp_1_cfg_x = _ptw_io_requestor_0_pmp_1_cfg_x;
    assign dcache_io_ptw_pmp_1_cfg_w = _ptw_io_requestor_0_pmp_1_cfg_w;
    assign dcache_io_ptw_pmp_1_cfg_r = _ptw_io_requestor_0_pmp_1_cfg_r;
    assign dcache_io_ptw_pmp_1_addr = _ptw_io_requestor_0_pmp_1_addr;
    assign dcache_io_ptw_pmp_1_mask = _ptw_io_requestor_0_pmp_1_mask;
    assign dcache_io_ptw_pmp_2_cfg_l = _ptw_io_requestor_0_pmp_2_cfg_l;
    assign dcache_io_ptw_pmp_2_cfg_res = _ptw_io_requestor_0_pmp_2_cfg_res;
    assign dcache_io_ptw_pmp_2_cfg_a = _ptw_io_requestor_0_pmp_2_cfg_a;
    assign dcache_io_ptw_pmp_2_cfg_x = _ptw_io_requestor_0_pmp_2_cfg_x;
    assign dcache_io_ptw_pmp_2_cfg_w = _ptw_io_requestor_0_pmp_2_cfg_w;
    assign dcache_io_ptw_pmp_2_cfg_r = _ptw_io_requestor_0_pmp_2_cfg_r;
    assign dcache_io_ptw_pmp_2_addr = _ptw_io_requestor_0_pmp_2_addr;
    assign dcache_io_ptw_pmp_2_mask = _ptw_io_requestor_0_pmp_2_mask;
    assign dcache_io_ptw_pmp_3_cfg_l = _ptw_io_requestor_0_pmp_3_cfg_l;
    assign dcache_io_ptw_pmp_3_cfg_res = _ptw_io_requestor_0_pmp_3_cfg_res;
    assign dcache_io_ptw_pmp_3_cfg_a = _ptw_io_requestor_0_pmp_3_cfg_a;
    assign dcache_io_ptw_pmp_3_cfg_x = _ptw_io_requestor_0_pmp_3_cfg_x;
    assign dcache_io_ptw_pmp_3_cfg_w = _ptw_io_requestor_0_pmp_3_cfg_w;
    assign dcache_io_ptw_pmp_3_cfg_r = _ptw_io_requestor_0_pmp_3_cfg_r;
    assign dcache_io_ptw_pmp_3_addr = _ptw_io_requestor_0_pmp_3_addr;
    assign dcache_io_ptw_pmp_3_mask = _ptw_io_requestor_0_pmp_3_mask;
    assign dcache_io_ptw_pmp_4_cfg_l = _ptw_io_requestor_0_pmp_4_cfg_l;
    assign dcache_io_ptw_pmp_4_cfg_res = _ptw_io_requestor_0_pmp_4_cfg_res;
    assign dcache_io_ptw_pmp_4_cfg_a = _ptw_io_requestor_0_pmp_4_cfg_a;
    assign dcache_io_ptw_pmp_4_cfg_x = _ptw_io_requestor_0_pmp_4_cfg_x;
    assign dcache_io_ptw_pmp_4_cfg_w = _ptw_io_requestor_0_pmp_4_cfg_w;
    assign dcache_io_ptw_pmp_4_cfg_r = _ptw_io_requestor_0_pmp_4_cfg_r;
    assign dcache_io_ptw_pmp_4_addr = _ptw_io_requestor_0_pmp_4_addr;
    assign dcache_io_ptw_pmp_4_mask = _ptw_io_requestor_0_pmp_4_mask;
    assign dcache_io_ptw_pmp_5_cfg_l = _ptw_io_requestor_0_pmp_5_cfg_l;
    assign dcache_io_ptw_pmp_5_cfg_res = _ptw_io_requestor_0_pmp_5_cfg_res;
    assign dcache_io_ptw_pmp_5_cfg_a = _ptw_io_requestor_0_pmp_5_cfg_a;
    assign dcache_io_ptw_pmp_5_cfg_x = _ptw_io_requestor_0_pmp_5_cfg_x;
    assign dcache_io_ptw_pmp_5_cfg_w = _ptw_io_requestor_0_pmp_5_cfg_w;
    assign dcache_io_ptw_pmp_5_cfg_r = _ptw_io_requestor_0_pmp_5_cfg_r;
    assign dcache_io_ptw_pmp_5_addr = _ptw_io_requestor_0_pmp_5_addr;
    assign dcache_io_ptw_pmp_5_mask = _ptw_io_requestor_0_pmp_5_mask;
    assign dcache_io_ptw_pmp_6_cfg_l = _ptw_io_requestor_0_pmp_6_cfg_l;
    assign dcache_io_ptw_pmp_6_cfg_res = _ptw_io_requestor_0_pmp_6_cfg_res;
    assign dcache_io_ptw_pmp_6_cfg_a = _ptw_io_requestor_0_pmp_6_cfg_a;
    assign dcache_io_ptw_pmp_6_cfg_x = _ptw_io_requestor_0_pmp_6_cfg_x;
    assign dcache_io_ptw_pmp_6_cfg_w = _ptw_io_requestor_0_pmp_6_cfg_w;
    assign dcache_io_ptw_pmp_6_cfg_r = _ptw_io_requestor_0_pmp_6_cfg_r;
    assign dcache_io_ptw_pmp_6_addr = _ptw_io_requestor_0_pmp_6_addr;
    assign dcache_io_ptw_pmp_6_mask = _ptw_io_requestor_0_pmp_6_mask;
    assign dcache_io_ptw_pmp_7_cfg_l = _ptw_io_requestor_0_pmp_7_cfg_l;
    assign dcache_io_ptw_pmp_7_cfg_res = _ptw_io_requestor_0_pmp_7_cfg_res;
    assign dcache_io_ptw_pmp_7_cfg_a = _ptw_io_requestor_0_pmp_7_cfg_a;
    assign dcache_io_ptw_pmp_7_cfg_x = _ptw_io_requestor_0_pmp_7_cfg_x;
    assign dcache_io_ptw_pmp_7_cfg_w = _ptw_io_requestor_0_pmp_7_cfg_w;
    assign dcache_io_ptw_pmp_7_cfg_r = _ptw_io_requestor_0_pmp_7_cfg_r;
    assign dcache_io_ptw_pmp_7_addr = _ptw_io_requestor_0_pmp_7_addr;
    assign dcache_io_ptw_pmp_7_mask = _ptw_io_requestor_0_pmp_7_mask;
    assign dcache_io_ptw_customCSRs_csrs_0_ren = _ptw_io_requestor_0_customCSRs_csrs_0_ren;
    assign dcache_io_ptw_customCSRs_csrs_0_wen = _ptw_io_requestor_0_customCSRs_csrs_0_wen;
    assign dcache_io_ptw_customCSRs_csrs_0_wdata = _ptw_io_requestor_0_customCSRs_csrs_0_wdata;
    assign dcache_io_ptw_customCSRs_csrs_0_value = _ptw_io_requestor_0_customCSRs_csrs_0_value;
    assign _dcache_io_ptw_customCSRs_csrs_0_stall = dcache_io_ptw_customCSRs_csrs_0_stall;
    assign _dcache_io_ptw_customCSRs_csrs_0_set = dcache_io_ptw_customCSRs_csrs_0_set;
    assign _dcache_io_ptw_customCSRs_csrs_0_sdata = dcache_io_ptw_customCSRs_csrs_0_sdata;
    assign dcache_io_ptw_customCSRs_csrs_1_ren = _ptw_io_requestor_0_customCSRs_csrs_1_ren;
    assign dcache_io_ptw_customCSRs_csrs_1_wen = _ptw_io_requestor_0_customCSRs_csrs_1_wen;
    assign dcache_io_ptw_customCSRs_csrs_1_wdata = _ptw_io_requestor_0_customCSRs_csrs_1_wdata;
    assign dcache_io_ptw_customCSRs_csrs_1_value = _ptw_io_requestor_0_customCSRs_csrs_1_value;
    assign _dcache_io_ptw_customCSRs_csrs_1_stall = dcache_io_ptw_customCSRs_csrs_1_stall;
    assign _dcache_io_ptw_customCSRs_csrs_1_set = dcache_io_ptw_customCSRs_csrs_1_set;
    assign _dcache_io_ptw_customCSRs_csrs_1_sdata = dcache_io_ptw_customCSRs_csrs_1_sdata;
    assign dcache_io_ptw_customCSRs_csrs_2_ren = _ptw_io_requestor_0_customCSRs_csrs_2_ren;
    assign dcache_io_ptw_customCSRs_csrs_2_wen = _ptw_io_requestor_0_customCSRs_csrs_2_wen;
    assign dcache_io_ptw_customCSRs_csrs_2_wdata = _ptw_io_requestor_0_customCSRs_csrs_2_wdata;
    assign dcache_io_ptw_customCSRs_csrs_2_value = _ptw_io_requestor_0_customCSRs_csrs_2_value;
    assign _dcache_io_ptw_customCSRs_csrs_2_stall = dcache_io_ptw_customCSRs_csrs_2_stall;
    assign _dcache_io_ptw_customCSRs_csrs_2_set = dcache_io_ptw_customCSRs_csrs_2_set;
    assign _dcache_io_ptw_customCSRs_csrs_2_sdata = dcache_io_ptw_customCSRs_csrs_2_sdata;
    assign dcache_io_ptw_customCSRs_csrs_3_ren = _ptw_io_requestor_0_customCSRs_csrs_3_ren;
    assign dcache_io_ptw_customCSRs_csrs_3_wen = _ptw_io_requestor_0_customCSRs_csrs_3_wen;
    assign dcache_io_ptw_customCSRs_csrs_3_wdata = _ptw_io_requestor_0_customCSRs_csrs_3_wdata;
    assign dcache_io_ptw_customCSRs_csrs_3_value = _ptw_io_requestor_0_customCSRs_csrs_3_value;
    assign _dcache_io_ptw_customCSRs_csrs_3_stall = dcache_io_ptw_customCSRs_csrs_3_stall;
    assign _dcache_io_ptw_customCSRs_csrs_3_set = dcache_io_ptw_customCSRs_csrs_3_set;
    assign _dcache_io_ptw_customCSRs_csrs_3_sdata = dcache_io_ptw_customCSRs_csrs_3_sdata;
    assign dcache_tlb_port_req_valid = 1'h0;
    assign dcache_tlb_port_req_bits_vaddr = 34'h0;
    assign dcache_tlb_port_req_bits_passthrough = 1'h0;
    assign dcache_tlb_port_req_bits_size = 2'h0;
    assign dcache_tlb_port_req_bits_cmd = 5'h0;
    assign dcache_tlb_port_req_bits_prv = 2'h0;
    assign dcache_tlb_port_req_bits_v = 1'h0;
    assign dcache_tlb_port_s2_kill = 1'h0;
    
  wire        widget_1_auto_in_a_ready;
  wire        widget_1_auto_in_d_valid;
  wire [2:0]  widget_1_auto_in_d_bits_opcode;
  wire [1:0]  widget_1_auto_in_d_bits_param;
  wire [3:0]  widget_1_auto_in_d_bits_size;
  wire        widget_1_auto_in_d_bits_source;
  wire [1:0]  widget_1_auto_in_d_bits_sink;
  wire        widget_1_auto_in_d_bits_denied;
  wire [63:0] widget_1_auto_in_d_bits_data;
  wire        widget_1_auto_in_d_bits_corrupt;
  wire frontend_clock;
    wire frontend_reset;
    wire frontend_auto_icache_master_out_a_ready;
    wire frontend_auto_icache_master_out_a_valid;
    wire[2:0] frontend_auto_icache_master_out_a_bits_opcode;
    wire[2:0] frontend_auto_icache_master_out_a_bits_param;
    wire[3:0] frontend_auto_icache_master_out_a_bits_size;
    wire frontend_auto_icache_master_out_a_bits_source;
    wire[31:0] frontend_auto_icache_master_out_a_bits_address;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_bufferable;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_modifiable;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_privileged;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_secure;
    wire frontend_auto_icache_master_out_a_bits_user_amba_prot_fetch;
    wire[7:0] frontend_auto_icache_master_out_a_bits_mask;
    wire[63:0] frontend_auto_icache_master_out_a_bits_data;
    wire frontend_auto_icache_master_out_a_bits_corrupt;
    wire frontend_auto_icache_master_out_d_ready;
    wire frontend_auto_icache_master_out_d_valid;
    wire[2:0] frontend_auto_icache_master_out_d_bits_opcode;
    wire[1:0] frontend_auto_icache_master_out_d_bits_param;
    wire[3:0] frontend_auto_icache_master_out_d_bits_size;
    wire frontend_auto_icache_master_out_d_bits_source;
    wire[1:0] frontend_auto_icache_master_out_d_bits_sink;
    wire frontend_auto_icache_master_out_d_bits_denied;
    wire[63:0] frontend_auto_icache_master_out_d_bits_data;
    wire frontend_auto_icache_master_out_d_bits_corrupt;
    wire[31:0] frontend_auto_reset_vector_sink_in;
    wire frontend_io_cpu_might_request;
    wire frontend_io_cpu_clock_enabled;
    wire frontend_io_cpu_req_valid;
    wire[33:0] frontend_io_cpu_req_bits_pc;
    wire frontend_io_cpu_req_bits_speculative;
    wire frontend_io_cpu_sfence_valid;
    wire frontend_io_cpu_sfence_bits_rs1;
    wire frontend_io_cpu_sfence_bits_rs2;
    wire[32:0] frontend_io_cpu_sfence_bits_addr;
    wire frontend_io_cpu_sfence_bits_asid;
    wire frontend_io_cpu_sfence_bits_hv;
    wire frontend_io_cpu_sfence_bits_hg;
    wire frontend_io_cpu_resp_ready;
    wire frontend_io_cpu_resp_valid;
    wire[1:0] frontend_io_cpu_resp_bits_btb_cfiType;
    wire frontend_io_cpu_resp_bits_btb_taken;
    wire[1:0] frontend_io_cpu_resp_bits_btb_mask;
    wire frontend_io_cpu_resp_bits_btb_bridx;
    wire[32:0] frontend_io_cpu_resp_bits_btb_target;
    wire frontend_io_cpu_resp_bits_btb_entry;
    wire[7:0] frontend_io_cpu_resp_bits_btb_bht_history;
    wire frontend_io_cpu_resp_bits_btb_bht_value;
    wire[33:0] frontend_io_cpu_resp_bits_pc;
    wire[31:0] frontend_io_cpu_resp_bits_data;
    wire[1:0] frontend_io_cpu_resp_bits_mask;
    wire frontend_io_cpu_resp_bits_xcpt_pf_inst;
    wire frontend_io_cpu_resp_bits_xcpt_gf_inst;
    wire frontend_io_cpu_resp_bits_xcpt_ae_inst;
    wire frontend_io_cpu_resp_bits_replay;
    wire frontend_io_cpu_gpa_valid;
    wire[33:0] frontend_io_cpu_gpa_bits;
    wire frontend_io_cpu_btb_update_valid;
    wire[1:0] frontend_io_cpu_btb_update_bits_prediction_cfiType;
    wire frontend_io_cpu_btb_update_bits_prediction_taken;
    wire[1:0] frontend_io_cpu_btb_update_bits_prediction_mask;
    wire frontend_io_cpu_btb_update_bits_prediction_bridx;
    wire[32:0] frontend_io_cpu_btb_update_bits_prediction_target;
    wire frontend_io_cpu_btb_update_bits_prediction_entry;
    wire[7:0] frontend_io_cpu_btb_update_bits_prediction_bht_history;
    wire frontend_io_cpu_btb_update_bits_prediction_bht_value;
    wire[32:0] frontend_io_cpu_btb_update_bits_pc;
    wire[32:0] frontend_io_cpu_btb_update_bits_target;
    wire frontend_io_cpu_btb_update_bits_taken;
    wire frontend_io_cpu_btb_update_bits_isValid;
    wire[32:0] frontend_io_cpu_btb_update_bits_br_pc;
    wire[1:0] frontend_io_cpu_btb_update_bits_cfiType;
    wire frontend_io_cpu_bht_update_valid;
    wire[7:0] frontend_io_cpu_bht_update_bits_prediction_history;
    wire frontend_io_cpu_bht_update_bits_prediction_value;
    wire[32:0] frontend_io_cpu_bht_update_bits_pc;
    wire frontend_io_cpu_bht_update_bits_branch;
    wire frontend_io_cpu_bht_update_bits_taken;
    wire frontend_io_cpu_bht_update_bits_mispredict;
    wire frontend_io_cpu_ras_update_valid;
    wire[1:0] frontend_io_cpu_ras_update_bits_cfiType;
    wire[32:0] frontend_io_cpu_ras_update_bits_returnAddr;
    wire frontend_io_cpu_flush_icache;
    wire[33:0] frontend_io_cpu_npc;
    wire frontend_io_cpu_perf_acquire;
    wire frontend_io_cpu_perf_tlbMiss;
    wire frontend_io_cpu_progress;
    wire frontend_io_ptw_req_ready;
    wire frontend_io_ptw_req_valid;
    wire frontend_io_ptw_req_bits_valid;
    wire[20:0] frontend_io_ptw_req_bits_bits_addr;
    wire frontend_io_ptw_req_bits_bits_need_gpa;
    wire frontend_io_ptw_req_bits_bits_vstage1;
    wire frontend_io_ptw_req_bits_bits_stage2;
    wire frontend_io_ptw_resp_valid;
    wire frontend_io_ptw_resp_bits_ae_ptw;
    wire frontend_io_ptw_resp_bits_ae_final;
    wire frontend_io_ptw_resp_bits_pf;
    wire frontend_io_ptw_resp_bits_gf;
    wire frontend_io_ptw_resp_bits_hr;
    wire frontend_io_ptw_resp_bits_hw;
    wire frontend_io_ptw_resp_bits_hx;
    wire[9:0] frontend_io_ptw_resp_bits_pte_reserved_for_future;
    wire[43:0] frontend_io_ptw_resp_bits_pte_ppn;
    wire[1:0] frontend_io_ptw_resp_bits_pte_reserved_for_software;
    wire frontend_io_ptw_resp_bits_pte_d;
    wire frontend_io_ptw_resp_bits_pte_a;
    wire frontend_io_ptw_resp_bits_pte_g;
    wire frontend_io_ptw_resp_bits_pte_u;
    wire frontend_io_ptw_resp_bits_pte_x;
    wire frontend_io_ptw_resp_bits_pte_w;
    wire frontend_io_ptw_resp_bits_pte_r;
    wire frontend_io_ptw_resp_bits_pte_v;
    wire[1:0] frontend_io_ptw_resp_bits_level;
    wire frontend_io_ptw_resp_bits_fragmented_superpage;
    wire frontend_io_ptw_resp_bits_homogeneous;
    wire frontend_io_ptw_resp_bits_gpa_valid;
    wire[32:0] frontend_io_ptw_resp_bits_gpa_bits;
    wire frontend_io_ptw_resp_bits_gpa_is_pte;
    wire[3:0] frontend_io_ptw_ptbr_mode;
    wire[15:0] frontend_io_ptw_ptbr_asid;
    wire[43:0] frontend_io_ptw_ptbr_ppn;
    wire[3:0] frontend_io_ptw_hgatp_mode;
    wire[15:0] frontend_io_ptw_hgatp_asid;
    wire[43:0] frontend_io_ptw_hgatp_ppn;
    wire[3:0] frontend_io_ptw_vsatp_mode;
    wire[15:0] frontend_io_ptw_vsatp_asid;
    wire[43:0] frontend_io_ptw_vsatp_ppn;
    wire frontend_io_ptw_status_debug;
    wire frontend_io_ptw_status_cease;
    wire frontend_io_ptw_status_wfi;
    wire[31:0] frontend_io_ptw_status_isa;
    wire[1:0] frontend_io_ptw_status_dprv;
    wire frontend_io_ptw_status_dv;
    wire[1:0] frontend_io_ptw_status_prv;
    wire frontend_io_ptw_status_v;
    wire frontend_io_ptw_status_sd;
    wire[22:0] frontend_io_ptw_status_zero2;
    wire frontend_io_ptw_status_mpv;
    wire frontend_io_ptw_status_gva;
    wire frontend_io_ptw_status_mbe;
    wire frontend_io_ptw_status_sbe;
    wire[1:0] frontend_io_ptw_status_sxl;
    wire[1:0] frontend_io_ptw_status_uxl;
    wire frontend_io_ptw_status_sd_rv32;
    wire[7:0] frontend_io_ptw_status_zero1;
    wire frontend_io_ptw_status_tsr;
    wire frontend_io_ptw_status_tw;
    wire frontend_io_ptw_status_tvm;
    wire frontend_io_ptw_status_mxr;
    wire frontend_io_ptw_status_sum;
    wire frontend_io_ptw_status_mprv;
    wire[1:0] frontend_io_ptw_status_xs;
    wire[1:0] frontend_io_ptw_status_fs;
    wire[1:0] frontend_io_ptw_status_mpp;
    wire[1:0] frontend_io_ptw_status_vs;
    wire frontend_io_ptw_status_spp;
    wire frontend_io_ptw_status_mpie;
    wire frontend_io_ptw_status_ube;
    wire frontend_io_ptw_status_spie;
    wire frontend_io_ptw_status_upie;
    wire frontend_io_ptw_status_mie;
    wire frontend_io_ptw_status_hie;
    wire frontend_io_ptw_status_sie;
    wire frontend_io_ptw_status_uie;
    wire[29:0] frontend_io_ptw_hstatus_zero6;
    wire[1:0] frontend_io_ptw_hstatus_vsxl;
    wire[8:0] frontend_io_ptw_hstatus_zero5;
    wire frontend_io_ptw_hstatus_vtsr;
    wire frontend_io_ptw_hstatus_vtw;
    wire frontend_io_ptw_hstatus_vtvm;
    wire[1:0] frontend_io_ptw_hstatus_zero3;
    wire[5:0] frontend_io_ptw_hstatus_vgein;
    wire[1:0] frontend_io_ptw_hstatus_zero2;
    wire frontend_io_ptw_hstatus_hu;
    wire frontend_io_ptw_hstatus_spvp;
    wire frontend_io_ptw_hstatus_spv;
    wire frontend_io_ptw_hstatus_gva;
    wire frontend_io_ptw_hstatus_vsbe;
    wire[4:0] frontend_io_ptw_hstatus_zero1;
    wire frontend_io_ptw_gstatus_debug;
    wire frontend_io_ptw_gstatus_cease;
    wire frontend_io_ptw_gstatus_wfi;
    wire[31:0] frontend_io_ptw_gstatus_isa;
    wire[1:0] frontend_io_ptw_gstatus_dprv;
    wire frontend_io_ptw_gstatus_dv;
    wire[1:0] frontend_io_ptw_gstatus_prv;
    wire frontend_io_ptw_gstatus_v;
    wire frontend_io_ptw_gstatus_sd;
    wire[22:0] frontend_io_ptw_gstatus_zero2;
    wire frontend_io_ptw_gstatus_mpv;
    wire frontend_io_ptw_gstatus_gva;
    wire frontend_io_ptw_gstatus_mbe;
    wire frontend_io_ptw_gstatus_sbe;
    wire[1:0] frontend_io_ptw_gstatus_sxl;
    wire[1:0] frontend_io_ptw_gstatus_uxl;
    wire frontend_io_ptw_gstatus_sd_rv32;
    wire[7:0] frontend_io_ptw_gstatus_zero1;
    wire frontend_io_ptw_gstatus_tsr;
    wire frontend_io_ptw_gstatus_tw;
    wire frontend_io_ptw_gstatus_tvm;
    wire frontend_io_ptw_gstatus_mxr;
    wire frontend_io_ptw_gstatus_sum;
    wire frontend_io_ptw_gstatus_mprv;
    wire[1:0] frontend_io_ptw_gstatus_xs;
    wire[1:0] frontend_io_ptw_gstatus_fs;
    wire[1:0] frontend_io_ptw_gstatus_mpp;
    wire[1:0] frontend_io_ptw_gstatus_vs;
    wire frontend_io_ptw_gstatus_spp;
    wire frontend_io_ptw_gstatus_mpie;
    wire frontend_io_ptw_gstatus_ube;
    wire frontend_io_ptw_gstatus_spie;
    wire frontend_io_ptw_gstatus_upie;
    wire frontend_io_ptw_gstatus_mie;
    wire frontend_io_ptw_gstatus_hie;
    wire frontend_io_ptw_gstatus_sie;
    wire frontend_io_ptw_gstatus_uie;
    wire frontend_io_ptw_pmp_0_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_0_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_0_cfg_a;
    wire frontend_io_ptw_pmp_0_cfg_x;
    wire frontend_io_ptw_pmp_0_cfg_w;
    wire frontend_io_ptw_pmp_0_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_0_addr;
    wire[31:0] frontend_io_ptw_pmp_0_mask;
    wire frontend_io_ptw_pmp_1_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_1_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_1_cfg_a;
    wire frontend_io_ptw_pmp_1_cfg_x;
    wire frontend_io_ptw_pmp_1_cfg_w;
    wire frontend_io_ptw_pmp_1_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_1_addr;
    wire[31:0] frontend_io_ptw_pmp_1_mask;
    wire frontend_io_ptw_pmp_2_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_2_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_2_cfg_a;
    wire frontend_io_ptw_pmp_2_cfg_x;
    wire frontend_io_ptw_pmp_2_cfg_w;
    wire frontend_io_ptw_pmp_2_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_2_addr;
    wire[31:0] frontend_io_ptw_pmp_2_mask;
    wire frontend_io_ptw_pmp_3_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_3_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_3_cfg_a;
    wire frontend_io_ptw_pmp_3_cfg_x;
    wire frontend_io_ptw_pmp_3_cfg_w;
    wire frontend_io_ptw_pmp_3_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_3_addr;
    wire[31:0] frontend_io_ptw_pmp_3_mask;
    wire frontend_io_ptw_pmp_4_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_4_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_4_cfg_a;
    wire frontend_io_ptw_pmp_4_cfg_x;
    wire frontend_io_ptw_pmp_4_cfg_w;
    wire frontend_io_ptw_pmp_4_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_4_addr;
    wire[31:0] frontend_io_ptw_pmp_4_mask;
    wire frontend_io_ptw_pmp_5_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_5_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_5_cfg_a;
    wire frontend_io_ptw_pmp_5_cfg_x;
    wire frontend_io_ptw_pmp_5_cfg_w;
    wire frontend_io_ptw_pmp_5_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_5_addr;
    wire[31:0] frontend_io_ptw_pmp_5_mask;
    wire frontend_io_ptw_pmp_6_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_6_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_6_cfg_a;
    wire frontend_io_ptw_pmp_6_cfg_x;
    wire frontend_io_ptw_pmp_6_cfg_w;
    wire frontend_io_ptw_pmp_6_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_6_addr;
    wire[31:0] frontend_io_ptw_pmp_6_mask;
    wire frontend_io_ptw_pmp_7_cfg_l;
    wire[1:0] frontend_io_ptw_pmp_7_cfg_res;
    wire[1:0] frontend_io_ptw_pmp_7_cfg_a;
    wire frontend_io_ptw_pmp_7_cfg_x;
    wire frontend_io_ptw_pmp_7_cfg_w;
    wire frontend_io_ptw_pmp_7_cfg_r;
    wire[29:0] frontend_io_ptw_pmp_7_addr;
    wire[31:0] frontend_io_ptw_pmp_7_mask;
    wire frontend_io_ptw_customCSRs_csrs_0_ren;
    wire frontend_io_ptw_customCSRs_csrs_0_wen;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_0_wdata;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_0_value;
    wire frontend_io_ptw_customCSRs_csrs_0_stall;
    wire frontend_io_ptw_customCSRs_csrs_0_set;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_0_sdata;
    wire frontend_io_ptw_customCSRs_csrs_1_ren;
    wire frontend_io_ptw_customCSRs_csrs_1_wen;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_1_wdata;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_1_value;
    wire frontend_io_ptw_customCSRs_csrs_1_stall;
    wire frontend_io_ptw_customCSRs_csrs_1_set;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_1_sdata;
    wire frontend_io_ptw_customCSRs_csrs_2_ren;
    wire frontend_io_ptw_customCSRs_csrs_2_wen;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_2_wdata;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_2_value;
    wire frontend_io_ptw_customCSRs_csrs_2_stall;
    wire frontend_io_ptw_customCSRs_csrs_2_set;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_2_sdata;
    wire frontend_io_ptw_customCSRs_csrs_3_ren;
    wire frontend_io_ptw_customCSRs_csrs_3_wen;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_3_wdata;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_3_value;
    wire frontend_io_ptw_customCSRs_csrs_3_stall;
    wire frontend_io_ptw_customCSRs_csrs_3_set;
    wire[63:0] frontend_io_ptw_customCSRs_csrs_3_sdata;
    wire frontend_io_errors_bus_valid;
    wire[31:0] frontend_io_errors_bus_bits;

    wire frontend__GEN ; 
    wire frontend__GEN_0 ; 
    wire[1:0] frontend__GEN_1 ; 
    wire frontend__GEN_2 ; 
    wire frontend__GEN_3 ; 
    wire frontend__GEN_4 ; 
    wire frontend__GEN_5 ; 
    wire[32:0] frontend__s2_pc_32to0 ; 
    wire[32:0] frontend___io_cpu_npc_output_32to0 ; 
    wire frontend__GEN_6 ; 
    wire frontend__GEN_7 ; 
    reg frontend_s2_tlb_resp_cacheable ; 
    reg frontend_s2_tlb_resp_gf_inst ; 
    reg frontend_s2_tlb_resp_pf_inst ; 
    reg frontend_s2_btb_resp_bits_bht_value ; reg[7:0] frontend_s2_btb_resp_bits_bht_history ; 
    reg frontend_s2_btb_resp_bits_entry ; reg[32:0] frontend_s2_btb_resp_bits_target ; 
    reg frontend_s2_btb_resp_bits_bridx ; reg[1:0] frontend_s2_btb_resp_bits_mask ; reg[1:0] frontend_s2_btb_resp_bits_cfiType ; reg[33:0] frontend_s2_pc ; reg[33:0] frontend_s1_pc ; 
    wire frontend__io_ptw_req_valid_output ; 
    wire frontend__tlb_io_req_ready ; 
    wire frontend__tlb_io_resp_miss ; 
    wire[31:0] frontend__tlb_io_resp_paddr ; 
    wire[33:0] frontend__tlb_io_resp_gpa ; 
    wire frontend__tlb_io_resp_gpa_is_pte ; 
    wire frontend__tlb_io_resp_pf_ld ; 
    wire frontend__tlb_io_resp_pf_st ; 
    wire frontend__tlb_io_resp_pf_inst ; 
    wire frontend__tlb_io_resp_gf_ld ; 
    wire frontend__tlb_io_resp_gf_st ; 
    wire frontend__tlb_io_resp_gf_inst ; 
    wire frontend__tlb_io_resp_ae_ld ; 
    wire frontend__tlb_io_resp_ae_st ; 
    wire frontend__tlb_io_resp_ae_inst ; 
    wire frontend__tlb_io_resp_ma_ld ; 
    wire frontend__tlb_io_resp_ma_st ; 
    wire frontend__tlb_io_resp_ma_inst ; 
    wire frontend__tlb_io_resp_cacheable ; 
    wire frontend__tlb_io_resp_must_alloc ; 
    wire frontend__tlb_io_resp_prefetchable ; 
    wire frontend__fq_io_enq_ready ; 
    wire[4:0] frontend__fq_io_mask ; 
    wire frontend__icache_io_resp_valid ; 
    wire[31:0] frontend__icache_io_resp_bits_data ; 
    wire frontend__icache_io_resp_bits_replay ; 
    wire frontend__icache_io_resp_bits_ae ; 
    wire[31:0] frontend_resetVectorSinkNodeIn = frontend_auto_reset_vector_sink_in ; 
    wire frontend_s2_redirect = frontend_io_cpu_req_valid ; 
    wire frontend_s2_btb_taken =1'h0; 
    wire frontend_predicted_taken =1'h0; 
    wire frontend_clock_en ; 
    wire frontend_s0_valid ;  
    wire frontend_icache_clock;
    wire frontend_icache_reset;
    wire frontend_icache_auto_master_out_a_ready;
    wire frontend_icache_auto_master_out_a_valid;
    wire[2:0] frontend_icache_auto_master_out_a_bits_opcode;
    wire[2:0] frontend_icache_auto_master_out_a_bits_param;
    wire[3:0] frontend_icache_auto_master_out_a_bits_size;
    wire frontend_icache_auto_master_out_a_bits_source;
    wire[31:0] frontend_icache_auto_master_out_a_bits_address;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_bufferable;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_modifiable;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_privileged;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_secure;
    wire frontend_icache_auto_master_out_a_bits_user_amba_prot_fetch;
    wire[7:0] frontend_icache_auto_master_out_a_bits_mask;
    wire[63:0] frontend_icache_auto_master_out_a_bits_data;
    wire frontend_icache_auto_master_out_a_bits_corrupt;
    wire frontend_icache_auto_master_out_d_ready;
    wire frontend_icache_auto_master_out_d_valid;
    wire[2:0] frontend_icache_auto_master_out_d_bits_opcode;
    wire[1:0] frontend_icache_auto_master_out_d_bits_param;
    wire[3:0] frontend_icache_auto_master_out_d_bits_size;
    wire frontend_icache_auto_master_out_d_bits_source;
    wire[1:0] frontend_icache_auto_master_out_d_bits_sink;
    wire frontend_icache_auto_master_out_d_bits_denied;
    wire[63:0] frontend_icache_auto_master_out_d_bits_data;
    wire frontend_icache_auto_master_out_d_bits_corrupt;
    wire frontend_icache_io_req_ready;
    wire frontend_icache_io_req_valid;
    wire[32:0] frontend_icache_io_req_bits_addr;
    wire[31:0] frontend_icache_io_s1_paddr;
    wire[32:0] frontend_icache_io_s2_vaddr;
    wire frontend_icache_io_s1_kill;
    wire frontend_icache_io_s2_kill;
    wire frontend_icache_io_s2_cacheable;
    wire frontend_icache_io_s2_prefetch;
    wire frontend_icache_io_resp_valid;
    wire[31:0] frontend_icache_io_resp_bits_data;
    wire frontend_icache_io_resp_bits_replay;
    wire frontend_icache_io_resp_bits_ae;
    wire frontend_icache_io_invalidate;
    wire frontend_icache_io_errors_bus_valid;
    wire[31:0] frontend_icache_io_errors_bus_bits;
    wire frontend_icache_io_perf_acquire;
    wire frontend_icache_io_clock_enabled;
    wire frontend_icache_io_keep_clock_enabled;

    wire frontend_icache__GEN ; 
    wire[31:0] frontend_icache_data_arrays_1_dout_1_data_0 ; 
    wire frontend_icache__GEN_0 ; 
    wire[31:0] frontend_icache_data_arrays_0_dout_data_0 ; 
    wire frontend_icache__GEN_1 ; 
    wire[20:0] frontend_icache_tag_array_tag_rdata_data_0 ; 
    wire frontend_icache_masterNodeOut_a_ready = frontend_icache_auto_master_out_a_ready ; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_readalloc = frontend_icache_io_s2_cacheable ; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_writealloc = frontend_icache_io_s2_cacheable ; 
    wire frontend_icache_masterNodeOut_d_valid = frontend_icache_auto_master_out_d_valid ; 
    wire[2:0] frontend_icache_masterNodeOut_d_bits_opcode = frontend_icache_auto_master_out_d_bits_opcode ; 
    wire[1:0] frontend_icache_masterNodeOut_d_bits_param = frontend_icache_auto_master_out_d_bits_param ; 
    wire[3:0] frontend_icache_masterNodeOut_d_bits_size = frontend_icache_auto_master_out_d_bits_size ; 
    wire frontend_icache_masterNodeOut_d_bits_source = frontend_icache_auto_master_out_d_bits_source ; 
    wire[1:0] frontend_icache_masterNodeOut_d_bits_sink = frontend_icache_auto_master_out_d_bits_sink ; 
    wire frontend_icache_masterNodeOut_d_bits_denied = frontend_icache_auto_master_out_d_bits_denied ; 
    wire[63:0] frontend_icache_masterNodeOut_d_bits_data = frontend_icache_auto_master_out_d_bits_data ; 
    wire frontend_icache_masterNodeOut_d_bits_corrupt = frontend_icache_auto_master_out_d_bits_corrupt ; 
    wire frontend_icache_tag_array_MPORT_clk = frontend_icache_clock ; 
    wire frontend_icache_tag_array_tag_rdata_clk = frontend_icache_clock ; 
    wire frontend_icache_data_arrays_0_MPORT_1_clk = frontend_icache_clock ; 
    wire frontend_icache_data_arrays_0_dout_clk = frontend_icache_clock ; 
    wire frontend_icache_data_arrays_1_MPORT_2_clk = frontend_icache_clock ; 
    wire frontend_icache_data_arrays_1_dout_1_clk = frontend_icache_clock ; 
    wire[31:0] frontend_icache__GEN_2 =32'h0; 
    wire[31:0] frontend_icache__GEN_3 =32'h0; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH_shiftAmount =2'h2; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_a_opcode =3'h4; 
    wire[3:0] frontend_icache__GEN_4 =4'h0; 
    wire[3:0] frontend_icache__GEN_5 =4'h0; 
    wire[1:0] frontend_icache__GEN_6 =2'h0; 
    wire[1:0] frontend_icache__GEN_7 =2'h0; 
    wire[2:0] frontend_icache__GEN_8 =3'h0; 
    wire[2:0] frontend_icache__GEN_9 =3'h0; 
    wire[2:0] frontend_icache__GEN_10 =3'h0; 
    wire[63:0] frontend_icache__GEN_11 =64'h0; 
    wire[63:0] frontend_icache__GEN_12 =64'h0; 
    wire[7:0] frontend_icache__GEN_13 =8'h0; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_bufferable =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_modifiable =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_privileged =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_secure =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_user_amba_prot_fetch =1'h1; 
    wire frontend_icache_tag_array_MPORT_mask_0 =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc =1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_1 =1'h1; 
    wire frontend_icache__GEN_14 =1'h1; 
    wire frontend_icache_s1_tag_disparity_0 =1'h0; 
    wire frontend_icache_scratchpadHit =1'h0; 
    wire frontend_icache_way =1'h0; 
    wire frontend_icache_way_1 =1'h0; 
    wire frontend_icache_s1s2_full_word_write =1'h0; 
    wire frontend_icache__s2_tag_hit_WIRE_0 =1'h0; 
    wire frontend_icache_s1_scratchpad_hit =1'h0; 
    wire frontend_icache_s2_report_uncorrectable_error =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_source =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_bufferable =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_modifiable =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_readalloc =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_writealloc =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_privileged =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_secure =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_user_amba_prot_fetch =1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_corrupt =1'h0; 
    wire frontend_icache__GEN_15 =1'h0; 
    wire frontend_icache__GEN_16 =1'h0; 
    wire frontend_icache__GEN_17 =1'h0; 
    wire frontend_icache__GEN_18 =1'h0; 
    wire frontend_icache__GEN_19 =1'h0; 
    wire frontend_icache__GEN_20 =1'h0; 
    wire frontend_icache__GEN_21 =1'h0; 
    wire frontend_icache__GEN_22 =1'h0; 
    wire frontend_icache__GEN_23 =1'h0; 
    wire frontend_icache__GEN_24 =1'h0; 
    wire frontend_icache__GEN_25 =1'h0; 
    wire frontend_icache__GEN_26 =1'h0; 
    wire frontend_icache__GEN_27 =1'h0; 
    wire frontend_icache__GEN_28 =1'h0; 
    wire frontend_icache__GEN_29 =1'h0; 
    wire frontend_icache__GEN_30 =1'h0; 
    wire frontend_icache__GEN_31 =1'h0; 
    wire frontend_icache__GEN_32 =1'h0; 
    wire frontend_icache__GEN_33 =1'h0; 
    wire frontend_icache_s2_request_refill ; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_a_param =3'h0; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_a_size =4'h6; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_a_address ; 
    wire[7:0] frontend_icache_masterNodeOut_a_bits_a_mask ; 
    wire[63:0] frontend_icache_masterNodeOut_a_bits_a_data =64'h0; 
    reg frontend_icache_scratchpadOn ; 
    reg frontend_icache_s1_slaveValid ; 
    reg frontend_icache_s2_slaveValid ; 
    reg frontend_icache_s3_slaveValid ; 
    wire frontend_icache__io_req_ready_output ; 
    wire frontend_icache_s0_valid = frontend_icache__io_req_ready_output & frontend_icache_io_req_valid ; 
    reg frontend_icache_s1_valid ; reg[32:0] frontend_icache_s1_vaddr ; 
    wire frontend_icache_s1_tag_hit_0 ; 
    wire frontend_icache_s1_hit = frontend_icache_s1_tag_hit_0 | frontend_icache_s1_slaveValid ; 
    reg frontend_icache_s2_valid ; 
    reg frontend_icache_s2_hit ; 
    reg frontend_icache_invalidated ; 
    reg frontend_icache_refill_valid ; 
    reg frontend_icache_send_hint ; 
    wire frontend_icache_masterNodeOut_a_valid ; 
    wire frontend_icache_refill_fire = frontend_icache_masterNodeOut_a_ready & frontend_icache_masterNodeOut_a_valid & frontend_icache_send_hint ==1'h0; 
    reg frontend_icache_hint_outstanding ; 
    wire frontend_icache_s2_miss = frontend_icache_s2_valid & frontend_icache_s2_hit ==1'h0& frontend_icache_io_s2_kill ==1'h0; 
    wire frontend_icache_s1_can_request_refill =( frontend_icache_s2_miss | frontend_icache_refill_valid )==1'h0; 
    reg frontend_icache_s2_request_refill_REG ; 
  assign  frontend_icache_s2_request_refill = frontend_icache_s2_miss & frontend_icache_s2_request_refill_REG ; 
  assign  frontend_icache_masterNodeOut_a_valid = frontend_icache_s2_request_refill ; 
    wire frontend_icache__GEN_34 = frontend_icache_s1_valid & frontend_icache_s1_can_request_refill ; reg[31:0] frontend_icache_refill_paddr ; 
    wire frontend_icache__GEN_35 = frontend_icache_s1_valid & frontend_icache_s1_can_request_refill ; reg[32:0] frontend_icache_refill_vaddr ; 
    wire[19:0] frontend_icache_refill_tag = frontend_icache_refill_paddr [31:12]; 
    wire[5:0] frontend_icache_refill_idx = frontend_icache_refill_paddr [11:6]; 
    wire frontend_icache_masterNodeOut_d_ready ; 
    wire[5:0] frontend_icache_tag_array_MPORT_addr = frontend_icache_refill_idx ; 
    wire frontend_icache_refill_one_beat_opdata = frontend_icache_masterNodeOut_d_bits_opcode [0]; 
    wire frontend_icache_refill_one_beat = frontend_icache_masterNodeOut_d_ready & frontend_icache_masterNodeOut_d_valid & frontend_icache_refill_one_beat_opdata ; 
  assign  frontend_icache__io_req_ready_output =( frontend_icache_refill_one_beat | frontend_icache_s3_slaveValid )==1'h0; 
    wire frontend_icache__GEN_36 = frontend_icache_masterNodeOut_d_ready & frontend_icache_masterNodeOut_d_valid ; 
    wire[26:0] frontend_icache__GEN_37 =27'hFFF<< frontend_icache_masterNodeOut_d_bits_size ; 
    wire[11:0] frontend_icache__GEN_38 =~( frontend_icache__GEN_37 [11:0]); 
    wire[8:0] frontend_icache_beats1_decode = frontend_icache__GEN_38 [11:3]; 
    wire frontend_icache_beats1_opdata = frontend_icache_masterNodeOut_d_bits_opcode [0]; 
    wire[8:0] frontend_icache_beats1 = frontend_icache_beats1_opdata  ?  frontend_icache_beats1_decode :9'h0; reg[8:0] frontend_icache_counter ; 
    wire[9:0] frontend_icache__GEN_39 ={1'h0, frontend_icache_counter }-10'h1; 
    wire[8:0] frontend_icache_counter1 = frontend_icache__GEN_39 [8:0]; 
    wire frontend_icache_first = frontend_icache_counter ==9'h0; 
    wire frontend_icache_last = frontend_icache_counter ==9'h1| frontend_icache_beats1 ==9'h0; 
    wire frontend_icache_d_done = frontend_icache_last & frontend_icache__GEN_36 ; 
    wire[8:0] frontend_icache_refill_cnt = frontend_icache_beats1 &~ frontend_icache_counter1 ; 
    wire frontend_icache_refill_done = frontend_icache_refill_one_beat & frontend_icache_d_done ; 
    wire frontend_icache_tag_array_MPORT_en = frontend_icache_refill_done ; 
  assign  frontend_icache_masterNodeOut_d_ready = frontend_icache_s3_slaveValid ==1'h0; 
    wire[20:0] frontend_icache__GEN_40 ; 
    wire[5:0] frontend_icache__tag_rdata_WIRE ; 
    wire[20:0] frontend_icache_tag_array_MPORT_data_0 ; 
    wire[5:0] frontend_icache_tag_array_tag_rdata_addr ; 
    wire frontend_icache_tag_array_tag_rdata_en ;  
    wire[5:0] frontend_icache_tag_array_0_ext_R0_addr;
    wire frontend_icache_tag_array_0_ext_R0_en;
    wire frontend_icache_tag_array_0_ext_R0_clk;
    wire[20:0] frontend_icache_tag_array_0_ext_R0_data;
    wire[5:0] frontend_icache_tag_array_0_ext_W0_addr;
    wire frontend_icache_tag_array_0_ext_W0_en;
    wire frontend_icache_tag_array_0_ext_W0_clk;
    wire[20:0] frontend_icache_tag_array_0_ext_W0_data;

    reg[20:0] frontend_icache_tag_array_0_ext_Memory [0:63]; 
    reg frontend_icache_tag_array_0_ext__R0_en_d0 ; reg[5:0] frontend_icache_tag_array_0_ext__R0_addr_d0 ; 
  always @( posedge  frontend_icache_tag_array_0_ext_R0_clk )
         begin  
             frontend_icache_tag_array_0_ext__R0_en_d0  <= frontend_icache_tag_array_0_ext_R0_en ; 
             frontend_icache_tag_array_0_ext__R0_addr_d0  <= frontend_icache_tag_array_0_ext_R0_addr ;
         end
  always @( posedge  frontend_icache_tag_array_0_ext_W0_clk )
         begin 
             if ( frontend_icache_tag_array_0_ext_W0_en &1'h1) 
                 frontend_icache_tag_array_0_ext_Memory  [ frontend_icache_tag_array_0_ext_W0_addr ]<= frontend_icache_tag_array_0_ext_W0_data ;
         end
  assign  frontend_icache_tag_array_0_ext_R0_data = frontend_icache_tag_array_0_ext__R0_en_d0  ?  frontend_icache_tag_array_0_ext_Memory [ frontend_icache_tag_array_0_ext__R0_addr_d0 ]:21'bx;
    assign frontend_icache_tag_array_0_ext_R0_addr = frontend_icache_tag_array_tag_rdata_addr;
    assign frontend_icache_tag_array_0_ext_R0_en = frontend_icache_tag_array_tag_rdata_en;
    assign frontend_icache_tag_array_0_ext_R0_clk = frontend_icache_tag_array_tag_rdata_clk;
    assign frontend_icache_tag_array_tag_rdata_data_0 = frontend_icache_tag_array_0_ext_R0_data;
    assign frontend_icache_tag_array_0_ext_W0_addr = frontend_icache_tag_array_MPORT_addr;
    assign frontend_icache_tag_array_0_ext_W0_en = frontend_icache__GEN_1;
    assign frontend_icache_tag_array_0_ext_W0_clk = frontend_icache_tag_array_MPORT_clk;
    assign frontend_icache_tag_array_0_ext_W0_data = frontend_icache_tag_array_MPORT_data_0;
     
  assign  frontend_icache__GEN_1 = frontend_icache_tag_array_MPORT_en & frontend_icache_tag_array_MPORT_mask_0 ; 
  assign  frontend_icache__tag_rdata_WIRE = frontend_icache_io_req_bits_addr [11:6]; 
  assign  frontend_icache_tag_array_tag_rdata_en = frontend_icache_refill_done ==1'h0& frontend_icache_s0_valid ; 
  assign  frontend_icache_tag_array_tag_rdata_addr = frontend_icache__tag_rdata_WIRE ; 
    reg frontend_icache_accruedRefillError ; 
    wire frontend_icache_refillError = frontend_icache_masterNodeOut_d_bits_corrupt | frontend_icache_refill_cnt >9'h0& frontend_icache_accruedRefillError ; 
    wire[20:0] frontend_icache_enc_tag ={ frontend_icache_refillError , frontend_icache_refill_tag }; 
  assign  frontend_icache__GEN_40 = frontend_icache_enc_tag ; 
  assign  frontend_icache_tag_array_MPORT_data_0 = frontend_icache__GEN_40 ; reg[63:0] frontend_icache_vb_array ; 
    wire[127:0] frontend_icache__GEN_41 =128'h1<<{1'h0, frontend_icache_refill_idx }; 
    wire[127:0] frontend_icache__GEN_42 = frontend_icache_refill_done & frontend_icache_invalidated ==1'h0 ? {64'h0, frontend_icache_vb_array }| frontend_icache__GEN_41 :~({64'h0,~ frontend_icache_vb_array }| frontend_icache__GEN_41 ); 
    wire frontend_icache_invalidate ; reg[11:0] frontend_icache_s1s3_slaveAddr ; reg[31:0] frontend_icache_s1s3_slaveData ; 
    wire[5:0] frontend_icache_s1_idx = frontend_icache_io_s1_paddr [11:6]; 
    wire[19:0] frontend_icache_s1_tag = frontend_icache_io_s1_paddr [31:12]; 
    wire[63:0] frontend_icache__GEN_43 = frontend_icache_vb_array >>{1'h0, frontend_icache_s1_idx }; 
    wire frontend_icache_s1_vb = frontend_icache__GEN_43 [0]& frontend_icache_s1_slaveValid ==1'h0; 
    wire frontend_icache_tl_error = frontend_icache_tag_array_tag_rdata_data_0 [20]; 
    wire[19:0] frontend_icache_tag = frontend_icache_tag_array_tag_rdata_data_0 [19:0]; 
    wire frontend_icache_tagMatch = frontend_icache_s1_vb & frontend_icache_tag == frontend_icache_s1_tag ; 
    wire frontend_icache_s1_tl_error_0 = frontend_icache_tagMatch & frontend_icache_tl_error ; 
  assign  frontend_icache_s1_tag_hit_0 = frontend_icache_tagMatch | frontend_icache_scratchpadHit ; 
    wire frontend_icache__GEN_44 =(( frontend_icache_s1_valid | frontend_icache_s1_slaveValid )==1'h0|( frontend_icache_s1_tag_hit_0 & frontend_icache_s1_tag_disparity_0 ==1'h0)<=1'h1)==1'h0; 
    wire[8:0] frontend_icache_mem_idx ; 
    wire frontend_icache_wen ; 
    wire[31:0] frontend_icache__GEN_45 ; 
    wire[8:0] frontend_icache__dout_WIRE ; 
    wire[8:0] frontend_icache_data_arrays_0_MPORT_1_addr ; 
    wire[31:0] frontend_icache_data_arrays_0_MPORT_1_data_0 ; 
    wire[8:0] frontend_icache_data_arrays_0_dout_addr ; 
    wire frontend_icache_data_arrays_0_dout_en ;  
    wire[8:0] frontend_icache_data_arrays_0_0_ext_R0_addr;
    wire frontend_icache_data_arrays_0_0_ext_R0_en;
    wire frontend_icache_data_arrays_0_0_ext_R0_clk;
    wire[31:0] frontend_icache_data_arrays_0_0_ext_R0_data;
    wire[8:0] frontend_icache_data_arrays_0_0_ext_W0_addr;
    wire frontend_icache_data_arrays_0_0_ext_W0_en;
    wire frontend_icache_data_arrays_0_0_ext_W0_clk;
    wire[31:0] frontend_icache_data_arrays_0_0_ext_W0_data;
    wire[8:0] frontend_icache_data_arrays_1_0_ext_R0_addr;
    wire frontend_icache_data_arrays_1_0_ext_R0_en;
    wire frontend_icache_data_arrays_1_0_ext_R0_clk;
    wire[31:0] frontend_icache_data_arrays_1_0_ext_R0_data;
    wire[8:0] frontend_icache_data_arrays_1_0_ext_W0_addr;
    wire frontend_icache_data_arrays_1_0_ext_W0_en;
    wire frontend_icache_data_arrays_1_0_ext_W0_clk;
    wire[31:0] frontend_icache_data_arrays_1_0_ext_W0_data;

    reg[31:0] frontend_icache_data_arrays_0_0_ext_Memory [0:511]; 
    reg frontend_icache_data_arrays_0_0_ext__R0_en_d0 ; reg[8:0] frontend_icache_data_arrays_0_0_ext__R0_addr_d0 ; 
  always @( posedge  frontend_icache_data_arrays_0_0_ext_R0_clk )
         begin  
             frontend_icache_data_arrays_0_0_ext__R0_en_d0  <= frontend_icache_data_arrays_0_0_ext_R0_en ; 
             frontend_icache_data_arrays_0_0_ext__R0_addr_d0  <= frontend_icache_data_arrays_0_0_ext_R0_addr ;
         end
  always @( posedge  frontend_icache_data_arrays_0_0_ext_W0_clk )
         begin 
             if ( frontend_icache_data_arrays_0_0_ext_W0_en &1'h1) 
                 frontend_icache_data_arrays_0_0_ext_Memory  [ frontend_icache_data_arrays_0_0_ext_W0_addr ]<= frontend_icache_data_arrays_0_0_ext_W0_data ;
         end
  assign  frontend_icache_data_arrays_0_0_ext_R0_data = frontend_icache_data_arrays_0_0_ext__R0_en_d0  ?  frontend_icache_data_arrays_0_0_ext_Memory [ frontend_icache_data_arrays_0_0_ext__R0_addr_d0 ]:32'bx;
     
    wire frontend_icache_data_arrays_0_MPORT_1_en ; 
    wire frontend_icache_data_arrays_0_MPORT_1_mask_0 ; 
  assign  frontend_icache__GEN_0 = frontend_icache_data_arrays_0_MPORT_1_en & frontend_icache_data_arrays_0_MPORT_1_mask_0 ; 
    wire[8:0] frontend_icache_mem_idx_1 ; 
    wire frontend_icache_wen_1 ; 
    wire[31:0] frontend_icache__GEN_46 ; 
    wire[8:0] frontend_icache__dout_WIRE_1 ; 
    wire[8:0] frontend_icache_data_arrays_1_MPORT_2_addr ; 
    wire[31:0] frontend_icache_data_arrays_1_MPORT_2_data_0 ; 
    wire[8:0] frontend_icache_data_arrays_1_dout_1_addr ; 
    wire frontend_icache_data_arrays_1_dout_1_en ;  
    
    reg[31:0] frontend_icache_data_arrays_1_0_ext_Memory [0:511]; 
    reg frontend_icache_data_arrays_1_0_ext__R0_en_d0 ; reg[8:0] frontend_icache_data_arrays_1_0_ext__R0_addr_d0 ; 
  always @( posedge  frontend_icache_data_arrays_1_0_ext_R0_clk )
         begin  
             frontend_icache_data_arrays_1_0_ext__R0_en_d0  <= frontend_icache_data_arrays_1_0_ext_R0_en ; 
             frontend_icache_data_arrays_1_0_ext__R0_addr_d0  <= frontend_icache_data_arrays_1_0_ext_R0_addr ;
         end
  always @( posedge  frontend_icache_data_arrays_1_0_ext_W0_clk )
         begin 
             if ( frontend_icache_data_arrays_1_0_ext_W0_en &1'h1) 
                 frontend_icache_data_arrays_1_0_ext_Memory  [ frontend_icache_data_arrays_1_0_ext_W0_addr ]<= frontend_icache_data_arrays_1_0_ext_W0_data ;
         end
  assign  frontend_icache_data_arrays_1_0_ext_R0_data = frontend_icache_data_arrays_1_0_ext__R0_en_d0  ?  frontend_icache_data_arrays_1_0_ext_Memory [ frontend_icache_data_arrays_1_0_ext__R0_addr_d0 ]:32'bx;
    assign frontend_icache_data_arrays_0_0_ext_R0_addr = frontend_icache_data_arrays_0_dout_addr;
    assign frontend_icache_data_arrays_0_0_ext_R0_en = frontend_icache_data_arrays_0_dout_en;
    assign frontend_icache_data_arrays_0_0_ext_R0_clk = frontend_icache_data_arrays_0_dout_clk;
    assign frontend_icache_data_arrays_0_dout_data_0 = frontend_icache_data_arrays_0_0_ext_R0_data;
    assign frontend_icache_data_arrays_0_0_ext_W0_addr = frontend_icache_data_arrays_0_MPORT_1_addr;
    assign frontend_icache_data_arrays_0_0_ext_W0_en = frontend_icache__GEN_0;
    assign frontend_icache_data_arrays_0_0_ext_W0_clk = frontend_icache_data_arrays_0_MPORT_1_clk;
    assign frontend_icache_data_arrays_0_0_ext_W0_data = frontend_icache_data_arrays_0_MPORT_1_data_0;
    assign frontend_icache_data_arrays_1_0_ext_R0_addr = frontend_icache_data_arrays_1_dout_1_addr;
    assign frontend_icache_data_arrays_1_0_ext_R0_en = frontend_icache_data_arrays_1_dout_1_en;
    assign frontend_icache_data_arrays_1_0_ext_R0_clk = frontend_icache_data_arrays_1_dout_1_clk;
    assign frontend_icache_data_arrays_1_dout_1_data_0 = frontend_icache_data_arrays_1_0_ext_R0_data;
    assign frontend_icache_data_arrays_1_0_ext_W0_addr = frontend_icache_data_arrays_1_MPORT_2_addr;
    assign frontend_icache_data_arrays_1_0_ext_W0_en = frontend_icache__GEN;
    assign frontend_icache_data_arrays_1_0_ext_W0_clk = frontend_icache_data_arrays_1_MPORT_2_clk;
    assign frontend_icache_data_arrays_1_0_ext_W0_data = frontend_icache_data_arrays_1_MPORT_2_data_0;
     
    wire frontend_icache_data_arrays_1_MPORT_2_en ; 
    wire frontend_icache_data_arrays_1_MPORT_2_mask_0 ; 
  assign  frontend_icache__GEN = frontend_icache_data_arrays_1_MPORT_2_en & frontend_icache_data_arrays_1_MPORT_2_mask_0 ; 
    wire frontend_icache_s0_ren = frontend_icache_s0_valid & frontend_icache_io_req_bits_addr [2]==1'h0; 
  assign  frontend_icache_wen = frontend_icache_refill_one_beat & frontend_icache_invalidated ==1'h0| frontend_icache_s3_slaveValid & frontend_icache_s1s3_slaveAddr [2]==1'h0; 
  assign  frontend_icache_data_arrays_0_MPORT_1_en = frontend_icache_wen ; 
  assign  frontend_icache_mem_idx = frontend_icache_refill_one_beat  ? { frontend_icache_refill_idx ,3'h0}| frontend_icache_refill_cnt : frontend_icache_s3_slaveValid  ?  frontend_icache_s1s3_slaveAddr [11:3]: frontend_icache_io_req_bits_addr [11:3]; 
  assign  frontend_icache_data_arrays_0_MPORT_1_addr = frontend_icache_mem_idx ; 
  assign  frontend_icache__dout_WIRE = frontend_icache_mem_idx ; 
    wire[31:0] frontend_icache_data = frontend_icache_s3_slaveValid  ?  frontend_icache_s1s3_slaveData : frontend_icache_masterNodeOut_d_bits_data [31:0]; 
  assign  frontend_icache__GEN_45 = frontend_icache_data ; 
  assign  frontend_icache_data_arrays_0_MPORT_1_data_0 = frontend_icache__GEN_45 ; 
  assign  frontend_icache_data_arrays_0_MPORT_1_mask_0 = frontend_icache_way ==1'h0; 
  assign  frontend_icache_data_arrays_0_dout_en = frontend_icache_wen ==1'h0& frontend_icache_s0_ren ; 
  assign  frontend_icache_data_arrays_0_dout_addr = frontend_icache__dout_WIRE ; 
    wire[31:0] frontend_icache__GEN_47 = frontend_icache_s1_slaveValid  ? {20'h0, frontend_icache_s1s3_slaveAddr }: frontend_icache_io_s1_paddr ; 
    wire frontend_icache_s0_ren_1 = frontend_icache_s0_valid &(&( frontend_icache_io_req_bits_addr [2])); 
  assign  frontend_icache_wen_1 = frontend_icache_refill_one_beat & frontend_icache_invalidated ==1'h0| frontend_icache_s3_slaveValid &(&( frontend_icache_s1s3_slaveAddr [2])); 
  assign  frontend_icache_data_arrays_1_MPORT_2_en = frontend_icache_wen_1 ; 
  assign  frontend_icache_mem_idx_1 = frontend_icache_refill_one_beat  ? { frontend_icache_refill_idx ,3'h0}| frontend_icache_refill_cnt : frontend_icache_s3_slaveValid  ?  frontend_icache_s1s3_slaveAddr [11:3]: frontend_icache_io_req_bits_addr [11:3]; 
  assign  frontend_icache_data_arrays_1_MPORT_2_addr = frontend_icache_mem_idx_1 ; 
  assign  frontend_icache__dout_WIRE_1 = frontend_icache_mem_idx_1 ; 
    wire[31:0] frontend_icache_data_1 = frontend_icache_s3_slaveValid  ?  frontend_icache_s1s3_slaveData : frontend_icache_masterNodeOut_d_bits_data [63:32]; 
  assign  frontend_icache__GEN_46 = frontend_icache_data_1 ; 
  assign  frontend_icache_data_arrays_1_MPORT_2_data_0 = frontend_icache__GEN_46 ; 
  assign  frontend_icache_data_arrays_1_MPORT_2_mask_0 = frontend_icache_way_1 ==1'h0; 
  assign  frontend_icache_data_arrays_1_dout_1_en = frontend_icache_wen_1 ==1'h0& frontend_icache_s0_ren_1 ; 
  assign  frontend_icache_data_arrays_1_dout_1_addr = frontend_icache__dout_WIRE_1 ; 
    wire[31:0] frontend_icache__GEN_48 = frontend_icache_s1_slaveValid  ? {20'h0, frontend_icache_s1s3_slaveAddr }: frontend_icache_io_s1_paddr ; 
    wire[31:0] frontend_icache_s1_dout_0 =(&( frontend_icache__GEN_48 [2])) ?  frontend_icache_data_arrays_1_dout_1_data_0 : frontend_icache_data_arrays_0_dout_data_0 ; 
    wire frontend_icache_s1_dont_read = frontend_icache_s1_slaveValid & frontend_icache_s1s2_full_word_write ; 
    wire frontend_icache_s1_clk_en = frontend_icache_s1_valid | frontend_icache_s1_slaveValid ; 
    wire frontend_icache__GEN_49 = frontend_icache_s1_dont_read  ?  frontend_icache__s2_tag_hit_WIRE_0 : frontend_icache_s1_tag_hit_0 ; 
    reg frontend_icache_s2_tag_hit_0 ; 
    wire[32:0] frontend_icache__GEN_50 = frontend_icache_s2_slaveValid  ? {21'h0, frontend_icache_s1s3_slaveAddr }: frontend_icache_io_s2_vaddr ; 
    wire[10:0] frontend_icache_s2_scratchpad_word_addr_hi ={1'h0, frontend_icache__GEN_50 [11:2]}; 
    wire[12:0] frontend_icache_s2_scratchpad_word_addr ={ frontend_icache_s2_scratchpad_word_addr_hi ,2'h0}; reg[31:0] frontend_icache_s2_dout_0 ; 
    reg frontend_icache_s2_tag_disparity_r_0 ; 
    wire frontend_icache_s2_tag_disparity =| frontend_icache_s2_tag_disparity_r_0 ; 
    wire frontend_icache_s2_disparity = frontend_icache_s2_tag_disparity ; 
    wire frontend_icache__GEN_51 =| frontend_icache_s1_tl_error_0 ; 
    reg frontend_icache_s2_tl_error ; 
    reg frontend_icache_s2_scratchpad_hit ; 
  assign  frontend_icache_invalidate = frontend_icache_s2_valid & frontend_icache_s2_disparity  ? 1'h1: frontend_icache_io_invalidate ; 
  assign  frontend_icache_masterNodeOut_a_bits_a_address ={ frontend_icache_refill_paddr [31:6],6'h0}; 
    wire frontend_icache_masterNodeOut_a_bits_legal =({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h2000}&33'hCA012000)==33'h0&1'h1|1'h0|(({1'h0, frontend_icache_masterNodeOut_a_bits_a_address }&33'hCA012000)==33'h0|({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h10000}&33'hCA010000)==33'h0|({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h2000000}&33'hCA010000)==33'h0|({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h8000000}&33'hC8000000)==33'h0|({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h40000000}&33'hC0000000)==33'h0|({1'h0, frontend_icache_masterNodeOut_a_bits_a_address ^32'h80000000}&33'hC0000000)==33'h0)&1'h1; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_opcode = frontend_icache_masterNodeOut_a_bits_a_opcode ; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_param = frontend_icache_masterNodeOut_a_bits_a_param ; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_size = frontend_icache_masterNodeOut_a_bits_a_size ; 
    wire frontend_icache_masterNodeOut_a_bits_source = frontend_icache_masterNodeOut_a_bits_a_source ; 
    wire[31:0] frontend_icache_masterNodeOut_a_bits_address = frontend_icache_masterNodeOut_a_bits_a_address ; 
    wire[7:0] frontend_icache_masterNodeOut_a_bits_mask = frontend_icache_masterNodeOut_a_bits_a_mask ; 
    wire[63:0] frontend_icache_masterNodeOut_a_bits_data = frontend_icache_masterNodeOut_a_bits_a_data ; 
    wire frontend_icache_masterNodeOut_a_bits_corrupt = frontend_icache_masterNodeOut_a_bits_a_corrupt ; 
    wire[3:0] frontend_icache__GEN_52 =4'h1<< frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH_shiftAmount ; 
    wire[2:0] frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH = frontend_icache__GEN_52 [2:0]|3'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_size = frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH [2]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_bit = frontend_icache_masterNodeOut_a_bits_a_address [2]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_nbit = frontend_icache_masterNodeOut_a_bits_a_mask_bit ==1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq = frontend_icache_masterNodeOut_a_bits_a_mask_nbit &1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 = frontend_icache_masterNodeOut_a_bits_a_mask_bit &1'h1; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_size_1 = frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH [1]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 = frontend_icache_masterNodeOut_a_bits_a_address [1]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 = frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ==1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_2 = frontend_icache_masterNodeOut_a_bits_a_mask_eq & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_2 = frontend_icache_masterNodeOut_a_bits_a_mask_acc | frontend_icache_masterNodeOut_a_bits_a_mask_size_1 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_3 = frontend_icache_masterNodeOut_a_bits_a_mask_eq & frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_3 = frontend_icache_masterNodeOut_a_bits_a_mask_acc | frontend_icache_masterNodeOut_a_bits_a_mask_size_1 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_3 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_4 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_4 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_1 | frontend_icache_masterNodeOut_a_bits_a_mask_size_1 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_4 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_5 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_1 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_1 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_5 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_1 | frontend_icache_masterNodeOut_a_bits_a_mask_size_1 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_5 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_size_2 = frontend_icache_masterNodeOut_a_bits_a_mask_sizeOH [0]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 = frontend_icache_masterNodeOut_a_bits_a_address [0]; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_nbit_2 = frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 ==1'h0; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_6 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_2 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_6 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_2 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_6 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_7 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_2 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_7 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_2 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_7 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_8 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_3 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_8 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_3 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_8 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_9 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_3 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_9 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_3 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_9 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_10 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_4 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_10 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_4 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_10 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_11 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_4 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_11 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_4 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_11 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_12 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_5 & frontend_icache_masterNodeOut_a_bits_a_mask_nbit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_12 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_5 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_12 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_eq_13 = frontend_icache_masterNodeOut_a_bits_a_mask_eq_5 & frontend_icache_masterNodeOut_a_bits_a_mask_bit_2 ; 
    wire frontend_icache_masterNodeOut_a_bits_a_mask_acc_13 = frontend_icache_masterNodeOut_a_bits_a_mask_acc_5 | frontend_icache_masterNodeOut_a_bits_a_mask_size_2 & frontend_icache_masterNodeOut_a_bits_a_mask_eq_13 ; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_lo_lo ={ frontend_icache_masterNodeOut_a_bits_a_mask_acc_7 , frontend_icache_masterNodeOut_a_bits_a_mask_acc_6 }; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_lo_hi ={ frontend_icache_masterNodeOut_a_bits_a_mask_acc_9 , frontend_icache_masterNodeOut_a_bits_a_mask_acc_8 }; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_a_mask_lo ={ frontend_icache_masterNodeOut_a_bits_a_mask_lo_hi , frontend_icache_masterNodeOut_a_bits_a_mask_lo_lo }; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_hi_lo ={ frontend_icache_masterNodeOut_a_bits_a_mask_acc_11 , frontend_icache_masterNodeOut_a_bits_a_mask_acc_10 }; 
    wire[1:0] frontend_icache_masterNodeOut_a_bits_a_mask_hi_hi ={ frontend_icache_masterNodeOut_a_bits_a_mask_acc_13 , frontend_icache_masterNodeOut_a_bits_a_mask_acc_12 }; 
    wire[3:0] frontend_icache_masterNodeOut_a_bits_a_mask_hi ={ frontend_icache_masterNodeOut_a_bits_a_mask_hi_hi , frontend_icache_masterNodeOut_a_bits_a_mask_hi_lo }; 
  assign  frontend_icache_masterNodeOut_a_bits_a_mask ={ frontend_icache_masterNodeOut_a_bits_a_mask_hi , frontend_icache_masterNodeOut_a_bits_a_mask_lo }; 
    wire frontend_icache__GEN_53 = frontend_icache__GEN_16 ; 
    wire[2:0] frontend_icache__GEN_54 = frontend_icache__GEN_8 ; 
    wire[1:0] frontend_icache__GEN_55 = frontend_icache__GEN_6 ; 
    wire[3:0] frontend_icache__GEN_56 = frontend_icache__GEN_4 ; 
    wire frontend_icache__GEN_57 = frontend_icache__GEN_17 ; 
    wire[31:0] frontend_icache__GEN_58 = frontend_icache__GEN_2 ; 
    wire[7:0] frontend_icache__GEN_59 = frontend_icache__GEN_13 ; 
    wire[63:0] frontend_icache__GEN_60 = frontend_icache__GEN_11 ; 
    wire frontend_icache__GEN_61 = frontend_icache__GEN_18 ; 
    wire frontend_icache__GEN_62 = frontend_icache__GEN_19 ; 
    wire[2:0] frontend_icache__GEN_63 = frontend_icache__GEN_9 ; 
    wire[2:0] frontend_icache__GEN_64 = frontend_icache__GEN_10 ; 
    wire[3:0] frontend_icache__GEN_65 = frontend_icache__GEN_5 ; 
    wire frontend_icache__GEN_66 = frontend_icache__GEN_21 ; 
    wire[31:0] frontend_icache__GEN_67 = frontend_icache__GEN_3 ; 
    wire frontend_icache__GEN_68 = frontend_icache__GEN_22 ; 
    wire frontend_icache__GEN_69 = frontend_icache__GEN_23 ; 
    wire frontend_icache__GEN_70 = frontend_icache__GEN_24 ; 
    wire frontend_icache__GEN_71 = frontend_icache__GEN_25 ; 
    wire frontend_icache__GEN_72 = frontend_icache__GEN_26 ; 
    wire frontend_icache__GEN_73 = frontend_icache__GEN_27 ; 
    wire frontend_icache__GEN_74 = frontend_icache__GEN_28 ; 
    wire[63:0] frontend_icache__GEN_75 = frontend_icache__GEN_12 ; 
    wire frontend_icache__GEN_76 = frontend_icache__GEN_29 ; 
    wire frontend_icache__GEN_77 = frontend_icache__GEN_31 ; 
    wire[1:0] frontend_icache__GEN_78 = frontend_icache__GEN_7 ; 
  always @( posedge  frontend_icache_clock )
         begin 
             if ( frontend_icache_reset ==1'h0& frontend_icache__GEN_44 )
                 begin 
                     if (1)$error("Assertion failed\n    at ICache.scala:513 assert(!(s1_valid || s1_slaveValid) || PopCount(s1_tag_hit zip s1_tag_disparity map { case (h, d) => h && !d }) <= 1.U)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed\n    at ICache.scala:818 assert(!(tl_out.a.valid && addrMaybeInScratchpad(tl_out.a.bits.address)))\n");
                     if (1)$fatal;
                 end 
         end
    wire frontend_icache__GEN_79 = frontend_icache_refill_valid ==1'h0; 
    wire frontend_icache__GEN_80 = frontend_icache_s2_slaveValid ==1'h0; 
    wire frontend_icache__GEN_81 = frontend_icache_s2_tag_disparity ==1'h0; 
    wire frontend_icache__GEN_82 = frontend_icache_s2_scratchpad_hit ==1'h0; 
  always @( posedge  frontend_icache_clock )
         begin 
             if ( frontend_icache_reset )
                 begin  
                     frontend_icache_scratchpadOn  <=1'h0; 
                     frontend_icache_s1_slaveValid  <=1'h0; 
                     frontend_icache_s2_slaveValid  <=1'h0; 
                     frontend_icache_s1_valid  <=1'h0; 
                     frontend_icache_s2_valid  <=1'h0; 
                     frontend_icache_refill_valid  <=1'h0; 
                     frontend_icache_send_hint  <=1'h0; 
                     frontend_icache_hint_outstanding  <=1'h0; 
                     frontend_icache_counter  <=9'h0; 
                     frontend_icache_vb_array  <=64'h0;
                 end 
              else 
                 begin  
                     frontend_icache_s1_slaveValid  <=1'h0; 
                     frontend_icache_s2_slaveValid  <= frontend_icache_s1_slaveValid ; 
                     frontend_icache_s1_valid  <= frontend_icache_s0_valid ; 
                     frontend_icache_s2_valid  <= frontend_icache_s1_valid & frontend_icache_io_s1_kill ==1'h0;
                     if ( frontend_icache_refill_done ) 
                         frontend_icache_refill_valid  <=1'h0;
                      else 
                         if ( frontend_icache_refill_fire ) 
                             frontend_icache_refill_valid  <=1'h1;
                          else 
                             begin 
                             end 
                     if ( frontend_icache__GEN_36 )
                         begin 
                             if ( frontend_icache_first ) 
                                 frontend_icache_counter  <= frontend_icache_beats1 ;
                              else  
                                 frontend_icache_counter  <= frontend_icache_counter1 ;
                         end 
                      else 
                         begin 
                         end 
                     if ( frontend_icache_invalidate ) 
                         frontend_icache_vb_array  <=64'h0;
                      else 
                         if ( frontend_icache_refill_one_beat ) 
                             frontend_icache_vb_array  <= frontend_icache__GEN_42 [63:0];
                          else 
                             begin 
                             end 
                 end 
         end
  always @( posedge  frontend_icache_clock )
         begin  
             frontend_icache_s3_slaveValid  <=1'h0;
             if ( frontend_icache_s0_valid ) 
                 frontend_icache_s1_vaddr  <= frontend_icache_io_req_bits_addr ;
              else 
                 begin 
                 end  
             frontend_icache_s2_hit  <= frontend_icache_s1_hit ;
             if ( frontend_icache__GEN_79 ) 
                 frontend_icache_invalidated  <=1'h0;
              else 
                 if ( frontend_icache_invalidate ) 
                     frontend_icache_invalidated  <=1'h1;
                  else 
                     begin 
                     end  
             frontend_icache_s2_request_refill_REG  <= frontend_icache_s1_can_request_refill ;
             if ( frontend_icache__GEN_34 ) 
                 frontend_icache_refill_paddr  <= frontend_icache_io_s1_paddr ;
              else 
                 begin 
                 end 
             if ( frontend_icache__GEN_35 ) 
                 frontend_icache_refill_vaddr  <= frontend_icache_s1_vaddr ;
              else 
                 begin 
                 end 
             if ( frontend_icache_refill_one_beat ) 
                 frontend_icache_accruedRefillError  <= frontend_icache_refillError ;
              else 
                 begin 
                 end 
             if ( frontend_icache_s1_clk_en )
                 begin  
                     frontend_icache_s2_tag_hit_0  <= frontend_icache__GEN_49 ; 
                     frontend_icache_s2_dout_0  <= frontend_icache_s1_dout_0 ; 
                     frontend_icache_s2_tag_disparity_r_0  <= frontend_icache_s1_tag_disparity_0 ; 
                     frontend_icache_s2_tl_error  <= frontend_icache__GEN_51 ; 
                     frontend_icache_s2_scratchpad_hit  <= frontend_icache_s1_scratchpad_hit ;
                 end 
              else 
                 begin 
                 end 
         end
  assign  frontend_icache_auto_master_out_a_valid = frontend_icache_masterNodeOut_a_valid ; 
  assign  frontend_icache_auto_master_out_a_bits_opcode = frontend_icache_masterNodeOut_a_bits_opcode ; 
  assign  frontend_icache_auto_master_out_a_bits_param = frontend_icache_masterNodeOut_a_bits_param ; 
  assign  frontend_icache_auto_master_out_a_bits_size = frontend_icache_masterNodeOut_a_bits_size ; 
  assign  frontend_icache_auto_master_out_a_bits_source = frontend_icache_masterNodeOut_a_bits_source ; 
  assign  frontend_icache_auto_master_out_a_bits_address = frontend_icache_masterNodeOut_a_bits_address ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_bufferable = frontend_icache_masterNodeOut_a_bits_user_amba_prot_bufferable ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_modifiable = frontend_icache_masterNodeOut_a_bits_user_amba_prot_modifiable ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc = frontend_icache_masterNodeOut_a_bits_user_amba_prot_readalloc ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc = frontend_icache_masterNodeOut_a_bits_user_amba_prot_writealloc ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_privileged = frontend_icache_masterNodeOut_a_bits_user_amba_prot_privileged ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_secure = frontend_icache_masterNodeOut_a_bits_user_amba_prot_secure ; 
  assign  frontend_icache_auto_master_out_a_bits_user_amba_prot_fetch = frontend_icache_masterNodeOut_a_bits_user_amba_prot_fetch ; 
  assign  frontend_icache_auto_master_out_a_bits_mask = frontend_icache_masterNodeOut_a_bits_mask ; 
  assign  frontend_icache_auto_master_out_a_bits_data = frontend_icache_masterNodeOut_a_bits_data ; 
  assign  frontend_icache_auto_master_out_a_bits_corrupt = frontend_icache_masterNodeOut_a_bits_corrupt ; 
  assign  frontend_icache_auto_master_out_d_ready = frontend_icache_masterNodeOut_d_ready ; 
  assign  frontend_icache_io_req_ready = frontend_icache__io_req_ready_output ; 
  assign  frontend_icache_io_resp_valid = frontend_icache_s2_valid & frontend_icache_s2_hit ; 
  assign  frontend_icache_io_resp_bits_data = frontend_icache_s2_dout_0 ; 
  assign  frontend_icache_io_resp_bits_replay = frontend_icache_s2_disparity ; 
  assign  frontend_icache_io_resp_bits_ae = frontend_icache_s2_tl_error ; 
  assign  frontend_icache_io_errors_bus_valid = frontend_icache_masterNodeOut_d_ready & frontend_icache_masterNodeOut_d_valid &( frontend_icache_masterNodeOut_d_bits_denied | frontend_icache_masterNodeOut_d_bits_corrupt ); 
  assign  frontend_icache_io_errors_bus_bits ={ frontend_icache_refill_paddr [31:6],6'h0}; 
  assign  frontend_icache_io_perf_acquire = frontend_icache_refill_fire ; 
  assign  frontend_icache_io_keep_clock_enabled = frontend_icache_s1_valid |1'h0| frontend_icache_s2_valid | frontend_icache_refill_valid | frontend_icache_send_hint | frontend_icache_hint_outstanding ;
    assign frontend_icache_clock = frontend_clock;
    assign frontend_icache_reset = frontend_reset;
    assign frontend_icache_auto_master_out_a_ready = frontend_auto_icache_master_out_a_ready;
    assign frontend_auto_icache_master_out_a_valid = frontend_icache_auto_master_out_a_valid;
    assign frontend_auto_icache_master_out_a_bits_opcode = frontend_icache_auto_master_out_a_bits_opcode;
    assign frontend_auto_icache_master_out_a_bits_param = frontend_icache_auto_master_out_a_bits_param;
    assign frontend_auto_icache_master_out_a_bits_size = frontend_icache_auto_master_out_a_bits_size;
    assign frontend_auto_icache_master_out_a_bits_source = frontend_icache_auto_master_out_a_bits_source;
    assign frontend_auto_icache_master_out_a_bits_address = frontend_icache_auto_master_out_a_bits_address;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_bufferable = frontend_icache_auto_master_out_a_bits_user_amba_prot_bufferable;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_modifiable = frontend_icache_auto_master_out_a_bits_user_amba_prot_modifiable;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc = frontend_icache_auto_master_out_a_bits_user_amba_prot_readalloc;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc = frontend_icache_auto_master_out_a_bits_user_amba_prot_writealloc;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_privileged = frontend_icache_auto_master_out_a_bits_user_amba_prot_privileged;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_secure = frontend_icache_auto_master_out_a_bits_user_amba_prot_secure;
    assign frontend_auto_icache_master_out_a_bits_user_amba_prot_fetch = frontend_icache_auto_master_out_a_bits_user_amba_prot_fetch;
    assign frontend_auto_icache_master_out_a_bits_mask = frontend_icache_auto_master_out_a_bits_mask;
    assign frontend_auto_icache_master_out_a_bits_data = frontend_icache_auto_master_out_a_bits_data;
    assign frontend_auto_icache_master_out_a_bits_corrupt = frontend_icache_auto_master_out_a_bits_corrupt;
    assign frontend_auto_icache_master_out_d_ready = frontend_icache_auto_master_out_d_ready;
    assign frontend_icache_auto_master_out_d_valid = frontend_auto_icache_master_out_d_valid;
    assign frontend_icache_auto_master_out_d_bits_opcode = frontend_auto_icache_master_out_d_bits_opcode;
    assign frontend_icache_auto_master_out_d_bits_param = frontend_auto_icache_master_out_d_bits_param;
    assign frontend_icache_auto_master_out_d_bits_size = frontend_auto_icache_master_out_d_bits_size;
    assign frontend_icache_auto_master_out_d_bits_source = frontend_auto_icache_master_out_d_bits_source;
    assign frontend_icache_auto_master_out_d_bits_sink = frontend_auto_icache_master_out_d_bits_sink;
    assign frontend_icache_auto_master_out_d_bits_denied = frontend_auto_icache_master_out_d_bits_denied;
    assign frontend_icache_auto_master_out_d_bits_data = frontend_auto_icache_master_out_d_bits_data;
    assign frontend_icache_auto_master_out_d_bits_corrupt = frontend_auto_icache_master_out_d_bits_corrupt;
    assign frontend_icache_io_req_valid = frontend_s0_valid;
    assign frontend_icache_io_req_bits_addr = frontend___io_cpu_npc_output_32to0;
    assign frontend_icache_io_s1_paddr = frontend__tlb_io_resp_paddr;
    assign frontend_icache_io_s2_vaddr = frontend__s2_pc_32to0;
    assign frontend_icache_io_s1_kill = frontend__GEN_5;
    assign frontend_icache_io_s2_kill = frontend__GEN_4;
    assign frontend_icache_io_s2_cacheable = frontend_s2_tlb_resp_cacheable;
    assign frontend_icache_io_s2_prefetch = frontend__GEN_3;
    assign frontend__icache_io_resp_valid = frontend_icache_io_resp_valid;
    assign frontend__icache_io_resp_bits_data = frontend_icache_io_resp_bits_data;
    assign frontend__icache_io_resp_bits_replay = frontend_icache_io_resp_bits_replay;
    assign frontend__icache_io_resp_bits_ae = frontend_icache_io_resp_bits_ae;
    assign frontend_icache_io_invalidate = frontend_io_cpu_flush_icache;
    assign frontend_io_errors_bus_valid = frontend_icache_io_errors_bus_valid;
    assign frontend_io_errors_bus_bits = frontend_icache_io_errors_bus_bits;
    assign frontend_io_cpu_perf_acquire = frontend_icache_io_perf_acquire;
    assign frontend_icache_io_clock_enabled = frontend_clock_en;
      
    wire frontend_fq_clock;
    wire frontend_fq_reset;
    wire frontend_fq_io_enq_ready;
    wire frontend_fq_io_enq_valid;
    wire[1:0] frontend_fq_io_enq_bits_btb_cfiType;
    wire frontend_fq_io_enq_bits_btb_taken;
    wire[1:0] frontend_fq_io_enq_bits_btb_mask;
    wire frontend_fq_io_enq_bits_btb_bridx;
    wire[32:0] frontend_fq_io_enq_bits_btb_target;
    wire frontend_fq_io_enq_bits_btb_entry;
    wire[7:0] frontend_fq_io_enq_bits_btb_bht_history;
    wire frontend_fq_io_enq_bits_btb_bht_value;
    wire[33:0] frontend_fq_io_enq_bits_pc;
    wire[31:0] frontend_fq_io_enq_bits_data;
    wire[1:0] frontend_fq_io_enq_bits_mask;
    wire frontend_fq_io_enq_bits_xcpt_pf_inst;
    wire frontend_fq_io_enq_bits_xcpt_gf_inst;
    wire frontend_fq_io_enq_bits_xcpt_ae_inst;
    wire frontend_fq_io_enq_bits_replay;
    wire frontend_fq_io_deq_ready;
    wire frontend_fq_io_deq_valid;
    wire[1:0] frontend_fq_io_deq_bits_btb_cfiType;
    wire frontend_fq_io_deq_bits_btb_taken;
    wire[1:0] frontend_fq_io_deq_bits_btb_mask;
    wire frontend_fq_io_deq_bits_btb_bridx;
    wire[32:0] frontend_fq_io_deq_bits_btb_target;
    wire frontend_fq_io_deq_bits_btb_entry;
    wire[7:0] frontend_fq_io_deq_bits_btb_bht_history;
    wire frontend_fq_io_deq_bits_btb_bht_value;
    wire[33:0] frontend_fq_io_deq_bits_pc;
    wire[31:0] frontend_fq_io_deq_bits_data;
    wire[1:0] frontend_fq_io_deq_bits_mask;
    wire frontend_fq_io_deq_bits_xcpt_pf_inst;
    wire frontend_fq_io_deq_bits_xcpt_gf_inst;
    wire frontend_fq_io_deq_bits_xcpt_ae_inst;
    wire frontend_fq_io_deq_bits_replay;
    wire[2:0] frontend_fq_io_count;
    wire[4:0] frontend_fq_io_mask;

    wire frontend_fq__valid_WIRE_0 =1'h0; 
    wire frontend_fq__valid_WIRE_1 =1'h0; 
    wire frontend_fq__valid_WIRE_2 =1'h0; 
    wire frontend_fq__valid_WIRE_3 =1'h0; 
    wire frontend_fq__valid_WIRE_4 =1'h0; 
    reg frontend_fq_valid_0 ; 
    reg frontend_fq_valid_1 ; 
    reg frontend_fq_valid_2 ; 
    reg frontend_fq_valid_3 ; 
    reg frontend_fq_valid_4 ; reg[1:0] frontend_fq_elts_0_btb_cfiType ; 
    reg frontend_fq_elts_0_btb_taken ; reg[1:0] frontend_fq_elts_0_btb_mask ; 
    reg frontend_fq_elts_0_btb_bridx ; reg[32:0] frontend_fq_elts_0_btb_target ; 
    reg frontend_fq_elts_0_btb_entry ; reg[7:0] frontend_fq_elts_0_btb_bht_history ; 
    reg frontend_fq_elts_0_btb_bht_value ; reg[33:0] frontend_fq_elts_0_pc ; reg[31:0] frontend_fq_elts_0_data ; reg[1:0] frontend_fq_elts_0_mask ; 
    reg frontend_fq_elts_0_xcpt_pf_inst ; 
    reg frontend_fq_elts_0_xcpt_gf_inst ; 
    reg frontend_fq_elts_0_xcpt_ae_inst ; 
    reg frontend_fq_elts_0_replay ; reg[1:0] frontend_fq_elts_1_btb_cfiType ; 
    reg frontend_fq_elts_1_btb_taken ; reg[1:0] frontend_fq_elts_1_btb_mask ; 
    reg frontend_fq_elts_1_btb_bridx ; reg[32:0] frontend_fq_elts_1_btb_target ; 
    reg frontend_fq_elts_1_btb_entry ; reg[7:0] frontend_fq_elts_1_btb_bht_history ; 
    reg frontend_fq_elts_1_btb_bht_value ; reg[33:0] frontend_fq_elts_1_pc ; reg[31:0] frontend_fq_elts_1_data ; reg[1:0] frontend_fq_elts_1_mask ; 
    reg frontend_fq_elts_1_xcpt_pf_inst ; 
    reg frontend_fq_elts_1_xcpt_gf_inst ; 
    reg frontend_fq_elts_1_xcpt_ae_inst ; 
    reg frontend_fq_elts_1_replay ; reg[1:0] frontend_fq_elts_2_btb_cfiType ; 
    reg frontend_fq_elts_2_btb_taken ; reg[1:0] frontend_fq_elts_2_btb_mask ; 
    reg frontend_fq_elts_2_btb_bridx ; reg[32:0] frontend_fq_elts_2_btb_target ; 
    reg frontend_fq_elts_2_btb_entry ; reg[7:0] frontend_fq_elts_2_btb_bht_history ; 
    reg frontend_fq_elts_2_btb_bht_value ; reg[33:0] frontend_fq_elts_2_pc ; reg[31:0] frontend_fq_elts_2_data ; reg[1:0] frontend_fq_elts_2_mask ; 
    reg frontend_fq_elts_2_xcpt_pf_inst ; 
    reg frontend_fq_elts_2_xcpt_gf_inst ; 
    reg frontend_fq_elts_2_xcpt_ae_inst ; 
    reg frontend_fq_elts_2_replay ; reg[1:0] frontend_fq_elts_3_btb_cfiType ; 
    reg frontend_fq_elts_3_btb_taken ; reg[1:0] frontend_fq_elts_3_btb_mask ; 
    reg frontend_fq_elts_3_btb_bridx ; reg[32:0] frontend_fq_elts_3_btb_target ; 
    reg frontend_fq_elts_3_btb_entry ; reg[7:0] frontend_fq_elts_3_btb_bht_history ; 
    reg frontend_fq_elts_3_btb_bht_value ; reg[33:0] frontend_fq_elts_3_pc ; reg[31:0] frontend_fq_elts_3_data ; reg[1:0] frontend_fq_elts_3_mask ; 
    reg frontend_fq_elts_3_xcpt_pf_inst ; 
    reg frontend_fq_elts_3_xcpt_gf_inst ; 
    reg frontend_fq_elts_3_xcpt_ae_inst ; 
    reg frontend_fq_elts_3_replay ; reg[1:0] frontend_fq_elts_4_btb_cfiType ; 
    reg frontend_fq_elts_4_btb_taken ; reg[1:0] frontend_fq_elts_4_btb_mask ; 
    reg frontend_fq_elts_4_btb_bridx ; reg[32:0] frontend_fq_elts_4_btb_target ; 
    reg frontend_fq_elts_4_btb_entry ; reg[7:0] frontend_fq_elts_4_btb_bht_history ; 
    reg frontend_fq_elts_4_btb_bht_value ; reg[33:0] frontend_fq_elts_4_pc ; reg[31:0] frontend_fq_elts_4_data ; reg[1:0] frontend_fq_elts_4_mask ; 
    reg frontend_fq_elts_4_xcpt_pf_inst ; 
    reg frontend_fq_elts_4_xcpt_gf_inst ; 
    reg frontend_fq_elts_4_xcpt_ae_inst ; 
    reg frontend_fq_elts_4_replay ; 
    wire[1:0] frontend_fq_wdata_btb_cfiType = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_btb_taken = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_taken : frontend_fq_io_enq_bits_btb_taken ; 
    wire[1:0] frontend_fq_wdata_btb_mask = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_btb_bridx = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[32:0] frontend_fq_wdata_btb_target = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_btb_entry = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_btb_bht_history = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_btb_bht_value = frontend_fq_valid_1  ?  frontend_fq_elts_1_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[33:0] frontend_fq_wdata_pc = frontend_fq_valid_1  ?  frontend_fq_elts_1_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_data = frontend_fq_valid_1  ?  frontend_fq_elts_1_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_mask = frontend_fq_valid_1  ?  frontend_fq_elts_1_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_xcpt_pf_inst = frontend_fq_valid_1  ?  frontend_fq_elts_1_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_xcpt_gf_inst = frontend_fq_valid_1  ?  frontend_fq_elts_1_xcpt_gf_inst : frontend_fq_io_enq_bits_xcpt_gf_inst ; 
    wire frontend_fq_wdata_xcpt_ae_inst = frontend_fq_valid_1  ?  frontend_fq_elts_1_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_replay = frontend_fq_valid_1  ?  frontend_fq_elts_1_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq__io_enq_ready_output ; 
    wire frontend_fq_wen = frontend_fq_io_deq_ready  ?  frontend_fq_valid_1 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_0 |1'h0): frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_0 ==1'h0; 
    wire frontend_fq__GEN = frontend_fq_valid_1 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_0 |1'h0); 
    wire frontend_fq__GEN_0 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid | frontend_fq_valid_0 ; 
    wire[1:0] frontend_fq_wdata_1_btb_cfiType = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_1_btb_taken = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_taken : frontend_fq_io_enq_bits_btb_taken ; 
    wire[1:0] frontend_fq_wdata_1_btb_mask = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_1_btb_bridx = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[32:0] frontend_fq_wdata_1_btb_target = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_1_btb_entry = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_1_btb_bht_history = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_1_btb_bht_value = frontend_fq_valid_2  ?  frontend_fq_elts_2_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[33:0] frontend_fq_wdata_1_pc = frontend_fq_valid_2  ?  frontend_fq_elts_2_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_1_data = frontend_fq_valid_2  ?  frontend_fq_elts_2_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_1_mask = frontend_fq_valid_2  ?  frontend_fq_elts_2_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_1_xcpt_pf_inst = frontend_fq_valid_2  ?  frontend_fq_elts_2_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_1_xcpt_gf_inst = frontend_fq_valid_2  ?  frontend_fq_elts_2_xcpt_gf_inst : frontend_fq_io_enq_bits_xcpt_gf_inst ; 
    wire frontend_fq_wdata_1_xcpt_ae_inst = frontend_fq_valid_2  ?  frontend_fq_elts_2_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_1_replay = frontend_fq_valid_2  ?  frontend_fq_elts_2_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_1 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_2 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_1 |1'h0): frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_0 & frontend_fq_valid_1 ==1'h0; 
    wire frontend_fq__GEN_1 = frontend_fq_valid_2 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_1 |1'h0); 
    wire frontend_fq__GEN_2 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_0 | frontend_fq_valid_1 ; 
    wire[1:0] frontend_fq_wdata_2_btb_cfiType = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_2_btb_taken = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_taken : frontend_fq_io_enq_bits_btb_taken ; 
    wire[1:0] frontend_fq_wdata_2_btb_mask = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_2_btb_bridx = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[32:0] frontend_fq_wdata_2_btb_target = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_2_btb_entry = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_2_btb_bht_history = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_2_btb_bht_value = frontend_fq_valid_3  ?  frontend_fq_elts_3_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[33:0] frontend_fq_wdata_2_pc = frontend_fq_valid_3  ?  frontend_fq_elts_3_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_2_data = frontend_fq_valid_3  ?  frontend_fq_elts_3_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_2_mask = frontend_fq_valid_3  ?  frontend_fq_elts_3_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_2_xcpt_pf_inst = frontend_fq_valid_3  ?  frontend_fq_elts_3_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_2_xcpt_gf_inst = frontend_fq_valid_3  ?  frontend_fq_elts_3_xcpt_gf_inst : frontend_fq_io_enq_bits_xcpt_gf_inst ; 
    wire frontend_fq_wdata_2_xcpt_ae_inst = frontend_fq_valid_3  ?  frontend_fq_elts_3_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_2_replay = frontend_fq_valid_3  ?  frontend_fq_elts_3_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_2 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_3 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_2 |1'h0): frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_1 & frontend_fq_valid_2 ==1'h0; 
    wire frontend_fq__GEN_3 = frontend_fq_valid_3 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_2 |1'h0); 
    wire frontend_fq__GEN_4 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_1 | frontend_fq_valid_2 ; 
    wire[1:0] frontend_fq_wdata_3_btb_cfiType = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_cfiType : frontend_fq_io_enq_bits_btb_cfiType ; 
    wire frontend_fq_wdata_3_btb_taken = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_taken : frontend_fq_io_enq_bits_btb_taken ; 
    wire[1:0] frontend_fq_wdata_3_btb_mask = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_mask : frontend_fq_io_enq_bits_btb_mask ; 
    wire frontend_fq_wdata_3_btb_bridx = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bridx : frontend_fq_io_enq_bits_btb_bridx ; 
    wire[32:0] frontend_fq_wdata_3_btb_target = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_target : frontend_fq_io_enq_bits_btb_target ; 
    wire frontend_fq_wdata_3_btb_entry = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_entry : frontend_fq_io_enq_bits_btb_entry ; 
    wire[7:0] frontend_fq_wdata_3_btb_bht_history = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bht_history : frontend_fq_io_enq_bits_btb_bht_history ; 
    wire frontend_fq_wdata_3_btb_bht_value = frontend_fq_valid_4  ?  frontend_fq_elts_4_btb_bht_value : frontend_fq_io_enq_bits_btb_bht_value ; 
    wire[33:0] frontend_fq_wdata_3_pc = frontend_fq_valid_4  ?  frontend_fq_elts_4_pc : frontend_fq_io_enq_bits_pc ; 
    wire[31:0] frontend_fq_wdata_3_data = frontend_fq_valid_4  ?  frontend_fq_elts_4_data : frontend_fq_io_enq_bits_data ; 
    wire[1:0] frontend_fq_wdata_3_mask = frontend_fq_valid_4  ?  frontend_fq_elts_4_mask : frontend_fq_io_enq_bits_mask ; 
    wire frontend_fq_wdata_3_xcpt_pf_inst = frontend_fq_valid_4  ?  frontend_fq_elts_4_xcpt_pf_inst : frontend_fq_io_enq_bits_xcpt_pf_inst ; 
    wire frontend_fq_wdata_3_xcpt_gf_inst = frontend_fq_valid_4  ?  frontend_fq_elts_4_xcpt_gf_inst : frontend_fq_io_enq_bits_xcpt_gf_inst ; 
    wire frontend_fq_wdata_3_xcpt_ae_inst = frontend_fq_valid_4  ?  frontend_fq_elts_4_xcpt_ae_inst : frontend_fq_io_enq_bits_xcpt_ae_inst ; 
    wire frontend_fq_wdata_3_replay = frontend_fq_valid_4  ?  frontend_fq_elts_4_replay : frontend_fq_io_enq_bits_replay ; 
    wire frontend_fq_wen_3 = frontend_fq_io_deq_ready  ?  frontend_fq_valid_4 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_3 |1'h0): frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_2 & frontend_fq_valid_3 ==1'h0; 
    wire frontend_fq__GEN_5 = frontend_fq_valid_4 | frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_3 |1'h0); 
    wire frontend_fq__GEN_6 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_2 | frontend_fq_valid_3 ; 
    wire frontend_fq_wen_4 = frontend_fq_io_deq_ready  ?  frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_4 |1'h0)|1'h0: frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_3 & frontend_fq_valid_4 ==1'h0; 
    wire frontend_fq__GEN_7 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid &( frontend_fq_valid_4 |1'h0)|1'h0; 
    wire frontend_fq__GEN_8 = frontend_fq__io_enq_ready_output & frontend_fq_io_enq_valid & frontend_fq_valid_3 | frontend_fq_valid_4 ; 
  assign  frontend_fq__io_enq_ready_output = frontend_fq_valid_4 ==1'h0; 
    wire frontend_fq__GEN_9 = frontend_fq_valid_0 ==1'h0; 
    wire[1:0] frontend_fq_io_mask_lo ={ frontend_fq_valid_1 , frontend_fq_valid_0 }; 
    wire[1:0] frontend_fq_io_mask_hi_hi ={ frontend_fq_valid_4 , frontend_fq_valid_3 }; 
    wire[2:0] frontend_fq_io_mask_hi ={ frontend_fq_io_mask_hi_hi , frontend_fq_valid_2 }; 
    wire[4:0] frontend_fq__io_mask_output ={ frontend_fq_io_mask_hi , frontend_fq_io_mask_lo }; 
    wire[2:0] frontend_fq__GEN_10 ={2'h0, frontend_fq__io_mask_output [2]}+{1'h0,{1'h0, frontend_fq__io_mask_output [3]}+{1'h0, frontend_fq__io_mask_output [4]}}; 
  always @( posedge  frontend_fq_clock )
         begin 
             if ( frontend_fq_reset )
                 begin  
                     frontend_fq_valid_0  <= frontend_fq__valid_WIRE_0 ; 
                     frontend_fq_valid_1  <= frontend_fq__valid_WIRE_1 ; 
                     frontend_fq_valid_2  <= frontend_fq__valid_WIRE_2 ; 
                     frontend_fq_valid_3  <= frontend_fq__valid_WIRE_3 ; 
                     frontend_fq_valid_4  <= frontend_fq__valid_WIRE_4 ;
                 end 
              else 
                 if ( frontend_fq_io_deq_ready )
                     begin  
                         frontend_fq_valid_0  <= frontend_fq__GEN ; 
                         frontend_fq_valid_1  <= frontend_fq__GEN_1 ; 
                         frontend_fq_valid_2  <= frontend_fq__GEN_3 ; 
                         frontend_fq_valid_3  <= frontend_fq__GEN_5 ; 
                         frontend_fq_valid_4  <= frontend_fq__GEN_7 ;
                     end 
                  else 
                     begin  
                         frontend_fq_valid_0  <= frontend_fq__GEN_0 ; 
                         frontend_fq_valid_1  <= frontend_fq__GEN_2 ; 
                         frontend_fq_valid_2  <= frontend_fq__GEN_4 ; 
                         frontend_fq_valid_3  <= frontend_fq__GEN_6 ; 
                         frontend_fq_valid_4  <= frontend_fq__GEN_8 ;
                     end 
         end
  always @( posedge  frontend_fq_clock )
         begin 
             if ( frontend_fq_wen )
                 begin  
                     frontend_fq_elts_0_btb_cfiType  <= frontend_fq_wdata_btb_cfiType ; 
                     frontend_fq_elts_0_btb_taken  <= frontend_fq_wdata_btb_taken ; 
                     frontend_fq_elts_0_btb_mask  <= frontend_fq_wdata_btb_mask ; 
                     frontend_fq_elts_0_btb_bridx  <= frontend_fq_wdata_btb_bridx ; 
                     frontend_fq_elts_0_btb_target  <= frontend_fq_wdata_btb_target ; 
                     frontend_fq_elts_0_btb_entry  <= frontend_fq_wdata_btb_entry ; 
                     frontend_fq_elts_0_btb_bht_history  <= frontend_fq_wdata_btb_bht_history ; 
                     frontend_fq_elts_0_btb_bht_value  <= frontend_fq_wdata_btb_bht_value ; 
                     frontend_fq_elts_0_pc  <= frontend_fq_wdata_pc ; 
                     frontend_fq_elts_0_data  <= frontend_fq_wdata_data ; 
                     frontend_fq_elts_0_mask  <= frontend_fq_wdata_mask ; 
                     frontend_fq_elts_0_xcpt_pf_inst  <= frontend_fq_wdata_xcpt_pf_inst ; 
                     frontend_fq_elts_0_xcpt_gf_inst  <= frontend_fq_wdata_xcpt_gf_inst ; 
                     frontend_fq_elts_0_xcpt_ae_inst  <= frontend_fq_wdata_xcpt_ae_inst ; 
                     frontend_fq_elts_0_replay  <= frontend_fq_wdata_replay ;
                 end 
              else 
                 begin 
                 end 
             if ( frontend_fq_wen_1 )
                 begin  
                     frontend_fq_elts_1_btb_cfiType  <= frontend_fq_wdata_1_btb_cfiType ; 
                     frontend_fq_elts_1_btb_taken  <= frontend_fq_wdata_1_btb_taken ; 
                     frontend_fq_elts_1_btb_mask  <= frontend_fq_wdata_1_btb_mask ; 
                     frontend_fq_elts_1_btb_bridx  <= frontend_fq_wdata_1_btb_bridx ; 
                     frontend_fq_elts_1_btb_target  <= frontend_fq_wdata_1_btb_target ; 
                     frontend_fq_elts_1_btb_entry  <= frontend_fq_wdata_1_btb_entry ; 
                     frontend_fq_elts_1_btb_bht_history  <= frontend_fq_wdata_1_btb_bht_history ; 
                     frontend_fq_elts_1_btb_bht_value  <= frontend_fq_wdata_1_btb_bht_value ; 
                     frontend_fq_elts_1_pc  <= frontend_fq_wdata_1_pc ; 
                     frontend_fq_elts_1_data  <= frontend_fq_wdata_1_data ; 
                     frontend_fq_elts_1_mask  <= frontend_fq_wdata_1_mask ; 
                     frontend_fq_elts_1_xcpt_pf_inst  <= frontend_fq_wdata_1_xcpt_pf_inst ; 
                     frontend_fq_elts_1_xcpt_gf_inst  <= frontend_fq_wdata_1_xcpt_gf_inst ; 
                     frontend_fq_elts_1_xcpt_ae_inst  <= frontend_fq_wdata_1_xcpt_ae_inst ; 
                     frontend_fq_elts_1_replay  <= frontend_fq_wdata_1_replay ;
                 end 
              else 
                 begin 
                 end 
             if ( frontend_fq_wen_2 )
                 begin  
                     frontend_fq_elts_2_btb_cfiType  <= frontend_fq_wdata_2_btb_cfiType ; 
                     frontend_fq_elts_2_btb_taken  <= frontend_fq_wdata_2_btb_taken ; 
                     frontend_fq_elts_2_btb_mask  <= frontend_fq_wdata_2_btb_mask ; 
                     frontend_fq_elts_2_btb_bridx  <= frontend_fq_wdata_2_btb_bridx ; 
                     frontend_fq_elts_2_btb_target  <= frontend_fq_wdata_2_btb_target ; 
                     frontend_fq_elts_2_btb_entry  <= frontend_fq_wdata_2_btb_entry ; 
                     frontend_fq_elts_2_btb_bht_history  <= frontend_fq_wdata_2_btb_bht_history ; 
                     frontend_fq_elts_2_btb_bht_value  <= frontend_fq_wdata_2_btb_bht_value ; 
                     frontend_fq_elts_2_pc  <= frontend_fq_wdata_2_pc ; 
                     frontend_fq_elts_2_data  <= frontend_fq_wdata_2_data ; 
                     frontend_fq_elts_2_mask  <= frontend_fq_wdata_2_mask ; 
                     frontend_fq_elts_2_xcpt_pf_inst  <= frontend_fq_wdata_2_xcpt_pf_inst ; 
                     frontend_fq_elts_2_xcpt_gf_inst  <= frontend_fq_wdata_2_xcpt_gf_inst ; 
                     frontend_fq_elts_2_xcpt_ae_inst  <= frontend_fq_wdata_2_xcpt_ae_inst ; 
                     frontend_fq_elts_2_replay  <= frontend_fq_wdata_2_replay ;
                 end 
              else 
                 begin 
                 end 
             if ( frontend_fq_wen_3 )
                 begin  
                     frontend_fq_elts_3_btb_cfiType  <= frontend_fq_wdata_3_btb_cfiType ; 
                     frontend_fq_elts_3_btb_taken  <= frontend_fq_wdata_3_btb_taken ; 
                     frontend_fq_elts_3_btb_mask  <= frontend_fq_wdata_3_btb_mask ; 
                     frontend_fq_elts_3_btb_bridx  <= frontend_fq_wdata_3_btb_bridx ; 
                     frontend_fq_elts_3_btb_target  <= frontend_fq_wdata_3_btb_target ; 
                     frontend_fq_elts_3_btb_entry  <= frontend_fq_wdata_3_btb_entry ; 
                     frontend_fq_elts_3_btb_bht_history  <= frontend_fq_wdata_3_btb_bht_history ; 
                     frontend_fq_elts_3_btb_bht_value  <= frontend_fq_wdata_3_btb_bht_value ; 
                     frontend_fq_elts_3_pc  <= frontend_fq_wdata_3_pc ; 
                     frontend_fq_elts_3_data  <= frontend_fq_wdata_3_data ; 
                     frontend_fq_elts_3_mask  <= frontend_fq_wdata_3_mask ; 
                     frontend_fq_elts_3_xcpt_pf_inst  <= frontend_fq_wdata_3_xcpt_pf_inst ; 
                     frontend_fq_elts_3_xcpt_gf_inst  <= frontend_fq_wdata_3_xcpt_gf_inst ; 
                     frontend_fq_elts_3_xcpt_ae_inst  <= frontend_fq_wdata_3_xcpt_ae_inst ; 
                     frontend_fq_elts_3_replay  <= frontend_fq_wdata_3_replay ;
                 end 
              else 
                 begin 
                 end 
             if ( frontend_fq_wen_4 )
                 begin  
                     frontend_fq_elts_4_btb_cfiType  <= frontend_fq_io_enq_bits_btb_cfiType ; 
                     frontend_fq_elts_4_btb_taken  <= frontend_fq_io_enq_bits_btb_taken ; 
                     frontend_fq_elts_4_btb_mask  <= frontend_fq_io_enq_bits_btb_mask ; 
                     frontend_fq_elts_4_btb_bridx  <= frontend_fq_io_enq_bits_btb_bridx ; 
                     frontend_fq_elts_4_btb_target  <= frontend_fq_io_enq_bits_btb_target ; 
                     frontend_fq_elts_4_btb_entry  <= frontend_fq_io_enq_bits_btb_entry ; 
                     frontend_fq_elts_4_btb_bht_history  <= frontend_fq_io_enq_bits_btb_bht_history ; 
                     frontend_fq_elts_4_btb_bht_value  <= frontend_fq_io_enq_bits_btb_bht_value ; 
                     frontend_fq_elts_4_pc  <= frontend_fq_io_enq_bits_pc ; 
                     frontend_fq_elts_4_data  <= frontend_fq_io_enq_bits_data ; 
                     frontend_fq_elts_4_mask  <= frontend_fq_io_enq_bits_mask ; 
                     frontend_fq_elts_4_xcpt_pf_inst  <= frontend_fq_io_enq_bits_xcpt_pf_inst ; 
                     frontend_fq_elts_4_xcpt_gf_inst  <= frontend_fq_io_enq_bits_xcpt_gf_inst ; 
                     frontend_fq_elts_4_xcpt_ae_inst  <= frontend_fq_io_enq_bits_xcpt_ae_inst ; 
                     frontend_fq_elts_4_replay  <= frontend_fq_io_enq_bits_replay ;
                 end 
              else 
                 begin 
                 end 
         end
  assign  frontend_fq_io_enq_ready = frontend_fq__io_enq_ready_output ; 
  assign  frontend_fq_io_deq_valid = frontend_fq_io_enq_valid  ? 1'h1: frontend_fq_valid_0 ; 
  assign  frontend_fq_io_deq_bits_btb_cfiType = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_cfiType : frontend_fq_elts_0_btb_cfiType ; 
  assign  frontend_fq_io_deq_bits_btb_taken = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_taken : frontend_fq_elts_0_btb_taken ; 
  assign  frontend_fq_io_deq_bits_btb_mask = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_mask : frontend_fq_elts_0_btb_mask ; 
  assign  frontend_fq_io_deq_bits_btb_bridx = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_bridx : frontend_fq_elts_0_btb_bridx ; 
  assign  frontend_fq_io_deq_bits_btb_target = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_target : frontend_fq_elts_0_btb_target ; 
  assign  frontend_fq_io_deq_bits_btb_entry = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_entry : frontend_fq_elts_0_btb_entry ; 
  assign  frontend_fq_io_deq_bits_btb_bht_history = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_bht_history : frontend_fq_elts_0_btb_bht_history ; 
  assign  frontend_fq_io_deq_bits_btb_bht_value = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_btb_bht_value : frontend_fq_elts_0_btb_bht_value ; 
  assign  frontend_fq_io_deq_bits_pc = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_pc : frontend_fq_elts_0_pc ; 
  assign  frontend_fq_io_deq_bits_data = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_data : frontend_fq_elts_0_data ; 
  assign  frontend_fq_io_deq_bits_mask = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_mask : frontend_fq_elts_0_mask ; 
  assign  frontend_fq_io_deq_bits_xcpt_pf_inst = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_xcpt_pf_inst : frontend_fq_elts_0_xcpt_pf_inst ; 
  assign  frontend_fq_io_deq_bits_xcpt_gf_inst = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_xcpt_gf_inst : frontend_fq_elts_0_xcpt_gf_inst ; 
  assign  frontend_fq_io_deq_bits_xcpt_ae_inst = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_xcpt_ae_inst : frontend_fq_elts_0_xcpt_ae_inst ; 
  assign  frontend_fq_io_deq_bits_replay = frontend_fq__GEN_9  ?  frontend_fq_io_enq_bits_replay : frontend_fq_elts_0_replay ; 
  assign  frontend_fq_io_count ={1'h0,{1'h0, frontend_fq__io_mask_output [0]}+{1'h0, frontend_fq__io_mask_output [1]}}+{1'h0, frontend_fq__GEN_10 [1:0]}; 
  assign  frontend_fq_io_mask = frontend_fq__io_mask_output ;
    assign frontend_fq_clock = frontend_clock;
    assign frontend_fq_reset = frontend_reset|frontend_io_cpu_req_valid;
    assign frontend__fq_io_enq_ready = frontend_fq_io_enq_ready;
    assign frontend_fq_io_enq_valid = frontend__GEN_2;
    assign frontend_fq_io_enq_bits_btb_cfiType = frontend_s2_btb_resp_bits_cfiType;
    assign frontend_fq_io_enq_bits_btb_taken = frontend_s2_btb_taken;
    assign frontend_fq_io_enq_bits_btb_mask = frontend_s2_btb_resp_bits_mask;
    assign frontend_fq_io_enq_bits_btb_bridx = frontend_s2_btb_resp_bits_bridx;
    assign frontend_fq_io_enq_bits_btb_target = frontend_s2_btb_resp_bits_target;
    assign frontend_fq_io_enq_bits_btb_entry = frontend_s2_btb_resp_bits_entry;
    assign frontend_fq_io_enq_bits_btb_bht_history = frontend_s2_btb_resp_bits_bht_history;
    assign frontend_fq_io_enq_bits_btb_bht_value = frontend_s2_btb_resp_bits_bht_value;
    assign frontend_fq_io_enq_bits_pc = frontend_s2_pc;
    assign frontend_fq_io_enq_bits_data = frontend__icache_io_resp_bits_data;
    assign frontend_fq_io_enq_bits_mask = frontend__GEN_1;
    assign frontend_fq_io_enq_bits_xcpt_pf_inst = frontend_s2_tlb_resp_pf_inst;
    assign frontend_fq_io_enq_bits_xcpt_gf_inst = frontend_s2_tlb_resp_gf_inst;
    assign frontend_fq_io_enq_bits_xcpt_ae_inst = frontend__GEN;
    assign frontend_fq_io_enq_bits_replay = frontend__GEN_0;
    assign frontend_fq_io_deq_ready = frontend_io_cpu_resp_ready;
    assign frontend_io_cpu_resp_valid = frontend_fq_io_deq_valid;
    assign frontend_io_cpu_resp_bits_btb_cfiType = frontend_fq_io_deq_bits_btb_cfiType;
    assign frontend_io_cpu_resp_bits_btb_taken = frontend_fq_io_deq_bits_btb_taken;
    assign frontend_io_cpu_resp_bits_btb_mask = frontend_fq_io_deq_bits_btb_mask;
    assign frontend_io_cpu_resp_bits_btb_bridx = frontend_fq_io_deq_bits_btb_bridx;
    assign frontend_io_cpu_resp_bits_btb_target = frontend_fq_io_deq_bits_btb_target;
    assign frontend_io_cpu_resp_bits_btb_entry = frontend_fq_io_deq_bits_btb_entry;
    assign frontend_io_cpu_resp_bits_btb_bht_history = frontend_fq_io_deq_bits_btb_bht_history;
    assign frontend_io_cpu_resp_bits_btb_bht_value = frontend_fq_io_deq_bits_btb_bht_value;
    assign frontend_io_cpu_resp_bits_pc = frontend_fq_io_deq_bits_pc;
    assign frontend_io_cpu_resp_bits_data = frontend_fq_io_deq_bits_data;
    assign frontend_io_cpu_resp_bits_mask = frontend_fq_io_deq_bits_mask;
    assign frontend_io_cpu_resp_bits_xcpt_pf_inst = frontend_fq_io_deq_bits_xcpt_pf_inst;
    assign frontend_io_cpu_resp_bits_xcpt_gf_inst = frontend_fq_io_deq_bits_xcpt_gf_inst;
    assign frontend_io_cpu_resp_bits_xcpt_ae_inst = frontend_fq_io_deq_bits_xcpt_ae_inst;
    assign frontend_io_cpu_resp_bits_replay = frontend_fq_io_deq_bits_replay;
    assign frontend__fq_io_mask = frontend_fq_io_mask;
     
    reg frontend_clock_en_reg ; 
  assign  frontend_clock_en = frontend_clock_en_reg | frontend_io_cpu_might_request ; 
    wire frontend__GEN_8 =(( frontend_io_cpu_req_valid | frontend_io_cpu_sfence_valid | frontend_io_cpu_flush_icache | frontend_io_cpu_bht_update_valid | frontend_io_cpu_btb_update_valid )==1'h0| frontend_io_cpu_might_request )==1'h0;  
    wire frontend_tlb_clock;
    wire frontend_tlb_reset;
    wire frontend_tlb_io_req_ready;
    wire frontend_tlb_io_req_valid;
    wire[33:0] frontend_tlb_io_req_bits_vaddr;
    wire frontend_tlb_io_req_bits_passthrough;
    wire[1:0] frontend_tlb_io_req_bits_size;
    wire[4:0] frontend_tlb_io_req_bits_cmd;
    wire[1:0] frontend_tlb_io_req_bits_prv;
    wire frontend_tlb_io_req_bits_v;
    wire frontend_tlb_io_resp_miss;
    wire[31:0] frontend_tlb_io_resp_paddr;
    wire[33:0] frontend_tlb_io_resp_gpa;
    wire frontend_tlb_io_resp_gpa_is_pte;
    wire frontend_tlb_io_resp_pf_ld;
    wire frontend_tlb_io_resp_pf_st;
    wire frontend_tlb_io_resp_pf_inst;
    wire frontend_tlb_io_resp_gf_ld;
    wire frontend_tlb_io_resp_gf_st;
    wire frontend_tlb_io_resp_gf_inst;
    wire frontend_tlb_io_resp_ae_ld;
    wire frontend_tlb_io_resp_ae_st;
    wire frontend_tlb_io_resp_ae_inst;
    wire frontend_tlb_io_resp_ma_ld;
    wire frontend_tlb_io_resp_ma_st;
    wire frontend_tlb_io_resp_ma_inst;
    wire frontend_tlb_io_resp_cacheable;
    wire frontend_tlb_io_resp_must_alloc;
    wire frontend_tlb_io_resp_prefetchable;
    wire frontend_tlb_io_sfence_valid;
    wire frontend_tlb_io_sfence_bits_rs1;
    wire frontend_tlb_io_sfence_bits_rs2;
    wire[32:0] frontend_tlb_io_sfence_bits_addr;
    wire frontend_tlb_io_sfence_bits_asid;
    wire frontend_tlb_io_sfence_bits_hv;
    wire frontend_tlb_io_sfence_bits_hg;
    wire frontend_tlb_io_ptw_req_ready;
    wire frontend_tlb_io_ptw_req_valid;
    wire frontend_tlb_io_ptw_req_bits_valid;
    wire[20:0] frontend_tlb_io_ptw_req_bits_bits_addr;
    wire frontend_tlb_io_ptw_req_bits_bits_need_gpa;
    wire frontend_tlb_io_ptw_req_bits_bits_vstage1;
    wire frontend_tlb_io_ptw_req_bits_bits_stage2;
    wire frontend_tlb_io_ptw_resp_valid;
    wire frontend_tlb_io_ptw_resp_bits_ae_ptw;
    wire frontend_tlb_io_ptw_resp_bits_ae_final;
    wire frontend_tlb_io_ptw_resp_bits_pf;
    wire frontend_tlb_io_ptw_resp_bits_gf;
    wire frontend_tlb_io_ptw_resp_bits_hr;
    wire frontend_tlb_io_ptw_resp_bits_hw;
    wire frontend_tlb_io_ptw_resp_bits_hx;
    wire[9:0] frontend_tlb_io_ptw_resp_bits_pte_reserved_for_future;
    wire[43:0] frontend_tlb_io_ptw_resp_bits_pte_ppn;
    wire[1:0] frontend_tlb_io_ptw_resp_bits_pte_reserved_for_software;
    wire frontend_tlb_io_ptw_resp_bits_pte_d;
    wire frontend_tlb_io_ptw_resp_bits_pte_a;
    wire frontend_tlb_io_ptw_resp_bits_pte_g;
    wire frontend_tlb_io_ptw_resp_bits_pte_u;
    wire frontend_tlb_io_ptw_resp_bits_pte_x;
    wire frontend_tlb_io_ptw_resp_bits_pte_w;
    wire frontend_tlb_io_ptw_resp_bits_pte_r;
    wire frontend_tlb_io_ptw_resp_bits_pte_v;
    wire[1:0] frontend_tlb_io_ptw_resp_bits_level;
    wire frontend_tlb_io_ptw_resp_bits_fragmented_superpage;
    wire frontend_tlb_io_ptw_resp_bits_homogeneous;
    wire frontend_tlb_io_ptw_resp_bits_gpa_valid;
    wire[32:0] frontend_tlb_io_ptw_resp_bits_gpa_bits;
    wire frontend_tlb_io_ptw_resp_bits_gpa_is_pte;
    wire[3:0] frontend_tlb_io_ptw_ptbr_mode;
    wire[15:0] frontend_tlb_io_ptw_ptbr_asid;
    wire[43:0] frontend_tlb_io_ptw_ptbr_ppn;
    wire[3:0] frontend_tlb_io_ptw_hgatp_mode;
    wire[15:0] frontend_tlb_io_ptw_hgatp_asid;
    wire[43:0] frontend_tlb_io_ptw_hgatp_ppn;
    wire[3:0] frontend_tlb_io_ptw_vsatp_mode;
    wire[15:0] frontend_tlb_io_ptw_vsatp_asid;
    wire[43:0] frontend_tlb_io_ptw_vsatp_ppn;
    wire frontend_tlb_io_ptw_status_debug;
    wire frontend_tlb_io_ptw_status_cease;
    wire frontend_tlb_io_ptw_status_wfi;
    wire[31:0] frontend_tlb_io_ptw_status_isa;
    wire[1:0] frontend_tlb_io_ptw_status_dprv;
    wire frontend_tlb_io_ptw_status_dv;
    wire[1:0] frontend_tlb_io_ptw_status_prv;
    wire frontend_tlb_io_ptw_status_v;
    wire frontend_tlb_io_ptw_status_sd;
    wire[22:0] frontend_tlb_io_ptw_status_zero2;
    wire frontend_tlb_io_ptw_status_mpv;
    wire frontend_tlb_io_ptw_status_gva;
    wire frontend_tlb_io_ptw_status_mbe;
    wire frontend_tlb_io_ptw_status_sbe;
    wire[1:0] frontend_tlb_io_ptw_status_sxl;
    wire[1:0] frontend_tlb_io_ptw_status_uxl;
    wire frontend_tlb_io_ptw_status_sd_rv32;
    wire[7:0] frontend_tlb_io_ptw_status_zero1;
    wire frontend_tlb_io_ptw_status_tsr;
    wire frontend_tlb_io_ptw_status_tw;
    wire frontend_tlb_io_ptw_status_tvm;
    wire frontend_tlb_io_ptw_status_mxr;
    wire frontend_tlb_io_ptw_status_sum;
    wire frontend_tlb_io_ptw_status_mprv;
    wire[1:0] frontend_tlb_io_ptw_status_xs;
    wire[1:0] frontend_tlb_io_ptw_status_fs;
    wire[1:0] frontend_tlb_io_ptw_status_mpp;
    wire[1:0] frontend_tlb_io_ptw_status_vs;
    wire frontend_tlb_io_ptw_status_spp;
    wire frontend_tlb_io_ptw_status_mpie;
    wire frontend_tlb_io_ptw_status_ube;
    wire frontend_tlb_io_ptw_status_spie;
    wire frontend_tlb_io_ptw_status_upie;
    wire frontend_tlb_io_ptw_status_mie;
    wire frontend_tlb_io_ptw_status_hie;
    wire frontend_tlb_io_ptw_status_sie;
    wire frontend_tlb_io_ptw_status_uie;
    wire[29:0] frontend_tlb_io_ptw_hstatus_zero6;
    wire[1:0] frontend_tlb_io_ptw_hstatus_vsxl;
    wire[8:0] frontend_tlb_io_ptw_hstatus_zero5;
    wire frontend_tlb_io_ptw_hstatus_vtsr;
    wire frontend_tlb_io_ptw_hstatus_vtw;
    wire frontend_tlb_io_ptw_hstatus_vtvm;
    wire[1:0] frontend_tlb_io_ptw_hstatus_zero3;
    wire[5:0] frontend_tlb_io_ptw_hstatus_vgein;
    wire[1:0] frontend_tlb_io_ptw_hstatus_zero2;
    wire frontend_tlb_io_ptw_hstatus_hu;
    wire frontend_tlb_io_ptw_hstatus_spvp;
    wire frontend_tlb_io_ptw_hstatus_spv;
    wire frontend_tlb_io_ptw_hstatus_gva;
    wire frontend_tlb_io_ptw_hstatus_vsbe;
    wire[4:0] frontend_tlb_io_ptw_hstatus_zero1;
    wire frontend_tlb_io_ptw_gstatus_debug;
    wire frontend_tlb_io_ptw_gstatus_cease;
    wire frontend_tlb_io_ptw_gstatus_wfi;
    wire[31:0] frontend_tlb_io_ptw_gstatus_isa;
    wire[1:0] frontend_tlb_io_ptw_gstatus_dprv;
    wire frontend_tlb_io_ptw_gstatus_dv;
    wire[1:0] frontend_tlb_io_ptw_gstatus_prv;
    wire frontend_tlb_io_ptw_gstatus_v;
    wire frontend_tlb_io_ptw_gstatus_sd;
    wire[22:0] frontend_tlb_io_ptw_gstatus_zero2;
    wire frontend_tlb_io_ptw_gstatus_mpv;
    wire frontend_tlb_io_ptw_gstatus_gva;
    wire frontend_tlb_io_ptw_gstatus_mbe;
    wire frontend_tlb_io_ptw_gstatus_sbe;
    wire[1:0] frontend_tlb_io_ptw_gstatus_sxl;
    wire[1:0] frontend_tlb_io_ptw_gstatus_uxl;
    wire frontend_tlb_io_ptw_gstatus_sd_rv32;
    wire[7:0] frontend_tlb_io_ptw_gstatus_zero1;
    wire frontend_tlb_io_ptw_gstatus_tsr;
    wire frontend_tlb_io_ptw_gstatus_tw;
    wire frontend_tlb_io_ptw_gstatus_tvm;
    wire frontend_tlb_io_ptw_gstatus_mxr;
    wire frontend_tlb_io_ptw_gstatus_sum;
    wire frontend_tlb_io_ptw_gstatus_mprv;
    wire[1:0] frontend_tlb_io_ptw_gstatus_xs;
    wire[1:0] frontend_tlb_io_ptw_gstatus_fs;
    wire[1:0] frontend_tlb_io_ptw_gstatus_mpp;
    wire[1:0] frontend_tlb_io_ptw_gstatus_vs;
    wire frontend_tlb_io_ptw_gstatus_spp;
    wire frontend_tlb_io_ptw_gstatus_mpie;
    wire frontend_tlb_io_ptw_gstatus_ube;
    wire frontend_tlb_io_ptw_gstatus_spie;
    wire frontend_tlb_io_ptw_gstatus_upie;
    wire frontend_tlb_io_ptw_gstatus_mie;
    wire frontend_tlb_io_ptw_gstatus_hie;
    wire frontend_tlb_io_ptw_gstatus_sie;
    wire frontend_tlb_io_ptw_gstatus_uie;
    wire frontend_tlb_io_ptw_pmp_0_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_0_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_0_cfg_a;
    wire frontend_tlb_io_ptw_pmp_0_cfg_x;
    wire frontend_tlb_io_ptw_pmp_0_cfg_w;
    wire frontend_tlb_io_ptw_pmp_0_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_0_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_0_mask;
    wire frontend_tlb_io_ptw_pmp_1_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_1_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_1_cfg_a;
    wire frontend_tlb_io_ptw_pmp_1_cfg_x;
    wire frontend_tlb_io_ptw_pmp_1_cfg_w;
    wire frontend_tlb_io_ptw_pmp_1_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_1_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_1_mask;
    wire frontend_tlb_io_ptw_pmp_2_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_2_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_2_cfg_a;
    wire frontend_tlb_io_ptw_pmp_2_cfg_x;
    wire frontend_tlb_io_ptw_pmp_2_cfg_w;
    wire frontend_tlb_io_ptw_pmp_2_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_2_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_2_mask;
    wire frontend_tlb_io_ptw_pmp_3_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_3_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_3_cfg_a;
    wire frontend_tlb_io_ptw_pmp_3_cfg_x;
    wire frontend_tlb_io_ptw_pmp_3_cfg_w;
    wire frontend_tlb_io_ptw_pmp_3_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_3_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_3_mask;
    wire frontend_tlb_io_ptw_pmp_4_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_4_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_4_cfg_a;
    wire frontend_tlb_io_ptw_pmp_4_cfg_x;
    wire frontend_tlb_io_ptw_pmp_4_cfg_w;
    wire frontend_tlb_io_ptw_pmp_4_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_4_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_4_mask;
    wire frontend_tlb_io_ptw_pmp_5_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_5_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_5_cfg_a;
    wire frontend_tlb_io_ptw_pmp_5_cfg_x;
    wire frontend_tlb_io_ptw_pmp_5_cfg_w;
    wire frontend_tlb_io_ptw_pmp_5_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_5_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_5_mask;
    wire frontend_tlb_io_ptw_pmp_6_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_6_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_6_cfg_a;
    wire frontend_tlb_io_ptw_pmp_6_cfg_x;
    wire frontend_tlb_io_ptw_pmp_6_cfg_w;
    wire frontend_tlb_io_ptw_pmp_6_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_6_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_6_mask;
    wire frontend_tlb_io_ptw_pmp_7_cfg_l;
    wire[1:0] frontend_tlb_io_ptw_pmp_7_cfg_res;
    wire[1:0] frontend_tlb_io_ptw_pmp_7_cfg_a;
    wire frontend_tlb_io_ptw_pmp_7_cfg_x;
    wire frontend_tlb_io_ptw_pmp_7_cfg_w;
    wire frontend_tlb_io_ptw_pmp_7_cfg_r;
    wire[29:0] frontend_tlb_io_ptw_pmp_7_addr;
    wire[31:0] frontend_tlb_io_ptw_pmp_7_mask;
    wire frontend_tlb_io_ptw_customCSRs_csrs_0_ren;
    wire frontend_tlb_io_ptw_customCSRs_csrs_0_wen;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_0_wdata;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_0_value;
    wire frontend_tlb_io_ptw_customCSRs_csrs_0_stall;
    wire frontend_tlb_io_ptw_customCSRs_csrs_0_set;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_0_sdata;
    wire frontend_tlb_io_ptw_customCSRs_csrs_1_ren;
    wire frontend_tlb_io_ptw_customCSRs_csrs_1_wen;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_1_wdata;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_1_value;
    wire frontend_tlb_io_ptw_customCSRs_csrs_1_stall;
    wire frontend_tlb_io_ptw_customCSRs_csrs_1_set;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_1_sdata;
    wire frontend_tlb_io_ptw_customCSRs_csrs_2_ren;
    wire frontend_tlb_io_ptw_customCSRs_csrs_2_wen;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_2_wdata;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_2_value;
    wire frontend_tlb_io_ptw_customCSRs_csrs_2_stall;
    wire frontend_tlb_io_ptw_customCSRs_csrs_2_set;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_2_sdata;
    wire frontend_tlb_io_ptw_customCSRs_csrs_3_ren;
    wire frontend_tlb_io_ptw_customCSRs_csrs_3_wen;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_3_wdata;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_3_value;
    wire frontend_tlb_io_ptw_customCSRs_csrs_3_stall;
    wire frontend_tlb_io_ptw_customCSRs_csrs_3_set;
    wire[63:0] frontend_tlb_io_ptw_customCSRs_csrs_3_sdata;
    wire frontend_tlb_io_kill;

    wire[1:0] frontend_tlb__mpu_priv_1to0 ; 
    wire[31:0] frontend_tlb__mpu_physaddr_31to0 ; 
    wire[19:0] frontend_tlb__entries_barrier_5_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_5_io_y_u ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_5_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_5_io_y_pf ; 
    wire frontend_tlb__entries_barrier_5_io_y_gf ; 
    wire frontend_tlb__entries_barrier_5_io_y_sw ; 
    wire frontend_tlb__entries_barrier_5_io_y_sx ; 
    wire frontend_tlb__entries_barrier_5_io_y_sr ; 
    wire frontend_tlb__entries_barrier_5_io_y_hw ; 
    wire frontend_tlb__entries_barrier_5_io_y_hx ; 
    wire frontend_tlb__entries_barrier_5_io_y_hr ; 
    wire[19:0] frontend_tlb__entries_barrier_4_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_4_io_y_u ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_4_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_4_io_y_pf ; 
    wire frontend_tlb__entries_barrier_4_io_y_gf ; 
    wire frontend_tlb__entries_barrier_4_io_y_sw ; 
    wire frontend_tlb__entries_barrier_4_io_y_sx ; 
    wire frontend_tlb__entries_barrier_4_io_y_sr ; 
    wire frontend_tlb__entries_barrier_4_io_y_hw ; 
    wire frontend_tlb__entries_barrier_4_io_y_hx ; 
    wire frontend_tlb__entries_barrier_4_io_y_hr ; 
    wire frontend_tlb__entries_barrier_4_io_y_pw ; 
    wire frontend_tlb__entries_barrier_4_io_y_px ; 
    wire frontend_tlb__entries_barrier_4_io_y_pr ; 
    wire frontend_tlb__entries_barrier_4_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_4_io_y_pal ; 
    wire frontend_tlb__entries_barrier_4_io_y_paa ; 
    wire frontend_tlb__entries_barrier_4_io_y_eff ; 
    wire frontend_tlb__entries_barrier_4_io_y_c ; 
    wire[19:0] frontend_tlb__entries_barrier_3_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_3_io_y_u ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_3_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_3_io_y_pf ; 
    wire frontend_tlb__entries_barrier_3_io_y_gf ; 
    wire frontend_tlb__entries_barrier_3_io_y_sw ; 
    wire frontend_tlb__entries_barrier_3_io_y_sx ; 
    wire frontend_tlb__entries_barrier_3_io_y_sr ; 
    wire frontend_tlb__entries_barrier_3_io_y_hw ; 
    wire frontend_tlb__entries_barrier_3_io_y_hx ; 
    wire frontend_tlb__entries_barrier_3_io_y_hr ; 
    wire frontend_tlb__entries_barrier_3_io_y_pw ; 
    wire frontend_tlb__entries_barrier_3_io_y_px ; 
    wire frontend_tlb__entries_barrier_3_io_y_pr ; 
    wire frontend_tlb__entries_barrier_3_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_3_io_y_pal ; 
    wire frontend_tlb__entries_barrier_3_io_y_paa ; 
    wire frontend_tlb__entries_barrier_3_io_y_eff ; 
    wire frontend_tlb__entries_barrier_3_io_y_c ; 
    wire[19:0] frontend_tlb__entries_barrier_2_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_2_io_y_u ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_2_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_2_io_y_pf ; 
    wire frontend_tlb__entries_barrier_2_io_y_gf ; 
    wire frontend_tlb__entries_barrier_2_io_y_sw ; 
    wire frontend_tlb__entries_barrier_2_io_y_sx ; 
    wire frontend_tlb__entries_barrier_2_io_y_sr ; 
    wire frontend_tlb__entries_barrier_2_io_y_hw ; 
    wire frontend_tlb__entries_barrier_2_io_y_hx ; 
    wire frontend_tlb__entries_barrier_2_io_y_hr ; 
    wire frontend_tlb__entries_barrier_2_io_y_pw ; 
    wire frontend_tlb__entries_barrier_2_io_y_px ; 
    wire frontend_tlb__entries_barrier_2_io_y_pr ; 
    wire frontend_tlb__entries_barrier_2_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_2_io_y_pal ; 
    wire frontend_tlb__entries_barrier_2_io_y_paa ; 
    wire frontend_tlb__entries_barrier_2_io_y_eff ; 
    wire frontend_tlb__entries_barrier_2_io_y_c ; 
    wire[19:0] frontend_tlb__entries_barrier_1_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_1_io_y_u ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_1_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_1_io_y_pf ; 
    wire frontend_tlb__entries_barrier_1_io_y_gf ; 
    wire frontend_tlb__entries_barrier_1_io_y_sw ; 
    wire frontend_tlb__entries_barrier_1_io_y_sx ; 
    wire frontend_tlb__entries_barrier_1_io_y_sr ; 
    wire frontend_tlb__entries_barrier_1_io_y_hw ; 
    wire frontend_tlb__entries_barrier_1_io_y_hx ; 
    wire frontend_tlb__entries_barrier_1_io_y_hr ; 
    wire frontend_tlb__entries_barrier_1_io_y_pw ; 
    wire frontend_tlb__entries_barrier_1_io_y_px ; 
    wire frontend_tlb__entries_barrier_1_io_y_pr ; 
    wire frontend_tlb__entries_barrier_1_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_1_io_y_pal ; 
    wire frontend_tlb__entries_barrier_1_io_y_paa ; 
    wire frontend_tlb__entries_barrier_1_io_y_eff ; 
    wire frontend_tlb__entries_barrier_1_io_y_c ; 
    wire[19:0] frontend_tlb__entries_barrier_io_y_ppn ; 
    wire frontend_tlb__entries_barrier_io_y_u ; 
    wire frontend_tlb__entries_barrier_io_y_ae_ptw ; 
    wire frontend_tlb__entries_barrier_io_y_ae_final ; 
    wire frontend_tlb__entries_barrier_io_y_ae_stage2 ; 
    wire frontend_tlb__entries_barrier_io_y_pf ; 
    wire frontend_tlb__entries_barrier_io_y_gf ; 
    wire frontend_tlb__entries_barrier_io_y_sw ; 
    wire frontend_tlb__entries_barrier_io_y_sx ; 
    wire frontend_tlb__entries_barrier_io_y_sr ; 
    wire frontend_tlb__entries_barrier_io_y_hw ; 
    wire frontend_tlb__entries_barrier_io_y_hx ; 
    wire frontend_tlb__entries_barrier_io_y_hr ; 
    wire frontend_tlb__entries_barrier_io_y_pw ; 
    wire frontend_tlb__entries_barrier_io_y_px ; 
    wire frontend_tlb__entries_barrier_io_y_pr ; 
    wire frontend_tlb__entries_barrier_io_y_ppp ; 
    wire frontend_tlb__entries_barrier_io_y_pal ; 
    wire frontend_tlb__entries_barrier_io_y_paa ; 
    wire frontend_tlb__entries_barrier_io_y_eff ; 
    wire frontend_tlb__entries_barrier_io_y_c ; 
    wire frontend_tlb__pmp_io_r ; 
    wire frontend_tlb__pmp_io_w ; 
    wire frontend_tlb__pmp_io_x ; 
    wire[19:0] frontend_tlb__mpu_ppn_barrier_io_y_ppn ; 
    wire frontend_tlb_newEntry_u = frontend_tlb_io_ptw_resp_bits_pte_u ; 
    wire frontend_tlb_newEntry_ae_ptw = frontend_tlb_io_ptw_resp_bits_ae_ptw ; 
    wire frontend_tlb_newEntry_ae_final = frontend_tlb_io_ptw_resp_bits_ae_final ; 
    wire frontend_tlb_newEntry_pf = frontend_tlb_io_ptw_resp_bits_pf ; 
    wire frontend_tlb_newEntry_gf = frontend_tlb_io_ptw_resp_bits_gf ; 
    wire frontend_tlb_newEntry_hw = frontend_tlb_io_ptw_resp_bits_hw ; 
    wire frontend_tlb_newEntry_hx = frontend_tlb_io_ptw_resp_bits_hx ; 
    wire frontend_tlb_newEntry_hr = frontend_tlb_io_ptw_resp_bits_hr ; 
    wire frontend_tlb_newEntry_fragmented_superpage = frontend_tlb_io_ptw_resp_bits_fragmented_superpage ; 
    wire[5:0] frontend_tlb_stage1_bypass =6'h0; 
    wire frontend_tlb_priv_v =1'h0; 
    wire frontend_tlb_stage1_en =1'h0; 
    wire frontend_tlb_vstage1_en =1'h0; 
    wire frontend_tlb_stage2_en =1'h0; 
    wire frontend_tlb_do_refill =1'h0; 
    wire frontend_tlb_cmd_readx =1'h0; 
    wire[20:0] frontend_tlb_vpn = frontend_tlb_io_req_bits_vaddr [32:12]; reg[1:0] frontend_tlb_sectored_entries_0_0_level ; reg[20:0] frontend_tlb_sectored_entries_0_0_tag_vpn ; 
    reg frontend_tlb_sectored_entries_0_0_tag_v ; reg[41:0] frontend_tlb_sectored_entries_0_0_data_0 ; reg[41:0] frontend_tlb_sectored_entries_0_0_data_1 ; reg[41:0] frontend_tlb_sectored_entries_0_0_data_2 ; reg[41:0] frontend_tlb_sectored_entries_0_0_data_3 ; 
    reg frontend_tlb_sectored_entries_0_0_valid_0 ; 
    reg frontend_tlb_sectored_entries_0_0_valid_1 ; 
    reg frontend_tlb_sectored_entries_0_0_valid_2 ; 
    reg frontend_tlb_sectored_entries_0_0_valid_3 ; reg[1:0] frontend_tlb_superpage_entries_0_level ; reg[20:0] frontend_tlb_superpage_entries_0_tag_vpn ; 
    reg frontend_tlb_superpage_entries_0_tag_v ; reg[41:0] frontend_tlb_superpage_entries_0_data_0 ; 
    wire[41:0] frontend_tlb__entries_WIRE_3 = frontend_tlb_superpage_entries_0_data_0 ; 
    reg frontend_tlb_superpage_entries_0_valid_0 ; reg[1:0] frontend_tlb_superpage_entries_1_level ; reg[20:0] frontend_tlb_superpage_entries_1_tag_vpn ; 
    reg frontend_tlb_superpage_entries_1_tag_v ; reg[41:0] frontend_tlb_superpage_entries_1_data_0 ; 
    wire[41:0] frontend_tlb__entries_WIRE_5 = frontend_tlb_superpage_entries_1_data_0 ; 
    reg frontend_tlb_superpage_entries_1_valid_0 ; reg[1:0] frontend_tlb_superpage_entries_2_level ; reg[20:0] frontend_tlb_superpage_entries_2_tag_vpn ; 
    reg frontend_tlb_superpage_entries_2_tag_v ; reg[41:0] frontend_tlb_superpage_entries_2_data_0 ; 
    wire[41:0] frontend_tlb__entries_WIRE_7 = frontend_tlb_superpage_entries_2_data_0 ; 
    reg frontend_tlb_superpage_entries_2_valid_0 ; reg[1:0] frontend_tlb_superpage_entries_3_level ; reg[20:0] frontend_tlb_superpage_entries_3_tag_vpn ; 
    reg frontend_tlb_superpage_entries_3_tag_v ; reg[41:0] frontend_tlb_superpage_entries_3_data_0 ; 
    wire[41:0] frontend_tlb__entries_WIRE_9 = frontend_tlb_superpage_entries_3_data_0 ; 
    reg frontend_tlb_superpage_entries_3_valid_0 ; reg[1:0] frontend_tlb_special_entry_level ; reg[20:0] frontend_tlb_special_entry_tag_vpn ; 
    reg frontend_tlb_special_entry_tag_v ; reg[41:0] frontend_tlb_special_entry_data_0 ; 
    wire[41:0] frontend_tlb__mpu_ppn_WIRE_1 = frontend_tlb_special_entry_data_0 ; 
    wire[41:0] frontend_tlb__entries_WIRE_11 = frontend_tlb_special_entry_data_0 ; 
    reg frontend_tlb_special_entry_valid_0 ; reg[1:0] frontend_tlb_state ; reg[20:0] frontend_tlb_r_refill_tag ; reg[1:0] frontend_tlb_r_superpage_repl_addr ; 
    wire[1:0] frontend_tlb_waddr = frontend_tlb_r_superpage_repl_addr ; 
    reg frontend_tlb_r_sectored_hit_valid ; 
    reg frontend_tlb_r_superpage_hit_valid ; reg[1:0] frontend_tlb_r_superpage_hit_bits ; 
    reg frontend_tlb_r_vstage1_en ; 
    reg frontend_tlb_r_stage2_en ; 
    reg frontend_tlb_r_need_gpa ; 
    reg frontend_tlb_r_gpa_valid ; reg[32:0] frontend_tlb_r_gpa ; reg[20:0] frontend_tlb_r_gpa_vpn ; 
    reg frontend_tlb_r_gpa_is_pte ; 
    wire frontend_tlb_priv_s = frontend_tlb_io_req_bits_prv [0]; 
    wire frontend_tlb_priv_uses_vm = frontend_tlb_io_req_bits_prv <=2'h1; 
    wire[3:0] frontend_tlb_satp_mode = frontend_tlb_priv_v  ?  frontend_tlb_io_ptw_vsatp_mode : frontend_tlb_io_ptw_ptbr_mode ; 
    wire[15:0] frontend_tlb_satp_asid = frontend_tlb_priv_v  ?  frontend_tlb_io_ptw_vsatp_asid : frontend_tlb_io_ptw_ptbr_asid ; 
    wire[43:0] frontend_tlb_satp_ppn = frontend_tlb_priv_v  ?  frontend_tlb_io_ptw_vsatp_ppn : frontend_tlb_io_ptw_ptbr_ppn ; 
    wire frontend_tlb_vm_enabled =( frontend_tlb_stage1_en | frontend_tlb_stage2_en )& frontend_tlb_priv_uses_vm & frontend_tlb_io_req_bits_passthrough ==1'h0; 
    reg frontend_tlb_v_entries_use_stage1 ; 
    wire frontend_tlb_vsatp_mode_mismatch = frontend_tlb_priv_v & frontend_tlb_vstage1_en != frontend_tlb_v_entries_use_stage1 & frontend_tlb_io_req_bits_passthrough ==1'h0; 
    wire[19:0] frontend_tlb_refill_ppn = frontend_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire frontend_tlb_invalidate_refill = frontend_tlb_state ==2'h1|(& frontend_tlb_state )| frontend_tlb_io_sfence_valid ; 
    wire frontend_tlb__mpu_ppn_WIRE_fragmented_superpage = frontend_tlb__mpu_ppn_WIRE_1 [0]; 
    wire frontend_tlb__mpu_ppn_WIRE_c = frontend_tlb__mpu_ppn_WIRE_1 [1]; 
    wire frontend_tlb__mpu_ppn_WIRE_eff = frontend_tlb__mpu_ppn_WIRE_1 [2]; 
    wire frontend_tlb__mpu_ppn_WIRE_paa = frontend_tlb__mpu_ppn_WIRE_1 [3]; 
    wire frontend_tlb__mpu_ppn_WIRE_pal = frontend_tlb__mpu_ppn_WIRE_1 [4]; 
    wire frontend_tlb__mpu_ppn_WIRE_ppp = frontend_tlb__mpu_ppn_WIRE_1 [5]; 
    wire frontend_tlb__mpu_ppn_WIRE_pr = frontend_tlb__mpu_ppn_WIRE_1 [6]; 
    wire frontend_tlb__mpu_ppn_WIRE_px = frontend_tlb__mpu_ppn_WIRE_1 [7]; 
    wire frontend_tlb__mpu_ppn_WIRE_pw = frontend_tlb__mpu_ppn_WIRE_1 [8]; 
    wire frontend_tlb__mpu_ppn_WIRE_hr = frontend_tlb__mpu_ppn_WIRE_1 [9]; 
    wire frontend_tlb__mpu_ppn_WIRE_hx = frontend_tlb__mpu_ppn_WIRE_1 [10]; 
    wire frontend_tlb__mpu_ppn_WIRE_hw = frontend_tlb__mpu_ppn_WIRE_1 [11]; 
    wire frontend_tlb__mpu_ppn_WIRE_sr = frontend_tlb__mpu_ppn_WIRE_1 [12]; 
    wire frontend_tlb__mpu_ppn_WIRE_sx = frontend_tlb__mpu_ppn_WIRE_1 [13]; 
    wire frontend_tlb__mpu_ppn_WIRE_sw = frontend_tlb__mpu_ppn_WIRE_1 [14]; 
    wire frontend_tlb__mpu_ppn_WIRE_gf = frontend_tlb__mpu_ppn_WIRE_1 [15]; 
    wire frontend_tlb__mpu_ppn_WIRE_pf = frontend_tlb__mpu_ppn_WIRE_1 [16]; 
    wire frontend_tlb__mpu_ppn_WIRE_ae_stage2 = frontend_tlb__mpu_ppn_WIRE_1 [17]; 
    wire frontend_tlb__mpu_ppn_WIRE_ae_final = frontend_tlb__mpu_ppn_WIRE_1 [18]; 
    wire frontend_tlb__mpu_ppn_WIRE_ae_ptw = frontend_tlb__mpu_ppn_WIRE_1 [19]; 
    wire frontend_tlb__mpu_ppn_WIRE_g = frontend_tlb__mpu_ppn_WIRE_1 [20]; 
    wire frontend_tlb__mpu_ppn_WIRE_u = frontend_tlb__mpu_ppn_WIRE_1 [21]; 
    wire[19:0] frontend_tlb__mpu_ppn_WIRE_ppn = frontend_tlb__mpu_ppn_WIRE_1 [41:22];  
    wire frontend_tlb_mpu_ppn_barrier_clock;
    wire frontend_tlb_mpu_ppn_barrier_reset;
    wire[19:0] frontend_tlb_mpu_ppn_barrier_io_x_ppn;
    wire frontend_tlb_mpu_ppn_barrier_io_x_u;
    wire frontend_tlb_mpu_ppn_barrier_io_x_g;
    wire frontend_tlb_mpu_ppn_barrier_io_x_ae_ptw;
    wire frontend_tlb_mpu_ppn_barrier_io_x_ae_final;
    wire frontend_tlb_mpu_ppn_barrier_io_x_ae_stage2;
    wire frontend_tlb_mpu_ppn_barrier_io_x_pf;
    wire frontend_tlb_mpu_ppn_barrier_io_x_gf;
    wire frontend_tlb_mpu_ppn_barrier_io_x_sw;
    wire frontend_tlb_mpu_ppn_barrier_io_x_sx;
    wire frontend_tlb_mpu_ppn_barrier_io_x_sr;
    wire frontend_tlb_mpu_ppn_barrier_io_x_hw;
    wire frontend_tlb_mpu_ppn_barrier_io_x_hx;
    wire frontend_tlb_mpu_ppn_barrier_io_x_hr;
    wire frontend_tlb_mpu_ppn_barrier_io_x_pw;
    wire frontend_tlb_mpu_ppn_barrier_io_x_px;
    wire frontend_tlb_mpu_ppn_barrier_io_x_pr;
    wire frontend_tlb_mpu_ppn_barrier_io_x_ppp;
    wire frontend_tlb_mpu_ppn_barrier_io_x_pal;
    wire frontend_tlb_mpu_ppn_barrier_io_x_paa;
    wire frontend_tlb_mpu_ppn_barrier_io_x_eff;
    wire frontend_tlb_mpu_ppn_barrier_io_x_c;
    wire frontend_tlb_mpu_ppn_barrier_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_mpu_ppn_barrier_io_y_ppn;
    wire frontend_tlb_mpu_ppn_barrier_io_y_u;
    wire frontend_tlb_mpu_ppn_barrier_io_y_g;
    wire frontend_tlb_mpu_ppn_barrier_io_y_ae_ptw;
    wire frontend_tlb_mpu_ppn_barrier_io_y_ae_final;
    wire frontend_tlb_mpu_ppn_barrier_io_y_ae_stage2;
    wire frontend_tlb_mpu_ppn_barrier_io_y_pf;
    wire frontend_tlb_mpu_ppn_barrier_io_y_gf;
    wire frontend_tlb_mpu_ppn_barrier_io_y_sw;
    wire frontend_tlb_mpu_ppn_barrier_io_y_sx;
    wire frontend_tlb_mpu_ppn_barrier_io_y_sr;
    wire frontend_tlb_mpu_ppn_barrier_io_y_hw;
    wire frontend_tlb_mpu_ppn_barrier_io_y_hx;
    wire frontend_tlb_mpu_ppn_barrier_io_y_hr;
    wire frontend_tlb_mpu_ppn_barrier_io_y_pw;
    wire frontend_tlb_mpu_ppn_barrier_io_y_px;
    wire frontend_tlb_mpu_ppn_barrier_io_y_pr;
    wire frontend_tlb_mpu_ppn_barrier_io_y_ppp;
    wire frontend_tlb_mpu_ppn_barrier_io_y_pal;
    wire frontend_tlb_mpu_ppn_barrier_io_y_paa;
    wire frontend_tlb_mpu_ppn_barrier_io_y_eff;
    wire frontend_tlb_mpu_ppn_barrier_io_y_c;
    wire frontend_tlb_mpu_ppn_barrier_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_clock;
    wire frontend_tlb_entries_barrier_reset;
    wire[19:0] frontend_tlb_entries_barrier_io_x_ppn;
    wire frontend_tlb_entries_barrier_io_x_u;
    wire frontend_tlb_entries_barrier_io_x_g;
    wire frontend_tlb_entries_barrier_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_io_x_ae_final;
    wire frontend_tlb_entries_barrier_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_io_x_pf;
    wire frontend_tlb_entries_barrier_io_x_gf;
    wire frontend_tlb_entries_barrier_io_x_sw;
    wire frontend_tlb_entries_barrier_io_x_sx;
    wire frontend_tlb_entries_barrier_io_x_sr;
    wire frontend_tlb_entries_barrier_io_x_hw;
    wire frontend_tlb_entries_barrier_io_x_hx;
    wire frontend_tlb_entries_barrier_io_x_hr;
    wire frontend_tlb_entries_barrier_io_x_pw;
    wire frontend_tlb_entries_barrier_io_x_px;
    wire frontend_tlb_entries_barrier_io_x_pr;
    wire frontend_tlb_entries_barrier_io_x_ppp;
    wire frontend_tlb_entries_barrier_io_x_pal;
    wire frontend_tlb_entries_barrier_io_x_paa;
    wire frontend_tlb_entries_barrier_io_x_eff;
    wire frontend_tlb_entries_barrier_io_x_c;
    wire frontend_tlb_entries_barrier_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_io_y_ppn;
    wire frontend_tlb_entries_barrier_io_y_u;
    wire frontend_tlb_entries_barrier_io_y_g;
    wire frontend_tlb_entries_barrier_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_io_y_ae_final;
    wire frontend_tlb_entries_barrier_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_io_y_pf;
    wire frontend_tlb_entries_barrier_io_y_gf;
    wire frontend_tlb_entries_barrier_io_y_sw;
    wire frontend_tlb_entries_barrier_io_y_sx;
    wire frontend_tlb_entries_barrier_io_y_sr;
    wire frontend_tlb_entries_barrier_io_y_hw;
    wire frontend_tlb_entries_barrier_io_y_hx;
    wire frontend_tlb_entries_barrier_io_y_hr;
    wire frontend_tlb_entries_barrier_io_y_pw;
    wire frontend_tlb_entries_barrier_io_y_px;
    wire frontend_tlb_entries_barrier_io_y_pr;
    wire frontend_tlb_entries_barrier_io_y_ppp;
    wire frontend_tlb_entries_barrier_io_y_pal;
    wire frontend_tlb_entries_barrier_io_y_paa;
    wire frontend_tlb_entries_barrier_io_y_eff;
    wire frontend_tlb_entries_barrier_io_y_c;
    wire frontend_tlb_entries_barrier_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_1_clock;
    wire frontend_tlb_entries_barrier_1_reset;
    wire[19:0] frontend_tlb_entries_barrier_1_io_x_ppn;
    wire frontend_tlb_entries_barrier_1_io_x_u;
    wire frontend_tlb_entries_barrier_1_io_x_g;
    wire frontend_tlb_entries_barrier_1_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_1_io_x_ae_final;
    wire frontend_tlb_entries_barrier_1_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_1_io_x_pf;
    wire frontend_tlb_entries_barrier_1_io_x_gf;
    wire frontend_tlb_entries_barrier_1_io_x_sw;
    wire frontend_tlb_entries_barrier_1_io_x_sx;
    wire frontend_tlb_entries_barrier_1_io_x_sr;
    wire frontend_tlb_entries_barrier_1_io_x_hw;
    wire frontend_tlb_entries_barrier_1_io_x_hx;
    wire frontend_tlb_entries_barrier_1_io_x_hr;
    wire frontend_tlb_entries_barrier_1_io_x_pw;
    wire frontend_tlb_entries_barrier_1_io_x_px;
    wire frontend_tlb_entries_barrier_1_io_x_pr;
    wire frontend_tlb_entries_barrier_1_io_x_ppp;
    wire frontend_tlb_entries_barrier_1_io_x_pal;
    wire frontend_tlb_entries_barrier_1_io_x_paa;
    wire frontend_tlb_entries_barrier_1_io_x_eff;
    wire frontend_tlb_entries_barrier_1_io_x_c;
    wire frontend_tlb_entries_barrier_1_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_1_io_y_ppn;
    wire frontend_tlb_entries_barrier_1_io_y_u;
    wire frontend_tlb_entries_barrier_1_io_y_g;
    wire frontend_tlb_entries_barrier_1_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_1_io_y_ae_final;
    wire frontend_tlb_entries_barrier_1_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_1_io_y_pf;
    wire frontend_tlb_entries_barrier_1_io_y_gf;
    wire frontend_tlb_entries_barrier_1_io_y_sw;
    wire frontend_tlb_entries_barrier_1_io_y_sx;
    wire frontend_tlb_entries_barrier_1_io_y_sr;
    wire frontend_tlb_entries_barrier_1_io_y_hw;
    wire frontend_tlb_entries_barrier_1_io_y_hx;
    wire frontend_tlb_entries_barrier_1_io_y_hr;
    wire frontend_tlb_entries_barrier_1_io_y_pw;
    wire frontend_tlb_entries_barrier_1_io_y_px;
    wire frontend_tlb_entries_barrier_1_io_y_pr;
    wire frontend_tlb_entries_barrier_1_io_y_ppp;
    wire frontend_tlb_entries_barrier_1_io_y_pal;
    wire frontend_tlb_entries_barrier_1_io_y_paa;
    wire frontend_tlb_entries_barrier_1_io_y_eff;
    wire frontend_tlb_entries_barrier_1_io_y_c;
    wire frontend_tlb_entries_barrier_1_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_2_clock;
    wire frontend_tlb_entries_barrier_2_reset;
    wire[19:0] frontend_tlb_entries_barrier_2_io_x_ppn;
    wire frontend_tlb_entries_barrier_2_io_x_u;
    wire frontend_tlb_entries_barrier_2_io_x_g;
    wire frontend_tlb_entries_barrier_2_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_2_io_x_ae_final;
    wire frontend_tlb_entries_barrier_2_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_2_io_x_pf;
    wire frontend_tlb_entries_barrier_2_io_x_gf;
    wire frontend_tlb_entries_barrier_2_io_x_sw;
    wire frontend_tlb_entries_barrier_2_io_x_sx;
    wire frontend_tlb_entries_barrier_2_io_x_sr;
    wire frontend_tlb_entries_barrier_2_io_x_hw;
    wire frontend_tlb_entries_barrier_2_io_x_hx;
    wire frontend_tlb_entries_barrier_2_io_x_hr;
    wire frontend_tlb_entries_barrier_2_io_x_pw;
    wire frontend_tlb_entries_barrier_2_io_x_px;
    wire frontend_tlb_entries_barrier_2_io_x_pr;
    wire frontend_tlb_entries_barrier_2_io_x_ppp;
    wire frontend_tlb_entries_barrier_2_io_x_pal;
    wire frontend_tlb_entries_barrier_2_io_x_paa;
    wire frontend_tlb_entries_barrier_2_io_x_eff;
    wire frontend_tlb_entries_barrier_2_io_x_c;
    wire frontend_tlb_entries_barrier_2_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_2_io_y_ppn;
    wire frontend_tlb_entries_barrier_2_io_y_u;
    wire frontend_tlb_entries_barrier_2_io_y_g;
    wire frontend_tlb_entries_barrier_2_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_2_io_y_ae_final;
    wire frontend_tlb_entries_barrier_2_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_2_io_y_pf;
    wire frontend_tlb_entries_barrier_2_io_y_gf;
    wire frontend_tlb_entries_barrier_2_io_y_sw;
    wire frontend_tlb_entries_barrier_2_io_y_sx;
    wire frontend_tlb_entries_barrier_2_io_y_sr;
    wire frontend_tlb_entries_barrier_2_io_y_hw;
    wire frontend_tlb_entries_barrier_2_io_y_hx;
    wire frontend_tlb_entries_barrier_2_io_y_hr;
    wire frontend_tlb_entries_barrier_2_io_y_pw;
    wire frontend_tlb_entries_barrier_2_io_y_px;
    wire frontend_tlb_entries_barrier_2_io_y_pr;
    wire frontend_tlb_entries_barrier_2_io_y_ppp;
    wire frontend_tlb_entries_barrier_2_io_y_pal;
    wire frontend_tlb_entries_barrier_2_io_y_paa;
    wire frontend_tlb_entries_barrier_2_io_y_eff;
    wire frontend_tlb_entries_barrier_2_io_y_c;
    wire frontend_tlb_entries_barrier_2_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_3_clock;
    wire frontend_tlb_entries_barrier_3_reset;
    wire[19:0] frontend_tlb_entries_barrier_3_io_x_ppn;
    wire frontend_tlb_entries_barrier_3_io_x_u;
    wire frontend_tlb_entries_barrier_3_io_x_g;
    wire frontend_tlb_entries_barrier_3_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_3_io_x_ae_final;
    wire frontend_tlb_entries_barrier_3_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_3_io_x_pf;
    wire frontend_tlb_entries_barrier_3_io_x_gf;
    wire frontend_tlb_entries_barrier_3_io_x_sw;
    wire frontend_tlb_entries_barrier_3_io_x_sx;
    wire frontend_tlb_entries_barrier_3_io_x_sr;
    wire frontend_tlb_entries_barrier_3_io_x_hw;
    wire frontend_tlb_entries_barrier_3_io_x_hx;
    wire frontend_tlb_entries_barrier_3_io_x_hr;
    wire frontend_tlb_entries_barrier_3_io_x_pw;
    wire frontend_tlb_entries_barrier_3_io_x_px;
    wire frontend_tlb_entries_barrier_3_io_x_pr;
    wire frontend_tlb_entries_barrier_3_io_x_ppp;
    wire frontend_tlb_entries_barrier_3_io_x_pal;
    wire frontend_tlb_entries_barrier_3_io_x_paa;
    wire frontend_tlb_entries_barrier_3_io_x_eff;
    wire frontend_tlb_entries_barrier_3_io_x_c;
    wire frontend_tlb_entries_barrier_3_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_3_io_y_ppn;
    wire frontend_tlb_entries_barrier_3_io_y_u;
    wire frontend_tlb_entries_barrier_3_io_y_g;
    wire frontend_tlb_entries_barrier_3_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_3_io_y_ae_final;
    wire frontend_tlb_entries_barrier_3_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_3_io_y_pf;
    wire frontend_tlb_entries_barrier_3_io_y_gf;
    wire frontend_tlb_entries_barrier_3_io_y_sw;
    wire frontend_tlb_entries_barrier_3_io_y_sx;
    wire frontend_tlb_entries_barrier_3_io_y_sr;
    wire frontend_tlb_entries_barrier_3_io_y_hw;
    wire frontend_tlb_entries_barrier_3_io_y_hx;
    wire frontend_tlb_entries_barrier_3_io_y_hr;
    wire frontend_tlb_entries_barrier_3_io_y_pw;
    wire frontend_tlb_entries_barrier_3_io_y_px;
    wire frontend_tlb_entries_barrier_3_io_y_pr;
    wire frontend_tlb_entries_barrier_3_io_y_ppp;
    wire frontend_tlb_entries_barrier_3_io_y_pal;
    wire frontend_tlb_entries_barrier_3_io_y_paa;
    wire frontend_tlb_entries_barrier_3_io_y_eff;
    wire frontend_tlb_entries_barrier_3_io_y_c;
    wire frontend_tlb_entries_barrier_3_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_4_clock;
    wire frontend_tlb_entries_barrier_4_reset;
    wire[19:0] frontend_tlb_entries_barrier_4_io_x_ppn;
    wire frontend_tlb_entries_barrier_4_io_x_u;
    wire frontend_tlb_entries_barrier_4_io_x_g;
    wire frontend_tlb_entries_barrier_4_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_4_io_x_ae_final;
    wire frontend_tlb_entries_barrier_4_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_4_io_x_pf;
    wire frontend_tlb_entries_barrier_4_io_x_gf;
    wire frontend_tlb_entries_barrier_4_io_x_sw;
    wire frontend_tlb_entries_barrier_4_io_x_sx;
    wire frontend_tlb_entries_barrier_4_io_x_sr;
    wire frontend_tlb_entries_barrier_4_io_x_hw;
    wire frontend_tlb_entries_barrier_4_io_x_hx;
    wire frontend_tlb_entries_barrier_4_io_x_hr;
    wire frontend_tlb_entries_barrier_4_io_x_pw;
    wire frontend_tlb_entries_barrier_4_io_x_px;
    wire frontend_tlb_entries_barrier_4_io_x_pr;
    wire frontend_tlb_entries_barrier_4_io_x_ppp;
    wire frontend_tlb_entries_barrier_4_io_x_pal;
    wire frontend_tlb_entries_barrier_4_io_x_paa;
    wire frontend_tlb_entries_barrier_4_io_x_eff;
    wire frontend_tlb_entries_barrier_4_io_x_c;
    wire frontend_tlb_entries_barrier_4_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_4_io_y_ppn;
    wire frontend_tlb_entries_barrier_4_io_y_u;
    wire frontend_tlb_entries_barrier_4_io_y_g;
    wire frontend_tlb_entries_barrier_4_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_4_io_y_ae_final;
    wire frontend_tlb_entries_barrier_4_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_4_io_y_pf;
    wire frontend_tlb_entries_barrier_4_io_y_gf;
    wire frontend_tlb_entries_barrier_4_io_y_sw;
    wire frontend_tlb_entries_barrier_4_io_y_sx;
    wire frontend_tlb_entries_barrier_4_io_y_sr;
    wire frontend_tlb_entries_barrier_4_io_y_hw;
    wire frontend_tlb_entries_barrier_4_io_y_hx;
    wire frontend_tlb_entries_barrier_4_io_y_hr;
    wire frontend_tlb_entries_barrier_4_io_y_pw;
    wire frontend_tlb_entries_barrier_4_io_y_px;
    wire frontend_tlb_entries_barrier_4_io_y_pr;
    wire frontend_tlb_entries_barrier_4_io_y_ppp;
    wire frontend_tlb_entries_barrier_4_io_y_pal;
    wire frontend_tlb_entries_barrier_4_io_y_paa;
    wire frontend_tlb_entries_barrier_4_io_y_eff;
    wire frontend_tlb_entries_barrier_4_io_y_c;
    wire frontend_tlb_entries_barrier_4_io_y_fragmented_superpage;
    wire frontend_tlb_entries_barrier_5_clock;
    wire frontend_tlb_entries_barrier_5_reset;
    wire[19:0] frontend_tlb_entries_barrier_5_io_x_ppn;
    wire frontend_tlb_entries_barrier_5_io_x_u;
    wire frontend_tlb_entries_barrier_5_io_x_g;
    wire frontend_tlb_entries_barrier_5_io_x_ae_ptw;
    wire frontend_tlb_entries_barrier_5_io_x_ae_final;
    wire frontend_tlb_entries_barrier_5_io_x_ae_stage2;
    wire frontend_tlb_entries_barrier_5_io_x_pf;
    wire frontend_tlb_entries_barrier_5_io_x_gf;
    wire frontend_tlb_entries_barrier_5_io_x_sw;
    wire frontend_tlb_entries_barrier_5_io_x_sx;
    wire frontend_tlb_entries_barrier_5_io_x_sr;
    wire frontend_tlb_entries_barrier_5_io_x_hw;
    wire frontend_tlb_entries_barrier_5_io_x_hx;
    wire frontend_tlb_entries_barrier_5_io_x_hr;
    wire frontend_tlb_entries_barrier_5_io_x_pw;
    wire frontend_tlb_entries_barrier_5_io_x_px;
    wire frontend_tlb_entries_barrier_5_io_x_pr;
    wire frontend_tlb_entries_barrier_5_io_x_ppp;
    wire frontend_tlb_entries_barrier_5_io_x_pal;
    wire frontend_tlb_entries_barrier_5_io_x_paa;
    wire frontend_tlb_entries_barrier_5_io_x_eff;
    wire frontend_tlb_entries_barrier_5_io_x_c;
    wire frontend_tlb_entries_barrier_5_io_x_fragmented_superpage;
    wire[19:0] frontend_tlb_entries_barrier_5_io_y_ppn;
    wire frontend_tlb_entries_barrier_5_io_y_u;
    wire frontend_tlb_entries_barrier_5_io_y_g;
    wire frontend_tlb_entries_barrier_5_io_y_ae_ptw;
    wire frontend_tlb_entries_barrier_5_io_y_ae_final;
    wire frontend_tlb_entries_barrier_5_io_y_ae_stage2;
    wire frontend_tlb_entries_barrier_5_io_y_pf;
    wire frontend_tlb_entries_barrier_5_io_y_gf;
    wire frontend_tlb_entries_barrier_5_io_y_sw;
    wire frontend_tlb_entries_barrier_5_io_y_sx;
    wire frontend_tlb_entries_barrier_5_io_y_sr;
    wire frontend_tlb_entries_barrier_5_io_y_hw;
    wire frontend_tlb_entries_barrier_5_io_y_hx;
    wire frontend_tlb_entries_barrier_5_io_y_hr;
    wire frontend_tlb_entries_barrier_5_io_y_pw;
    wire frontend_tlb_entries_barrier_5_io_y_px;
    wire frontend_tlb_entries_barrier_5_io_y_pr;
    wire frontend_tlb_entries_barrier_5_io_y_ppp;
    wire frontend_tlb_entries_barrier_5_io_y_pal;
    wire frontend_tlb_entries_barrier_5_io_y_paa;
    wire frontend_tlb_entries_barrier_5_io_y_eff;
    wire frontend_tlb_entries_barrier_5_io_y_c;
    wire frontend_tlb_entries_barrier_5_io_y_fragmented_superpage;

    assign  frontend_tlb_mpu_ppn_barrier_io_y_ppn = frontend_tlb_mpu_ppn_barrier_io_x_ppn ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_u = frontend_tlb_mpu_ppn_barrier_io_x_u ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_g = frontend_tlb_mpu_ppn_barrier_io_x_g ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_ae_ptw = frontend_tlb_mpu_ppn_barrier_io_x_ae_ptw ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_ae_final = frontend_tlb_mpu_ppn_barrier_io_x_ae_final ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_ae_stage2 = frontend_tlb_mpu_ppn_barrier_io_x_ae_stage2 ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_pf = frontend_tlb_mpu_ppn_barrier_io_x_pf ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_gf = frontend_tlb_mpu_ppn_barrier_io_x_gf ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_sw = frontend_tlb_mpu_ppn_barrier_io_x_sw ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_sx = frontend_tlb_mpu_ppn_barrier_io_x_sx ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_sr = frontend_tlb_mpu_ppn_barrier_io_x_sr ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_hw = frontend_tlb_mpu_ppn_barrier_io_x_hw ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_hx = frontend_tlb_mpu_ppn_barrier_io_x_hx ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_hr = frontend_tlb_mpu_ppn_barrier_io_x_hr ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_pw = frontend_tlb_mpu_ppn_barrier_io_x_pw ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_px = frontend_tlb_mpu_ppn_barrier_io_x_px ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_pr = frontend_tlb_mpu_ppn_barrier_io_x_pr ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_ppp = frontend_tlb_mpu_ppn_barrier_io_x_ppp ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_pal = frontend_tlb_mpu_ppn_barrier_io_x_pal ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_paa = frontend_tlb_mpu_ppn_barrier_io_x_paa ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_eff = frontend_tlb_mpu_ppn_barrier_io_x_eff ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_c = frontend_tlb_mpu_ppn_barrier_io_x_c ; 
  assign  frontend_tlb_mpu_ppn_barrier_io_y_fragmented_superpage = frontend_tlb_mpu_ppn_barrier_io_x_fragmented_superpage ;
     
    wire[21:0] frontend_tlb_mpu_ppn = frontend_tlb_do_refill  ? {2'h0, frontend_tlb_refill_ppn }: frontend_tlb_vm_enabled  ? {2'h0, frontend_tlb__mpu_ppn_barrier_io_y_ppn }: frontend_tlb_io_req_bits_vaddr [33:12]; 
    wire[33:0] frontend_tlb_mpu_physaddr ={ frontend_tlb_mpu_ppn , frontend_tlb_io_req_bits_vaddr [11:0]}; 
    wire[2:0] frontend_tlb_mpu_priv ={ frontend_tlb_io_ptw_status_debug , frontend_tlb_io_req_bits_prv };  
    wire frontend_tlb_pmp_clock;
    wire frontend_tlb_pmp_reset;
    wire[1:0] frontend_tlb_pmp_io_prv;
    wire frontend_tlb_pmp_io_pmp_0_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_0_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_0_cfg_a;
    wire frontend_tlb_pmp_io_pmp_0_cfg_x;
    wire frontend_tlb_pmp_io_pmp_0_cfg_w;
    wire frontend_tlb_pmp_io_pmp_0_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_0_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_0_mask;
    wire frontend_tlb_pmp_io_pmp_1_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_1_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_1_cfg_a;
    wire frontend_tlb_pmp_io_pmp_1_cfg_x;
    wire frontend_tlb_pmp_io_pmp_1_cfg_w;
    wire frontend_tlb_pmp_io_pmp_1_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_1_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_1_mask;
    wire frontend_tlb_pmp_io_pmp_2_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_2_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_2_cfg_a;
    wire frontend_tlb_pmp_io_pmp_2_cfg_x;
    wire frontend_tlb_pmp_io_pmp_2_cfg_w;
    wire frontend_tlb_pmp_io_pmp_2_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_2_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_2_mask;
    wire frontend_tlb_pmp_io_pmp_3_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_3_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_3_cfg_a;
    wire frontend_tlb_pmp_io_pmp_3_cfg_x;
    wire frontend_tlb_pmp_io_pmp_3_cfg_w;
    wire frontend_tlb_pmp_io_pmp_3_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_3_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_3_mask;
    wire frontend_tlb_pmp_io_pmp_4_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_4_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_4_cfg_a;
    wire frontend_tlb_pmp_io_pmp_4_cfg_x;
    wire frontend_tlb_pmp_io_pmp_4_cfg_w;
    wire frontend_tlb_pmp_io_pmp_4_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_4_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_4_mask;
    wire frontend_tlb_pmp_io_pmp_5_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_5_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_5_cfg_a;
    wire frontend_tlb_pmp_io_pmp_5_cfg_x;
    wire frontend_tlb_pmp_io_pmp_5_cfg_w;
    wire frontend_tlb_pmp_io_pmp_5_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_5_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_5_mask;
    wire frontend_tlb_pmp_io_pmp_6_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_6_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_6_cfg_a;
    wire frontend_tlb_pmp_io_pmp_6_cfg_x;
    wire frontend_tlb_pmp_io_pmp_6_cfg_w;
    wire frontend_tlb_pmp_io_pmp_6_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_6_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_6_mask;
    wire frontend_tlb_pmp_io_pmp_7_cfg_l;
    wire[1:0] frontend_tlb_pmp_io_pmp_7_cfg_res;
    wire[1:0] frontend_tlb_pmp_io_pmp_7_cfg_a;
    wire frontend_tlb_pmp_io_pmp_7_cfg_x;
    wire frontend_tlb_pmp_io_pmp_7_cfg_w;
    wire frontend_tlb_pmp_io_pmp_7_cfg_r;
    wire[29:0] frontend_tlb_pmp_io_pmp_7_addr;
    wire[31:0] frontend_tlb_pmp_io_pmp_7_mask;
    wire[31:0] frontend_tlb_pmp_io_addr;
    wire[1:0] frontend_tlb_pmp_io_size;
    wire frontend_tlb_pmp_io_r;
    wire frontend_tlb_pmp_io_w;
    wire frontend_tlb_pmp_io_x;

    wire frontend_tlb_pmp_res_cur_cfg_l = frontend_tlb_pmp_io_pmp_7_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_cfg_res = frontend_tlb_pmp_io_pmp_7_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_cfg_a = frontend_tlb_pmp_io_pmp_7_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_addr = frontend_tlb_pmp_io_pmp_7_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_mask = frontend_tlb_pmp_io_pmp_7_mask ; 
    wire frontend_tlb_pmp_res_cur_1_cfg_l = frontend_tlb_pmp_io_pmp_6_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_1_cfg_res = frontend_tlb_pmp_io_pmp_6_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_1_cfg_a = frontend_tlb_pmp_io_pmp_6_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_1_addr = frontend_tlb_pmp_io_pmp_6_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_1_mask = frontend_tlb_pmp_io_pmp_6_mask ; 
    wire frontend_tlb_pmp_res_cur_2_cfg_l = frontend_tlb_pmp_io_pmp_5_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_2_cfg_res = frontend_tlb_pmp_io_pmp_5_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_2_cfg_a = frontend_tlb_pmp_io_pmp_5_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_2_addr = frontend_tlb_pmp_io_pmp_5_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_2_mask = frontend_tlb_pmp_io_pmp_5_mask ; 
    wire frontend_tlb_pmp_res_cur_3_cfg_l = frontend_tlb_pmp_io_pmp_4_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_3_cfg_res = frontend_tlb_pmp_io_pmp_4_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_3_cfg_a = frontend_tlb_pmp_io_pmp_4_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_3_addr = frontend_tlb_pmp_io_pmp_4_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_3_mask = frontend_tlb_pmp_io_pmp_4_mask ; 
    wire frontend_tlb_pmp_res_cur_4_cfg_l = frontend_tlb_pmp_io_pmp_3_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_4_cfg_res = frontend_tlb_pmp_io_pmp_3_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_4_cfg_a = frontend_tlb_pmp_io_pmp_3_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_4_addr = frontend_tlb_pmp_io_pmp_3_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_4_mask = frontend_tlb_pmp_io_pmp_3_mask ; 
    wire frontend_tlb_pmp_res_cur_5_cfg_l = frontend_tlb_pmp_io_pmp_2_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_5_cfg_res = frontend_tlb_pmp_io_pmp_2_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_5_cfg_a = frontend_tlb_pmp_io_pmp_2_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_5_addr = frontend_tlb_pmp_io_pmp_2_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_5_mask = frontend_tlb_pmp_io_pmp_2_mask ; 
    wire frontend_tlb_pmp_res_cur_6_cfg_l = frontend_tlb_pmp_io_pmp_1_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_6_cfg_res = frontend_tlb_pmp_io_pmp_1_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_6_cfg_a = frontend_tlb_pmp_io_pmp_1_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_6_addr = frontend_tlb_pmp_io_pmp_1_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_6_mask = frontend_tlb_pmp_io_pmp_1_mask ; 
    wire frontend_tlb_pmp_res_cur_7_cfg_l = frontend_tlb_pmp_io_pmp_0_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cur_7_cfg_res = frontend_tlb_pmp_io_pmp_0_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cur_7_cfg_a = frontend_tlb_pmp_io_pmp_0_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_res_cur_7_addr = frontend_tlb_pmp_io_pmp_0_addr ; 
    wire[31:0] frontend_tlb_pmp_res_cur_7_mask = frontend_tlb_pmp_io_pmp_0_mask ; 
    wire[1:0] frontend_tlb_pmp__pmp0_WIRE_cfg_res =2'h0; 
    wire[1:0] frontend_tlb_pmp__pmp0_WIRE_cfg_a =2'h0; 
    wire[29:0] frontend_tlb_pmp__pmp0_WIRE_addr =30'h0; 
    wire[31:0] frontend_tlb_pmp__pmp0_WIRE_mask =32'h0; 
    wire frontend_tlb_pmp__pmp0_WIRE_cfg_l =1'h0; 
    wire frontend_tlb_pmp__pmp0_WIRE_cfg_x =1'h0; 
    wire frontend_tlb_pmp__pmp0_WIRE_cfg_w =1'h0; 
    wire frontend_tlb_pmp__pmp0_WIRE_cfg_r =1'h0; 
    wire frontend_tlb_pmp_default_0 = frontend_tlb_pmp_io_prv >2'h1; 
    wire frontend_tlb_pmp_pmp0_cfg_x = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_pmp0_cfg_w = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_pmp0_cfg_r = frontend_tlb_pmp_default_0 ; 
    wire frontend_tlb_pmp_pmp0_cfg_l = frontend_tlb_pmp__pmp0_WIRE_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_pmp0_cfg_res = frontend_tlb_pmp__pmp0_WIRE_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_pmp0_cfg_a = frontend_tlb_pmp__pmp0_WIRE_cfg_a ; 
    wire[29:0] frontend_tlb_pmp_pmp0_addr = frontend_tlb_pmp__pmp0_WIRE_addr ; 
    wire[31:0] frontend_tlb_pmp_pmp0_mask = frontend_tlb_pmp__pmp0_WIRE_mask ; 
    wire[4:0] frontend_tlb_pmp__GEN =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit = frontend_tlb_pmp_io_pmp_7_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_7_mask )==32'h0: frontend_tlb_pmp_io_pmp_7_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_7_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_7_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_1 ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_2 ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_3 ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_4 ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_5 ={ frontend_tlb_pmp_io_pmp_7_cfg_x , frontend_tlb_pmp_io_pmp_7_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_cfg_r =( frontend_tlb_pmp_io_pmp_7_cfg_r | frontend_tlb_pmp_res_ignore )&1'h1; 
    wire frontend_tlb_pmp_res_cur_cfg_w =( frontend_tlb_pmp_io_pmp_7_cfg_w | frontend_tlb_pmp_res_ignore )&1'h1; 
    wire frontend_tlb_pmp_res_cur_cfg_x =( frontend_tlb_pmp_io_pmp_7_cfg_x | frontend_tlb_pmp_res_ignore )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_0 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_1 = frontend_tlb_pmp_io_pmp_6_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_6_mask )==32'h0: frontend_tlb_pmp_io_pmp_6_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_6_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_1 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_6_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_6 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_7 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_8 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_9 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_10 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_11 ={ frontend_tlb_pmp_io_pmp_6_cfg_x , frontend_tlb_pmp_io_pmp_6_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_1_cfg_r =( frontend_tlb_pmp_io_pmp_6_cfg_r | frontend_tlb_pmp_res_ignore_1 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_1_cfg_w =( frontend_tlb_pmp_io_pmp_6_cfg_w | frontend_tlb_pmp_res_ignore_1 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_1_cfg_x =( frontend_tlb_pmp_io_pmp_6_cfg_x | frontend_tlb_pmp_res_ignore_1 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_1 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_2 = frontend_tlb_pmp_io_pmp_5_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_5_mask )==32'h0: frontend_tlb_pmp_io_pmp_5_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_5_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_2 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_5_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_12 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_13 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_14 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_15 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_16 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_17 ={ frontend_tlb_pmp_io_pmp_5_cfg_x , frontend_tlb_pmp_io_pmp_5_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_2_cfg_r =( frontend_tlb_pmp_io_pmp_5_cfg_r | frontend_tlb_pmp_res_ignore_2 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_2_cfg_w =( frontend_tlb_pmp_io_pmp_5_cfg_w | frontend_tlb_pmp_res_ignore_2 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_2_cfg_x =( frontend_tlb_pmp_io_pmp_5_cfg_x | frontend_tlb_pmp_res_ignore_2 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_2 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_3 = frontend_tlb_pmp_io_pmp_4_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_4_mask )==32'h0: frontend_tlb_pmp_io_pmp_4_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_4_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_3 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_4_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_18 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_19 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_20 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_21 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_22 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_23 ={ frontend_tlb_pmp_io_pmp_4_cfg_x , frontend_tlb_pmp_io_pmp_4_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_3_cfg_r =( frontend_tlb_pmp_io_pmp_4_cfg_r | frontend_tlb_pmp_res_ignore_3 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_3_cfg_w =( frontend_tlb_pmp_io_pmp_4_cfg_w | frontend_tlb_pmp_res_ignore_3 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_3_cfg_x =( frontend_tlb_pmp_io_pmp_4_cfg_x | frontend_tlb_pmp_res_ignore_3 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_3 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_4 = frontend_tlb_pmp_io_pmp_3_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_3_mask )==32'h0: frontend_tlb_pmp_io_pmp_3_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_3_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_4 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_3_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_24 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_25 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_26 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_27 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_28 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_29 ={ frontend_tlb_pmp_io_pmp_3_cfg_x , frontend_tlb_pmp_io_pmp_3_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_4_cfg_r =( frontend_tlb_pmp_io_pmp_3_cfg_r | frontend_tlb_pmp_res_ignore_4 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_4_cfg_w =( frontend_tlb_pmp_io_pmp_3_cfg_w | frontend_tlb_pmp_res_ignore_4 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_4_cfg_x =( frontend_tlb_pmp_io_pmp_3_cfg_x | frontend_tlb_pmp_res_ignore_4 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_4 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_5 = frontend_tlb_pmp_io_pmp_2_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_2_mask )==32'h0: frontend_tlb_pmp_io_pmp_2_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_2_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_5 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_2_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_30 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_31 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_32 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_33 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_34 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_35 ={ frontend_tlb_pmp_io_pmp_2_cfg_x , frontend_tlb_pmp_io_pmp_2_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_5_cfg_r =( frontend_tlb_pmp_io_pmp_2_cfg_r | frontend_tlb_pmp_res_ignore_5 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_5_cfg_w =( frontend_tlb_pmp_io_pmp_2_cfg_w | frontend_tlb_pmp_res_ignore_5 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_5_cfg_x =( frontend_tlb_pmp_io_pmp_2_cfg_x | frontend_tlb_pmp_res_ignore_5 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_5 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_6 = frontend_tlb_pmp_io_pmp_1_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_1_mask )==32'h0: frontend_tlb_pmp_io_pmp_1_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_1_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_6 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_1_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_36 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_37 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_38 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_39 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_40 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_41 ={ frontend_tlb_pmp_io_pmp_1_cfg_x , frontend_tlb_pmp_io_pmp_1_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_6_cfg_r =( frontend_tlb_pmp_io_pmp_1_cfg_r | frontend_tlb_pmp_res_ignore_6 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_6_cfg_w =( frontend_tlb_pmp_io_pmp_1_cfg_w | frontend_tlb_pmp_res_ignore_6 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_6_cfg_x =( frontend_tlb_pmp_io_pmp_1_cfg_x | frontend_tlb_pmp_res_ignore_6 )&1'h1; 
    wire[4:0] frontend_tlb_pmp__GEN_6 =5'h3<< frontend_tlb_pmp_io_size ; 
    wire frontend_tlb_pmp_res_hit_7 = frontend_tlb_pmp_io_pmp_0_cfg_a [1] ? (( frontend_tlb_pmp_io_addr ^~(~{ frontend_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3))&~ frontend_tlb_pmp_io_pmp_0_mask )==32'h0: frontend_tlb_pmp_io_pmp_0_cfg_a [0]& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_pmp0_addr ,2'h0}|32'h3)==1'h0& frontend_tlb_pmp_io_addr <~(~{ frontend_tlb_pmp_io_pmp_0_addr ,2'h0}|32'h3); 
    wire frontend_tlb_pmp_res_ignore_7 = frontend_tlb_pmp_default_0 & frontend_tlb_pmp_io_pmp_0_cfg_l ==1'h0; 
    wire[1:0] frontend_tlb_pmp_res_hi_42 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_43 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_44 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_45 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_46 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire[1:0] frontend_tlb_pmp_res_hi_47 ={ frontend_tlb_pmp_io_pmp_0_cfg_x , frontend_tlb_pmp_io_pmp_0_cfg_w }; 
    wire frontend_tlb_pmp_res_cur_7_cfg_r =( frontend_tlb_pmp_io_pmp_0_cfg_r | frontend_tlb_pmp_res_ignore_7 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_7_cfg_w =( frontend_tlb_pmp_io_pmp_0_cfg_w | frontend_tlb_pmp_res_ignore_7 )&1'h1; 
    wire frontend_tlb_pmp_res_cur_7_cfg_x =( frontend_tlb_pmp_io_pmp_0_cfg_x | frontend_tlb_pmp_res_ignore_7 )&1'h1; 
    wire frontend_tlb_pmp_res_cfg_l = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_l : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_l : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_l : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_l : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_l : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_l : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_l : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_l : frontend_tlb_pmp_pmp0_cfg_l ; 
    wire[1:0] frontend_tlb_pmp_res_cfg_res = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_res : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_res : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_res : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_res : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_res : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_res : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_res : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_res : frontend_tlb_pmp_pmp0_cfg_res ; 
    wire[1:0] frontend_tlb_pmp_res_cfg_a = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_a : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_a : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_a : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_a : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_a : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_a : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_a : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_a : frontend_tlb_pmp_pmp0_cfg_a ; 
    wire frontend_tlb_pmp_res_cfg_x = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_x : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_x : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_x : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_x : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_x : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_x : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_x : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_x : frontend_tlb_pmp_pmp0_cfg_x ; 
    wire frontend_tlb_pmp_res_cfg_w = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_w : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_w : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_w : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_w : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_w : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_w : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_w : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_w : frontend_tlb_pmp_pmp0_cfg_w ; 
    wire frontend_tlb_pmp_res_cfg_r = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_cfg_r : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_cfg_r : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_cfg_r : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_cfg_r : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_cfg_r : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_cfg_r : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_cfg_r : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_cfg_r : frontend_tlb_pmp_pmp0_cfg_r ; 
    wire[29:0] frontend_tlb_pmp_res_addr = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_addr : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_addr : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_addr : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_addr : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_addr : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_addr : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_addr : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_addr : frontend_tlb_pmp_pmp0_addr ; 
    wire[31:0] frontend_tlb_pmp_res_mask = frontend_tlb_pmp_res_hit_7  ?  frontend_tlb_pmp_res_cur_7_mask : frontend_tlb_pmp_res_hit_6  ?  frontend_tlb_pmp_res_cur_6_mask : frontend_tlb_pmp_res_hit_5  ?  frontend_tlb_pmp_res_cur_5_mask : frontend_tlb_pmp_res_hit_4  ?  frontend_tlb_pmp_res_cur_4_mask : frontend_tlb_pmp_res_hit_3  ?  frontend_tlb_pmp_res_cur_3_mask : frontend_tlb_pmp_res_hit_2  ?  frontend_tlb_pmp_res_cur_2_mask : frontend_tlb_pmp_res_hit_1  ?  frontend_tlb_pmp_res_cur_1_mask : frontend_tlb_pmp_res_hit  ?  frontend_tlb_pmp_res_cur_mask : frontend_tlb_pmp_pmp0_mask ; 
  assign  frontend_tlb_pmp_io_r = frontend_tlb_pmp_res_cfg_r ; 
  assign  frontend_tlb_pmp_io_w = frontend_tlb_pmp_res_cfg_w ; 
  assign  frontend_tlb_pmp_io_x = frontend_tlb_pmp_res_cfg_x ;
    assign frontend_tlb_pmp_clock = frontend_tlb_clock;
    assign frontend_tlb_pmp_reset = frontend_tlb_reset;
    assign frontend_tlb_pmp_io_prv = frontend_tlb__mpu_priv_1to0;
    assign frontend_tlb_pmp_io_pmp_0_cfg_l = frontend_tlb_io_ptw_pmp_0_cfg_l;
    assign frontend_tlb_pmp_io_pmp_0_cfg_res = frontend_tlb_io_ptw_pmp_0_cfg_res;
    assign frontend_tlb_pmp_io_pmp_0_cfg_a = frontend_tlb_io_ptw_pmp_0_cfg_a;
    assign frontend_tlb_pmp_io_pmp_0_cfg_x = frontend_tlb_io_ptw_pmp_0_cfg_x;
    assign frontend_tlb_pmp_io_pmp_0_cfg_w = frontend_tlb_io_ptw_pmp_0_cfg_w;
    assign frontend_tlb_pmp_io_pmp_0_cfg_r = frontend_tlb_io_ptw_pmp_0_cfg_r;
    assign frontend_tlb_pmp_io_pmp_0_addr = frontend_tlb_io_ptw_pmp_0_addr;
    assign frontend_tlb_pmp_io_pmp_0_mask = frontend_tlb_io_ptw_pmp_0_mask;
    assign frontend_tlb_pmp_io_pmp_1_cfg_l = frontend_tlb_io_ptw_pmp_1_cfg_l;
    assign frontend_tlb_pmp_io_pmp_1_cfg_res = frontend_tlb_io_ptw_pmp_1_cfg_res;
    assign frontend_tlb_pmp_io_pmp_1_cfg_a = frontend_tlb_io_ptw_pmp_1_cfg_a;
    assign frontend_tlb_pmp_io_pmp_1_cfg_x = frontend_tlb_io_ptw_pmp_1_cfg_x;
    assign frontend_tlb_pmp_io_pmp_1_cfg_w = frontend_tlb_io_ptw_pmp_1_cfg_w;
    assign frontend_tlb_pmp_io_pmp_1_cfg_r = frontend_tlb_io_ptw_pmp_1_cfg_r;
    assign frontend_tlb_pmp_io_pmp_1_addr = frontend_tlb_io_ptw_pmp_1_addr;
    assign frontend_tlb_pmp_io_pmp_1_mask = frontend_tlb_io_ptw_pmp_1_mask;
    assign frontend_tlb_pmp_io_pmp_2_cfg_l = frontend_tlb_io_ptw_pmp_2_cfg_l;
    assign frontend_tlb_pmp_io_pmp_2_cfg_res = frontend_tlb_io_ptw_pmp_2_cfg_res;
    assign frontend_tlb_pmp_io_pmp_2_cfg_a = frontend_tlb_io_ptw_pmp_2_cfg_a;
    assign frontend_tlb_pmp_io_pmp_2_cfg_x = frontend_tlb_io_ptw_pmp_2_cfg_x;
    assign frontend_tlb_pmp_io_pmp_2_cfg_w = frontend_tlb_io_ptw_pmp_2_cfg_w;
    assign frontend_tlb_pmp_io_pmp_2_cfg_r = frontend_tlb_io_ptw_pmp_2_cfg_r;
    assign frontend_tlb_pmp_io_pmp_2_addr = frontend_tlb_io_ptw_pmp_2_addr;
    assign frontend_tlb_pmp_io_pmp_2_mask = frontend_tlb_io_ptw_pmp_2_mask;
    assign frontend_tlb_pmp_io_pmp_3_cfg_l = frontend_tlb_io_ptw_pmp_3_cfg_l;
    assign frontend_tlb_pmp_io_pmp_3_cfg_res = frontend_tlb_io_ptw_pmp_3_cfg_res;
    assign frontend_tlb_pmp_io_pmp_3_cfg_a = frontend_tlb_io_ptw_pmp_3_cfg_a;
    assign frontend_tlb_pmp_io_pmp_3_cfg_x = frontend_tlb_io_ptw_pmp_3_cfg_x;
    assign frontend_tlb_pmp_io_pmp_3_cfg_w = frontend_tlb_io_ptw_pmp_3_cfg_w;
    assign frontend_tlb_pmp_io_pmp_3_cfg_r = frontend_tlb_io_ptw_pmp_3_cfg_r;
    assign frontend_tlb_pmp_io_pmp_3_addr = frontend_tlb_io_ptw_pmp_3_addr;
    assign frontend_tlb_pmp_io_pmp_3_mask = frontend_tlb_io_ptw_pmp_3_mask;
    assign frontend_tlb_pmp_io_pmp_4_cfg_l = frontend_tlb_io_ptw_pmp_4_cfg_l;
    assign frontend_tlb_pmp_io_pmp_4_cfg_res = frontend_tlb_io_ptw_pmp_4_cfg_res;
    assign frontend_tlb_pmp_io_pmp_4_cfg_a = frontend_tlb_io_ptw_pmp_4_cfg_a;
    assign frontend_tlb_pmp_io_pmp_4_cfg_x = frontend_tlb_io_ptw_pmp_4_cfg_x;
    assign frontend_tlb_pmp_io_pmp_4_cfg_w = frontend_tlb_io_ptw_pmp_4_cfg_w;
    assign frontend_tlb_pmp_io_pmp_4_cfg_r = frontend_tlb_io_ptw_pmp_4_cfg_r;
    assign frontend_tlb_pmp_io_pmp_4_addr = frontend_tlb_io_ptw_pmp_4_addr;
    assign frontend_tlb_pmp_io_pmp_4_mask = frontend_tlb_io_ptw_pmp_4_mask;
    assign frontend_tlb_pmp_io_pmp_5_cfg_l = frontend_tlb_io_ptw_pmp_5_cfg_l;
    assign frontend_tlb_pmp_io_pmp_5_cfg_res = frontend_tlb_io_ptw_pmp_5_cfg_res;
    assign frontend_tlb_pmp_io_pmp_5_cfg_a = frontend_tlb_io_ptw_pmp_5_cfg_a;
    assign frontend_tlb_pmp_io_pmp_5_cfg_x = frontend_tlb_io_ptw_pmp_5_cfg_x;
    assign frontend_tlb_pmp_io_pmp_5_cfg_w = frontend_tlb_io_ptw_pmp_5_cfg_w;
    assign frontend_tlb_pmp_io_pmp_5_cfg_r = frontend_tlb_io_ptw_pmp_5_cfg_r;
    assign frontend_tlb_pmp_io_pmp_5_addr = frontend_tlb_io_ptw_pmp_5_addr;
    assign frontend_tlb_pmp_io_pmp_5_mask = frontend_tlb_io_ptw_pmp_5_mask;
    assign frontend_tlb_pmp_io_pmp_6_cfg_l = frontend_tlb_io_ptw_pmp_6_cfg_l;
    assign frontend_tlb_pmp_io_pmp_6_cfg_res = frontend_tlb_io_ptw_pmp_6_cfg_res;
    assign frontend_tlb_pmp_io_pmp_6_cfg_a = frontend_tlb_io_ptw_pmp_6_cfg_a;
    assign frontend_tlb_pmp_io_pmp_6_cfg_x = frontend_tlb_io_ptw_pmp_6_cfg_x;
    assign frontend_tlb_pmp_io_pmp_6_cfg_w = frontend_tlb_io_ptw_pmp_6_cfg_w;
    assign frontend_tlb_pmp_io_pmp_6_cfg_r = frontend_tlb_io_ptw_pmp_6_cfg_r;
    assign frontend_tlb_pmp_io_pmp_6_addr = frontend_tlb_io_ptw_pmp_6_addr;
    assign frontend_tlb_pmp_io_pmp_6_mask = frontend_tlb_io_ptw_pmp_6_mask;
    assign frontend_tlb_pmp_io_pmp_7_cfg_l = frontend_tlb_io_ptw_pmp_7_cfg_l;
    assign frontend_tlb_pmp_io_pmp_7_cfg_res = frontend_tlb_io_ptw_pmp_7_cfg_res;
    assign frontend_tlb_pmp_io_pmp_7_cfg_a = frontend_tlb_io_ptw_pmp_7_cfg_a;
    assign frontend_tlb_pmp_io_pmp_7_cfg_x = frontend_tlb_io_ptw_pmp_7_cfg_x;
    assign frontend_tlb_pmp_io_pmp_7_cfg_w = frontend_tlb_io_ptw_pmp_7_cfg_w;
    assign frontend_tlb_pmp_io_pmp_7_cfg_r = frontend_tlb_io_ptw_pmp_7_cfg_r;
    assign frontend_tlb_pmp_io_pmp_7_addr = frontend_tlb_io_ptw_pmp_7_addr;
    assign frontend_tlb_pmp_io_pmp_7_mask = frontend_tlb_io_ptw_pmp_7_mask;
    assign frontend_tlb_pmp_io_addr = frontend_tlb__mpu_physaddr_31to0;
    assign frontend_tlb_pmp_io_size = frontend_tlb_io_req_bits_size;
    assign frontend_tlb__pmp_io_r = frontend_tlb_pmp_io_r;
    assign frontend_tlb__pmp_io_w = frontend_tlb_pmp_io_w;
    assign frontend_tlb__pmp_io_x = frontend_tlb_pmp_io_x;
     
  assign  frontend_tlb__mpu_physaddr_31to0 = frontend_tlb_mpu_physaddr [31:0]; 
  assign  frontend_tlb__mpu_priv_1to0 = frontend_tlb_mpu_priv [1:0]; 
    wire frontend_tlb__legal_address_WIRE_0 =({1'h0, frontend_tlb_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_1 =({1'h0, frontend_tlb_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_2 =({1'h0, frontend_tlb_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_3 =({1'h0, frontend_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_4 =({1'h0, frontend_tlb_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_5 =({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire frontend_tlb__legal_address_WIRE_6 =({1'h0, frontend_tlb_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0; 
    wire frontend_tlb_legal_address = frontend_tlb__legal_address_WIRE_0 | frontend_tlb__legal_address_WIRE_1 | frontend_tlb__legal_address_WIRE_2 | frontend_tlb__legal_address_WIRE_3 | frontend_tlb__legal_address_WIRE_4 | frontend_tlb__legal_address_WIRE_5 | frontend_tlb__legal_address_WIRE_6 ; 
    wire frontend_tlb__cacheable_WIRE =({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'h80000000)==35'h0|1'h0; 
    wire frontend_tlb_cacheable = frontend_tlb_legal_address & frontend_tlb__cacheable_WIRE ; 
    wire frontend_tlb_newEntry_c = frontend_tlb_cacheable ; 
    wire frontend_tlb_homogeneous =({1'h0, frontend_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0|1'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h3000}&35'h7FFFFF000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h10000}&35'h7FFFF0000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h2000000}&35'h7FFFF0000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'hC000000}&35'h7FC000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h60000000}&35'h7E0000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'h7F0000000)==35'h0; 
    wire frontend_tlb_deny_access_to_debug = frontend_tlb_mpu_priv <=3'h3&({1'h0, frontend_tlb_mpu_physaddr }&35'h7FFFFF000)==35'h0; 
    wire frontend_tlb_prot_r = frontend_tlb_legal_address & frontend_tlb_deny_access_to_debug ==1'h0& frontend_tlb__pmp_io_r ; 
    wire frontend_tlb_newEntry_pr = frontend_tlb_prot_r ; 
    wire frontend_tlb__prot_w_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire frontend_tlb_prot_w = frontend_tlb_legal_address & frontend_tlb__prot_w_WIRE & frontend_tlb_deny_access_to_debug ==1'h0& frontend_tlb__pmp_io_w ; 
    wire frontend_tlb_newEntry_pw = frontend_tlb_prot_w ; 
    wire frontend_tlb__prot_pp_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire frontend_tlb_prot_pp = frontend_tlb_legal_address & frontend_tlb__prot_pp_WIRE ; 
    wire frontend_tlb_newEntry_ppp = frontend_tlb_prot_pp ; 
    wire frontend_tlb__prot_al_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire frontend_tlb_prot_al = frontend_tlb_legal_address & frontend_tlb__prot_al_WIRE ; 
    wire frontend_tlb_newEntry_pal = frontend_tlb_prot_al ; 
    wire frontend_tlb__prot_aa_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hC8010000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0; 
    wire frontend_tlb_prot_aa = frontend_tlb_legal_address & frontend_tlb__prot_aa_WIRE ; 
    wire frontend_tlb_newEntry_paa = frontend_tlb_prot_aa ; 
    wire frontend_tlb__prot_x_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hCA000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h80000000}&35'hC0000000)==35'h0; 
    wire frontend_tlb_prot_x = frontend_tlb_legal_address & frontend_tlb__prot_x_WIRE & frontend_tlb_deny_access_to_debug ==1'h0& frontend_tlb__pmp_io_x ; 
    wire frontend_tlb_newEntry_px = frontend_tlb_prot_x ; 
    wire frontend_tlb__prot_eff_WIRE =({1'h0, frontend_tlb_mpu_physaddr }&35'hCA012000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h2000000}&35'hCA010000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h8000000}&35'hC8000000)==35'h0|({1'h0, frontend_tlb_mpu_physaddr ^34'h40000000}&35'hC0000000)==35'h0|1'h0; 
    wire frontend_tlb_prot_eff = frontend_tlb_legal_address & frontend_tlb__prot_eff_WIRE ; 
    wire frontend_tlb_newEntry_eff = frontend_tlb_prot_eff ; 
    wire[20:0] frontend_tlb__GEN = frontend_tlb_sectored_entries_0_0_tag_vpn ^ frontend_tlb_vpn ; 
    wire frontend_tlb_sector_hits_0 =( frontend_tlb_sectored_entries_0_0_valid_0 | frontend_tlb_sectored_entries_0_0_valid_1 | frontend_tlb_sectored_entries_0_0_valid_2 | frontend_tlb_sectored_entries_0_0_valid_3 )& frontend_tlb__GEN [20:2]==19'h0& frontend_tlb_sectored_entries_0_0_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_superpage_hits_0 = frontend_tlb_superpage_entries_0_valid_0 &( frontend_tlb_superpage_entries_0_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_0_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_superpage_hits_1 = frontend_tlb_superpage_entries_1_valid_0 &( frontend_tlb_superpage_entries_1_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_1_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_superpage_hits_2 = frontend_tlb_superpage_entries_2_valid_0 &( frontend_tlb_superpage_entries_2_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_2_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_superpage_hits_3 = frontend_tlb_superpage_entries_3_valid_0 &( frontend_tlb_superpage_entries_3_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_3_tag_v == frontend_tlb_priv_v ; 
    wire[1:0] frontend_tlb_hitsVec_idx = frontend_tlb_vpn [1:0]; 
    wire[20:0] frontend_tlb__GEN_0 = frontend_tlb_sectored_entries_0_0_tag_vpn ^ frontend_tlb_vpn ; 
    reg frontend_tlb_casez_tmp ; 
  always @(*)
         begin 
             casez ( frontend_tlb_hitsVec_idx )
              2 'b00: 
                  frontend_tlb_casez_tmp  = frontend_tlb_sectored_entries_0_0_valid_0 ;
              2 'b01: 
                  frontend_tlb_casez_tmp  = frontend_tlb_sectored_entries_0_0_valid_1 ;
              2 'b10: 
                  frontend_tlb_casez_tmp  = frontend_tlb_sectored_entries_0_0_valid_2 ;
              default : 
                  frontend_tlb_casez_tmp  = frontend_tlb_sectored_entries_0_0_valid_3 ;endcase
         end
    wire frontend_tlb_hitsVec_0 = frontend_tlb_vm_enabled & frontend_tlb_casez_tmp & frontend_tlb__GEN_0 [20:2]==19'h0& frontend_tlb_sectored_entries_0_0_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_hitsVec_1 = frontend_tlb_vm_enabled & frontend_tlb_superpage_entries_0_valid_0 &( frontend_tlb_superpage_entries_0_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_0_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_hitsVec_2 = frontend_tlb_vm_enabled & frontend_tlb_superpage_entries_1_valid_0 &( frontend_tlb_superpage_entries_1_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_1_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_hitsVec_3 = frontend_tlb_vm_enabled & frontend_tlb_superpage_entries_2_valid_0 &( frontend_tlb_superpage_entries_2_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_2_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_hitsVec_4 = frontend_tlb_vm_enabled & frontend_tlb_superpage_entries_3_valid_0 &( frontend_tlb_superpage_entries_3_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_superpage_entries_3_tag_v == frontend_tlb_priv_v ; 
    wire frontend_tlb_hitsVec_5 = frontend_tlb_vm_enabled & frontend_tlb_special_entry_valid_0 &( frontend_tlb_special_entry_tag_vpn ^ frontend_tlb_vpn )==21'h0& frontend_tlb_special_entry_tag_v == frontend_tlb_priv_v ; 
    wire[1:0] frontend_tlb_real_hits_lo_hi ={ frontend_tlb_hitsVec_2 , frontend_tlb_hitsVec_1 }; 
    wire[2:0] frontend_tlb_real_hits_lo ={ frontend_tlb_real_hits_lo_hi , frontend_tlb_hitsVec_0 }; 
    wire[1:0] frontend_tlb_real_hits_hi_hi ={ frontend_tlb_hitsVec_5 , frontend_tlb_hitsVec_4 }; 
    wire[2:0] frontend_tlb_real_hits_hi ={ frontend_tlb_real_hits_hi_hi , frontend_tlb_hitsVec_3 }; 
    wire[5:0] frontend_tlb_real_hits ={ frontend_tlb_real_hits_hi , frontend_tlb_real_hits_lo }; 
    wire[6:0] frontend_tlb_hits ={ frontend_tlb_vm_enabled ==1'h0, frontend_tlb_real_hits }; 
    wire frontend_tlb_refill_v = frontend_tlb_r_vstage1_en | frontend_tlb_r_stage2_en ; 
    wire[19:0] frontend_tlb_newEntry_ppn = frontend_tlb_io_ptw_resp_bits_pte_ppn [19:0]; 
    wire frontend_tlb_newEntry_g = frontend_tlb_io_ptw_resp_bits_pte_g & frontend_tlb_io_ptw_resp_bits_pte_v ; 
    wire frontend_tlb_newEntry_ae_stage2 = frontend_tlb_io_ptw_resp_bits_ae_final & frontend_tlb_io_ptw_resp_bits_gpa_is_pte & frontend_tlb_r_stage2_en ; 
    wire frontend_tlb_newEntry_sr = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x & frontend_tlb_io_ptw_resp_bits_pte_w ==1'h0)& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_r ; 
    wire frontend_tlb_newEntry_sw = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x & frontend_tlb_io_ptw_resp_bits_pte_w ==1'h0)& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_w & frontend_tlb_io_ptw_resp_bits_pte_d ; 
    wire frontend_tlb_newEntry_sx = frontend_tlb_io_ptw_resp_bits_pte_v &( frontend_tlb_io_ptw_resp_bits_pte_r | frontend_tlb_io_ptw_resp_bits_pte_x & frontend_tlb_io_ptw_resp_bits_pte_w ==1'h0)& frontend_tlb_io_ptw_resp_bits_pte_a & frontend_tlb_io_ptw_resp_bits_pte_x ; 
    wire frontend_tlb__GEN_1 = frontend_tlb_io_ptw_resp_bits_homogeneous ==1'h0&1'h1; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_lo_hi ={ frontend_tlb_special_entry_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_special_entry_data_0_lo_lo ={ frontend_tlb_special_entry_data_0_lo_lo_hi , frontend_tlb_special_entry_data_0_lo_lo_lo }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_hi_lo ={ frontend_tlb_special_entry_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_special_entry_data_0_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_special_entry_data_0_lo_hi_hi ={ frontend_tlb_special_entry_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_special_entry_data_0_lo_hi ={ frontend_tlb_special_entry_data_0_lo_hi_hi , frontend_tlb_special_entry_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_special_entry_data_0_lo ={ frontend_tlb_special_entry_data_0_lo_hi , frontend_tlb_special_entry_data_0_lo_lo }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_lo_lo ={ frontend_tlb_special_entry_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_lo_hi ={ frontend_tlb_special_entry_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_special_entry_data_0_hi_lo ={ frontend_tlb_special_entry_data_0_hi_lo_hi , frontend_tlb_special_entry_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb_special_entry_data_0_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_special_entry_data_0_hi_hi_lo ={ frontend_tlb_special_entry_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_special_entry_data_0_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_special_entry_data_0_hi_hi_hi ={ frontend_tlb_special_entry_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_special_entry_data_0_hi_hi ={ frontend_tlb_special_entry_data_0_hi_hi_hi , frontend_tlb_special_entry_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_special_entry_data_0_hi ={ frontend_tlb_special_entry_data_0_hi_hi , frontend_tlb_special_entry_data_0_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_2 ={ frontend_tlb_special_entry_data_0_hi , frontend_tlb_special_entry_data_0_lo }; 
    wire frontend_tlb__GEN_3 = frontend_tlb_do_refill &~ frontend_tlb__GEN_1 ; 
    wire frontend_tlb__GEN_4 = frontend_tlb_io_ptw_resp_bits_level <2'h2; 
    wire frontend_tlb__GEN_5 = frontend_tlb__GEN_3 & frontend_tlb__GEN_4 ; 
    wire frontend_tlb__GEN_6 = frontend_tlb_r_superpage_repl_addr ==2'h0; 
    wire[1:0] frontend_tlb__GEN_7 ={1'h0, frontend_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_0_data_0_lo_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_lo_hi , frontend_tlb_superpage_entries_0_data_0_lo_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_0_data_0_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_lo_hi_hi , frontend_tlb_superpage_entries_0_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_0_data_0_lo ={ frontend_tlb_superpage_entries_0_data_0_lo_hi , frontend_tlb_superpage_entries_0_data_0_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_0_data_0_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_lo_hi , frontend_tlb_superpage_entries_0_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_superpage_entries_0_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_0_data_0_hi_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi_hi , frontend_tlb_superpage_entries_0_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_0_data_0_hi ={ frontend_tlb_superpage_entries_0_data_0_hi_hi , frontend_tlb_superpage_entries_0_data_0_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_8 ={ frontend_tlb_superpage_entries_0_data_0_hi , frontend_tlb_superpage_entries_0_data_0_lo }; 
    wire frontend_tlb__GEN_9 = frontend_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire frontend_tlb__GEN_10 = frontend_tlb_r_superpage_repl_addr ==2'h1; 
    wire[1:0] frontend_tlb__GEN_11 ={1'h0, frontend_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_1_data_0_lo_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_lo_hi , frontend_tlb_superpage_entries_1_data_0_lo_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_1_data_0_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_lo_hi_hi , frontend_tlb_superpage_entries_1_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_1_data_0_lo ={ frontend_tlb_superpage_entries_1_data_0_lo_hi , frontend_tlb_superpage_entries_1_data_0_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_1_data_0_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_lo_hi , frontend_tlb_superpage_entries_1_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_superpage_entries_1_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_1_data_0_hi_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi_hi , frontend_tlb_superpage_entries_1_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_1_data_0_hi ={ frontend_tlb_superpage_entries_1_data_0_hi_hi , frontend_tlb_superpage_entries_1_data_0_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_12 ={ frontend_tlb_superpage_entries_1_data_0_hi , frontend_tlb_superpage_entries_1_data_0_lo }; 
    wire frontend_tlb__GEN_13 = frontend_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire frontend_tlb__GEN_14 = frontend_tlb_r_superpage_repl_addr ==2'h2; 
    wire[1:0] frontend_tlb__GEN_15 ={1'h0, frontend_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_2_data_0_lo_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_lo_hi , frontend_tlb_superpage_entries_2_data_0_lo_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_2_data_0_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_lo_hi_hi , frontend_tlb_superpage_entries_2_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_2_data_0_lo ={ frontend_tlb_superpage_entries_2_data_0_lo_hi , frontend_tlb_superpage_entries_2_data_0_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_2_data_0_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_lo_hi , frontend_tlb_superpage_entries_2_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_superpage_entries_2_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_2_data_0_hi_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi_hi , frontend_tlb_superpage_entries_2_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_2_data_0_hi ={ frontend_tlb_superpage_entries_2_data_0_hi_hi , frontend_tlb_superpage_entries_2_data_0_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_16 ={ frontend_tlb_superpage_entries_2_data_0_hi , frontend_tlb_superpage_entries_2_data_0_lo }; 
    wire frontend_tlb__GEN_17 = frontend_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire frontend_tlb__GEN_18 =& frontend_tlb_r_superpage_repl_addr ; 
    wire[1:0] frontend_tlb__GEN_19 ={1'h0, frontend_tlb_io_ptw_resp_bits_level [0]}; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_superpage_entries_3_data_0_lo_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_lo_hi , frontend_tlb_superpage_entries_3_data_0_lo_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_lo_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_superpage_entries_3_data_0_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_lo_hi_hi , frontend_tlb_superpage_entries_3_data_0_lo_hi_lo }; 
    wire[10:0] frontend_tlb_superpage_entries_3_data_0_lo ={ frontend_tlb_superpage_entries_3_data_0_lo_hi , frontend_tlb_superpage_entries_3_data_0_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_lo_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_superpage_entries_3_data_0_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_lo_hi , frontend_tlb_superpage_entries_3_data_0_hi_lo_lo }; 
    wire[1:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_lo ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_superpage_entries_3_data_0_hi_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_superpage_entries_3_data_0_hi_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi_hi , frontend_tlb_superpage_entries_3_data_0_hi_hi_lo }; 
    wire[30:0] frontend_tlb_superpage_entries_3_data_0_hi ={ frontend_tlb_superpage_entries_3_data_0_hi_hi , frontend_tlb_superpage_entries_3_data_0_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_20 ={ frontend_tlb_superpage_entries_3_data_0_hi , frontend_tlb_superpage_entries_3_data_0_lo }; 
    wire frontend_tlb__GEN_21 = frontend_tlb_invalidate_refill  ? 1'h0:1'h1; 
    wire frontend_tlb__GEN_22 = frontend_tlb__GEN_3 &~ frontend_tlb__GEN_4 ; 
    wire frontend_tlb__GEN_23 = frontend_tlb_r_sectored_hit_valid ==1'h0; 
    wire[1:0] frontend_tlb_idx = frontend_tlb_r_refill_tag [1:0]; 
    wire frontend_tlb__GEN_24 = frontend_tlb_idx ==2'h0; 
    wire frontend_tlb__GEN_25 = frontend_tlb_idx ==2'h1; 
    wire frontend_tlb__GEN_26 = frontend_tlb_idx ==2'h2; 
    wire frontend_tlb__GEN_27 =& frontend_tlb_idx ; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_lo ={ frontend_tlb_newEntry_c , frontend_tlb_newEntry_fragmented_superpage }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_hi_hi ={ frontend_tlb_newEntry_pal , frontend_tlb_newEntry_paa }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_lo_hi_hi , frontend_tlb_newEntry_eff }; 
    wire[4:0] frontend_tlb_sectored_entries_0_0_data_lo_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_lo_hi , frontend_tlb_sectored_entries_0_0_data_lo_lo_lo }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_lo_hi ={ frontend_tlb_newEntry_px , frontend_tlb_newEntry_pr }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_lo_hi , frontend_tlb_newEntry_ppp }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_hi_hi ={ frontend_tlb_newEntry_hx , frontend_tlb_newEntry_hr }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_lo_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_hi_hi , frontend_tlb_newEntry_pw }; 
    wire[5:0] frontend_tlb_sectored_entries_0_0_data_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_lo_hi_hi , frontend_tlb_sectored_entries_0_0_data_lo_hi_lo }; 
    wire[10:0] frontend_tlb_sectored_entries_0_0_data_lo ={ frontend_tlb_sectored_entries_0_0_data_lo_hi , frontend_tlb_sectored_entries_0_0_data_lo_lo }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_lo_hi ={ frontend_tlb_newEntry_sx , frontend_tlb_newEntry_sr }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_lo_hi , frontend_tlb_newEntry_hw }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_hi_hi ={ frontend_tlb_newEntry_pf , frontend_tlb_newEntry_gf }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_lo_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_hi_hi , frontend_tlb_newEntry_sw }; 
    wire[5:0] frontend_tlb_sectored_entries_0_0_data_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_lo_hi , frontend_tlb_sectored_entries_0_0_data_hi_lo_lo }; 
    wire[1:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_lo_hi ={ frontend_tlb_newEntry_ae_ptw , frontend_tlb_newEntry_ae_final }; 
    wire[2:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_lo ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_lo_hi , frontend_tlb_newEntry_ae_stage2 }; 
    wire[20:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_hi_hi ={ frontend_tlb_newEntry_ppn , frontend_tlb_newEntry_u }; 
    wire[21:0] frontend_tlb_sectored_entries_0_0_data_hi_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_hi_hi , frontend_tlb_newEntry_g }; 
    wire[24:0] frontend_tlb_sectored_entries_0_0_data_hi_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi_hi , frontend_tlb_sectored_entries_0_0_data_hi_hi_lo }; 
    wire[30:0] frontend_tlb_sectored_entries_0_0_data_hi ={ frontend_tlb_sectored_entries_0_0_data_hi_hi , frontend_tlb_sectored_entries_0_0_data_hi_lo }; 
    wire[41:0] frontend_tlb__GEN_28 ={ frontend_tlb_sectored_entries_0_0_data_hi , frontend_tlb_sectored_entries_0_0_data_lo }; 
    wire frontend_tlb__GEN_29 = frontend_tlb_idx ==2'h0; 
    wire frontend_tlb__GEN_30 = frontend_tlb_idx ==2'h1; 
    wire frontend_tlb__GEN_31 = frontend_tlb_idx ==2'h2; 
    wire frontend_tlb__GEN_32 =& frontend_tlb_idx ; reg[41:0] frontend_tlb_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( frontend_tlb_vpn [1:0])
              2 'b00: 
                  frontend_tlb_casez_tmp_0  = frontend_tlb_sectored_entries_0_0_data_0 ;
              2 'b01: 
                  frontend_tlb_casez_tmp_0  = frontend_tlb_sectored_entries_0_0_data_1 ;
              2 'b10: 
                  frontend_tlb_casez_tmp_0  = frontend_tlb_sectored_entries_0_0_data_2 ;
              default : 
                  frontend_tlb_casez_tmp_0  = frontend_tlb_sectored_entries_0_0_data_3 ;endcase
         end
    wire[41:0] frontend_tlb__entries_WIRE_1 = frontend_tlb_casez_tmp_0 ; 
    wire frontend_tlb__entries_WIRE_fragmented_superpage = frontend_tlb__entries_WIRE_1 [0]; 
    wire frontend_tlb__entries_WIRE_c = frontend_tlb__entries_WIRE_1 [1]; 
    wire frontend_tlb__entries_WIRE_eff = frontend_tlb__entries_WIRE_1 [2]; 
    wire frontend_tlb__entries_WIRE_paa = frontend_tlb__entries_WIRE_1 [3]; 
    wire frontend_tlb__entries_WIRE_pal = frontend_tlb__entries_WIRE_1 [4]; 
    wire frontend_tlb__entries_WIRE_ppp = frontend_tlb__entries_WIRE_1 [5]; 
    wire frontend_tlb__entries_WIRE_pr = frontend_tlb__entries_WIRE_1 [6]; 
    wire frontend_tlb__entries_WIRE_px = frontend_tlb__entries_WIRE_1 [7]; 
    wire frontend_tlb__entries_WIRE_pw = frontend_tlb__entries_WIRE_1 [8]; 
    wire frontend_tlb__entries_WIRE_hr = frontend_tlb__entries_WIRE_1 [9]; 
    wire frontend_tlb__entries_WIRE_hx = frontend_tlb__entries_WIRE_1 [10]; 
    wire frontend_tlb__entries_WIRE_hw = frontend_tlb__entries_WIRE_1 [11]; 
    wire frontend_tlb__entries_WIRE_sr = frontend_tlb__entries_WIRE_1 [12]; 
    wire frontend_tlb__entries_WIRE_sx = frontend_tlb__entries_WIRE_1 [13]; 
    wire frontend_tlb__entries_WIRE_sw = frontend_tlb__entries_WIRE_1 [14]; 
    wire frontend_tlb__entries_WIRE_gf = frontend_tlb__entries_WIRE_1 [15]; 
    wire frontend_tlb__entries_WIRE_pf = frontend_tlb__entries_WIRE_1 [16]; 
    wire frontend_tlb__entries_WIRE_ae_stage2 = frontend_tlb__entries_WIRE_1 [17]; 
    wire frontend_tlb__entries_WIRE_ae_final = frontend_tlb__entries_WIRE_1 [18]; 
    wire frontend_tlb__entries_WIRE_ae_ptw = frontend_tlb__entries_WIRE_1 [19]; 
    wire frontend_tlb__entries_WIRE_g = frontend_tlb__entries_WIRE_1 [20]; 
    wire frontend_tlb__entries_WIRE_u = frontend_tlb__entries_WIRE_1 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_ppn = frontend_tlb__entries_WIRE_1 [41:22];  
    
    assign  frontend_tlb_entries_barrier_io_y_ppn = frontend_tlb_entries_barrier_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_io_y_u = frontend_tlb_entries_barrier_io_x_u ; 
  assign  frontend_tlb_entries_barrier_io_y_g = frontend_tlb_entries_barrier_io_x_g ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_ptw = frontend_tlb_entries_barrier_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_final = frontend_tlb_entries_barrier_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_io_y_ae_stage2 = frontend_tlb_entries_barrier_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_io_y_pf = frontend_tlb_entries_barrier_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_io_y_gf = frontend_tlb_entries_barrier_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_io_y_sw = frontend_tlb_entries_barrier_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_io_y_sx = frontend_tlb_entries_barrier_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_io_y_sr = frontend_tlb_entries_barrier_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_io_y_hw = frontend_tlb_entries_barrier_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_io_y_hx = frontend_tlb_entries_barrier_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_io_y_hr = frontend_tlb_entries_barrier_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_io_y_pw = frontend_tlb_entries_barrier_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_io_y_px = frontend_tlb_entries_barrier_io_x_px ; 
  assign  frontend_tlb_entries_barrier_io_y_pr = frontend_tlb_entries_barrier_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_io_y_ppp = frontend_tlb_entries_barrier_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_io_y_pal = frontend_tlb_entries_barrier_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_io_y_paa = frontend_tlb_entries_barrier_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_io_y_eff = frontend_tlb_entries_barrier_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_io_y_c = frontend_tlb_entries_barrier_io_x_c ; 
  assign  frontend_tlb_entries_barrier_io_y_fragmented_superpage = frontend_tlb_entries_barrier_io_x_fragmented_superpage ;
     
    wire frontend_tlb__entries_WIRE_2_fragmented_superpage = frontend_tlb__entries_WIRE_3 [0]; 
    wire frontend_tlb__entries_WIRE_2_c = frontend_tlb__entries_WIRE_3 [1]; 
    wire frontend_tlb__entries_WIRE_2_eff = frontend_tlb__entries_WIRE_3 [2]; 
    wire frontend_tlb__entries_WIRE_2_paa = frontend_tlb__entries_WIRE_3 [3]; 
    wire frontend_tlb__entries_WIRE_2_pal = frontend_tlb__entries_WIRE_3 [4]; 
    wire frontend_tlb__entries_WIRE_2_ppp = frontend_tlb__entries_WIRE_3 [5]; 
    wire frontend_tlb__entries_WIRE_2_pr = frontend_tlb__entries_WIRE_3 [6]; 
    wire frontend_tlb__entries_WIRE_2_px = frontend_tlb__entries_WIRE_3 [7]; 
    wire frontend_tlb__entries_WIRE_2_pw = frontend_tlb__entries_WIRE_3 [8]; 
    wire frontend_tlb__entries_WIRE_2_hr = frontend_tlb__entries_WIRE_3 [9]; 
    wire frontend_tlb__entries_WIRE_2_hx = frontend_tlb__entries_WIRE_3 [10]; 
    wire frontend_tlb__entries_WIRE_2_hw = frontend_tlb__entries_WIRE_3 [11]; 
    wire frontend_tlb__entries_WIRE_2_sr = frontend_tlb__entries_WIRE_3 [12]; 
    wire frontend_tlb__entries_WIRE_2_sx = frontend_tlb__entries_WIRE_3 [13]; 
    wire frontend_tlb__entries_WIRE_2_sw = frontend_tlb__entries_WIRE_3 [14]; 
    wire frontend_tlb__entries_WIRE_2_gf = frontend_tlb__entries_WIRE_3 [15]; 
    wire frontend_tlb__entries_WIRE_2_pf = frontend_tlb__entries_WIRE_3 [16]; 
    wire frontend_tlb__entries_WIRE_2_ae_stage2 = frontend_tlb__entries_WIRE_3 [17]; 
    wire frontend_tlb__entries_WIRE_2_ae_final = frontend_tlb__entries_WIRE_3 [18]; 
    wire frontend_tlb__entries_WIRE_2_ae_ptw = frontend_tlb__entries_WIRE_3 [19]; 
    wire frontend_tlb__entries_WIRE_2_g = frontend_tlb__entries_WIRE_3 [20]; 
    wire frontend_tlb__entries_WIRE_2_u = frontend_tlb__entries_WIRE_3 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_2_ppn = frontend_tlb__entries_WIRE_3 [41:22];  
    
    assign  frontend_tlb_entries_barrier_1_io_y_ppn = frontend_tlb_entries_barrier_1_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_1_io_y_u = frontend_tlb_entries_barrier_1_io_x_u ; 
  assign  frontend_tlb_entries_barrier_1_io_y_g = frontend_tlb_entries_barrier_1_io_x_g ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_ptw = frontend_tlb_entries_barrier_1_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_final = frontend_tlb_entries_barrier_1_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ae_stage2 = frontend_tlb_entries_barrier_1_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pf = frontend_tlb_entries_barrier_1_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_1_io_y_gf = frontend_tlb_entries_barrier_1_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sw = frontend_tlb_entries_barrier_1_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sx = frontend_tlb_entries_barrier_1_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_1_io_y_sr = frontend_tlb_entries_barrier_1_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hw = frontend_tlb_entries_barrier_1_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hx = frontend_tlb_entries_barrier_1_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_1_io_y_hr = frontend_tlb_entries_barrier_1_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pw = frontend_tlb_entries_barrier_1_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_1_io_y_px = frontend_tlb_entries_barrier_1_io_x_px ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pr = frontend_tlb_entries_barrier_1_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_1_io_y_ppp = frontend_tlb_entries_barrier_1_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_1_io_y_pal = frontend_tlb_entries_barrier_1_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_1_io_y_paa = frontend_tlb_entries_barrier_1_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_1_io_y_eff = frontend_tlb_entries_barrier_1_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_1_io_y_c = frontend_tlb_entries_barrier_1_io_x_c ; 
  assign  frontend_tlb_entries_barrier_1_io_y_fragmented_superpage = frontend_tlb_entries_barrier_1_io_x_fragmented_superpage ;
     
    wire frontend_tlb__entries_WIRE_4_fragmented_superpage = frontend_tlb__entries_WIRE_5 [0]; 
    wire frontend_tlb__entries_WIRE_4_c = frontend_tlb__entries_WIRE_5 [1]; 
    wire frontend_tlb__entries_WIRE_4_eff = frontend_tlb__entries_WIRE_5 [2]; 
    wire frontend_tlb__entries_WIRE_4_paa = frontend_tlb__entries_WIRE_5 [3]; 
    wire frontend_tlb__entries_WIRE_4_pal = frontend_tlb__entries_WIRE_5 [4]; 
    wire frontend_tlb__entries_WIRE_4_ppp = frontend_tlb__entries_WIRE_5 [5]; 
    wire frontend_tlb__entries_WIRE_4_pr = frontend_tlb__entries_WIRE_5 [6]; 
    wire frontend_tlb__entries_WIRE_4_px = frontend_tlb__entries_WIRE_5 [7]; 
    wire frontend_tlb__entries_WIRE_4_pw = frontend_tlb__entries_WIRE_5 [8]; 
    wire frontend_tlb__entries_WIRE_4_hr = frontend_tlb__entries_WIRE_5 [9]; 
    wire frontend_tlb__entries_WIRE_4_hx = frontend_tlb__entries_WIRE_5 [10]; 
    wire frontend_tlb__entries_WIRE_4_hw = frontend_tlb__entries_WIRE_5 [11]; 
    wire frontend_tlb__entries_WIRE_4_sr = frontend_tlb__entries_WIRE_5 [12]; 
    wire frontend_tlb__entries_WIRE_4_sx = frontend_tlb__entries_WIRE_5 [13]; 
    wire frontend_tlb__entries_WIRE_4_sw = frontend_tlb__entries_WIRE_5 [14]; 
    wire frontend_tlb__entries_WIRE_4_gf = frontend_tlb__entries_WIRE_5 [15]; 
    wire frontend_tlb__entries_WIRE_4_pf = frontend_tlb__entries_WIRE_5 [16]; 
    wire frontend_tlb__entries_WIRE_4_ae_stage2 = frontend_tlb__entries_WIRE_5 [17]; 
    wire frontend_tlb__entries_WIRE_4_ae_final = frontend_tlb__entries_WIRE_5 [18]; 
    wire frontend_tlb__entries_WIRE_4_ae_ptw = frontend_tlb__entries_WIRE_5 [19]; 
    wire frontend_tlb__entries_WIRE_4_g = frontend_tlb__entries_WIRE_5 [20]; 
    wire frontend_tlb__entries_WIRE_4_u = frontend_tlb__entries_WIRE_5 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_4_ppn = frontend_tlb__entries_WIRE_5 [41:22];  
    
    assign  frontend_tlb_entries_barrier_2_io_y_ppn = frontend_tlb_entries_barrier_2_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_2_io_y_u = frontend_tlb_entries_barrier_2_io_x_u ; 
  assign  frontend_tlb_entries_barrier_2_io_y_g = frontend_tlb_entries_barrier_2_io_x_g ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_ptw = frontend_tlb_entries_barrier_2_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_final = frontend_tlb_entries_barrier_2_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ae_stage2 = frontend_tlb_entries_barrier_2_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pf = frontend_tlb_entries_barrier_2_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_2_io_y_gf = frontend_tlb_entries_barrier_2_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sw = frontend_tlb_entries_barrier_2_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sx = frontend_tlb_entries_barrier_2_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_2_io_y_sr = frontend_tlb_entries_barrier_2_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hw = frontend_tlb_entries_barrier_2_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hx = frontend_tlb_entries_barrier_2_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_2_io_y_hr = frontend_tlb_entries_barrier_2_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pw = frontend_tlb_entries_barrier_2_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_2_io_y_px = frontend_tlb_entries_barrier_2_io_x_px ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pr = frontend_tlb_entries_barrier_2_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_2_io_y_ppp = frontend_tlb_entries_barrier_2_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_2_io_y_pal = frontend_tlb_entries_barrier_2_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_2_io_y_paa = frontend_tlb_entries_barrier_2_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_2_io_y_eff = frontend_tlb_entries_barrier_2_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_2_io_y_c = frontend_tlb_entries_barrier_2_io_x_c ; 
  assign  frontend_tlb_entries_barrier_2_io_y_fragmented_superpage = frontend_tlb_entries_barrier_2_io_x_fragmented_superpage ;
     
    wire frontend_tlb__entries_WIRE_6_fragmented_superpage = frontend_tlb__entries_WIRE_7 [0]; 
    wire frontend_tlb__entries_WIRE_6_c = frontend_tlb__entries_WIRE_7 [1]; 
    wire frontend_tlb__entries_WIRE_6_eff = frontend_tlb__entries_WIRE_7 [2]; 
    wire frontend_tlb__entries_WIRE_6_paa = frontend_tlb__entries_WIRE_7 [3]; 
    wire frontend_tlb__entries_WIRE_6_pal = frontend_tlb__entries_WIRE_7 [4]; 
    wire frontend_tlb__entries_WIRE_6_ppp = frontend_tlb__entries_WIRE_7 [5]; 
    wire frontend_tlb__entries_WIRE_6_pr = frontend_tlb__entries_WIRE_7 [6]; 
    wire frontend_tlb__entries_WIRE_6_px = frontend_tlb__entries_WIRE_7 [7]; 
    wire frontend_tlb__entries_WIRE_6_pw = frontend_tlb__entries_WIRE_7 [8]; 
    wire frontend_tlb__entries_WIRE_6_hr = frontend_tlb__entries_WIRE_7 [9]; 
    wire frontend_tlb__entries_WIRE_6_hx = frontend_tlb__entries_WIRE_7 [10]; 
    wire frontend_tlb__entries_WIRE_6_hw = frontend_tlb__entries_WIRE_7 [11]; 
    wire frontend_tlb__entries_WIRE_6_sr = frontend_tlb__entries_WIRE_7 [12]; 
    wire frontend_tlb__entries_WIRE_6_sx = frontend_tlb__entries_WIRE_7 [13]; 
    wire frontend_tlb__entries_WIRE_6_sw = frontend_tlb__entries_WIRE_7 [14]; 
    wire frontend_tlb__entries_WIRE_6_gf = frontend_tlb__entries_WIRE_7 [15]; 
    wire frontend_tlb__entries_WIRE_6_pf = frontend_tlb__entries_WIRE_7 [16]; 
    wire frontend_tlb__entries_WIRE_6_ae_stage2 = frontend_tlb__entries_WIRE_7 [17]; 
    wire frontend_tlb__entries_WIRE_6_ae_final = frontend_tlb__entries_WIRE_7 [18]; 
    wire frontend_tlb__entries_WIRE_6_ae_ptw = frontend_tlb__entries_WIRE_7 [19]; 
    wire frontend_tlb__entries_WIRE_6_g = frontend_tlb__entries_WIRE_7 [20]; 
    wire frontend_tlb__entries_WIRE_6_u = frontend_tlb__entries_WIRE_7 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_6_ppn = frontend_tlb__entries_WIRE_7 [41:22];  
    
    assign  frontend_tlb_entries_barrier_3_io_y_ppn = frontend_tlb_entries_barrier_3_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_3_io_y_u = frontend_tlb_entries_barrier_3_io_x_u ; 
  assign  frontend_tlb_entries_barrier_3_io_y_g = frontend_tlb_entries_barrier_3_io_x_g ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_ptw = frontend_tlb_entries_barrier_3_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_final = frontend_tlb_entries_barrier_3_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ae_stage2 = frontend_tlb_entries_barrier_3_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pf = frontend_tlb_entries_barrier_3_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_3_io_y_gf = frontend_tlb_entries_barrier_3_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sw = frontend_tlb_entries_barrier_3_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sx = frontend_tlb_entries_barrier_3_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_3_io_y_sr = frontend_tlb_entries_barrier_3_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hw = frontend_tlb_entries_barrier_3_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hx = frontend_tlb_entries_barrier_3_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_3_io_y_hr = frontend_tlb_entries_barrier_3_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pw = frontend_tlb_entries_barrier_3_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_3_io_y_px = frontend_tlb_entries_barrier_3_io_x_px ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pr = frontend_tlb_entries_barrier_3_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_3_io_y_ppp = frontend_tlb_entries_barrier_3_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_3_io_y_pal = frontend_tlb_entries_barrier_3_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_3_io_y_paa = frontend_tlb_entries_barrier_3_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_3_io_y_eff = frontend_tlb_entries_barrier_3_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_3_io_y_c = frontend_tlb_entries_barrier_3_io_x_c ; 
  assign  frontend_tlb_entries_barrier_3_io_y_fragmented_superpage = frontend_tlb_entries_barrier_3_io_x_fragmented_superpage ;
     
    wire frontend_tlb__entries_WIRE_8_fragmented_superpage = frontend_tlb__entries_WIRE_9 [0]; 
    wire frontend_tlb__entries_WIRE_8_c = frontend_tlb__entries_WIRE_9 [1]; 
    wire frontend_tlb__entries_WIRE_8_eff = frontend_tlb__entries_WIRE_9 [2]; 
    wire frontend_tlb__entries_WIRE_8_paa = frontend_tlb__entries_WIRE_9 [3]; 
    wire frontend_tlb__entries_WIRE_8_pal = frontend_tlb__entries_WIRE_9 [4]; 
    wire frontend_tlb__entries_WIRE_8_ppp = frontend_tlb__entries_WIRE_9 [5]; 
    wire frontend_tlb__entries_WIRE_8_pr = frontend_tlb__entries_WIRE_9 [6]; 
    wire frontend_tlb__entries_WIRE_8_px = frontend_tlb__entries_WIRE_9 [7]; 
    wire frontend_tlb__entries_WIRE_8_pw = frontend_tlb__entries_WIRE_9 [8]; 
    wire frontend_tlb__entries_WIRE_8_hr = frontend_tlb__entries_WIRE_9 [9]; 
    wire frontend_tlb__entries_WIRE_8_hx = frontend_tlb__entries_WIRE_9 [10]; 
    wire frontend_tlb__entries_WIRE_8_hw = frontend_tlb__entries_WIRE_9 [11]; 
    wire frontend_tlb__entries_WIRE_8_sr = frontend_tlb__entries_WIRE_9 [12]; 
    wire frontend_tlb__entries_WIRE_8_sx = frontend_tlb__entries_WIRE_9 [13]; 
    wire frontend_tlb__entries_WIRE_8_sw = frontend_tlb__entries_WIRE_9 [14]; 
    wire frontend_tlb__entries_WIRE_8_gf = frontend_tlb__entries_WIRE_9 [15]; 
    wire frontend_tlb__entries_WIRE_8_pf = frontend_tlb__entries_WIRE_9 [16]; 
    wire frontend_tlb__entries_WIRE_8_ae_stage2 = frontend_tlb__entries_WIRE_9 [17]; 
    wire frontend_tlb__entries_WIRE_8_ae_final = frontend_tlb__entries_WIRE_9 [18]; 
    wire frontend_tlb__entries_WIRE_8_ae_ptw = frontend_tlb__entries_WIRE_9 [19]; 
    wire frontend_tlb__entries_WIRE_8_g = frontend_tlb__entries_WIRE_9 [20]; 
    wire frontend_tlb__entries_WIRE_8_u = frontend_tlb__entries_WIRE_9 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_8_ppn = frontend_tlb__entries_WIRE_9 [41:22];  
    
    assign  frontend_tlb_entries_barrier_4_io_y_ppn = frontend_tlb_entries_barrier_4_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_4_io_y_u = frontend_tlb_entries_barrier_4_io_x_u ; 
  assign  frontend_tlb_entries_barrier_4_io_y_g = frontend_tlb_entries_barrier_4_io_x_g ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_ptw = frontend_tlb_entries_barrier_4_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_final = frontend_tlb_entries_barrier_4_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ae_stage2 = frontend_tlb_entries_barrier_4_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pf = frontend_tlb_entries_barrier_4_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_4_io_y_gf = frontend_tlb_entries_barrier_4_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sw = frontend_tlb_entries_barrier_4_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sx = frontend_tlb_entries_barrier_4_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_4_io_y_sr = frontend_tlb_entries_barrier_4_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hw = frontend_tlb_entries_barrier_4_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hx = frontend_tlb_entries_barrier_4_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_4_io_y_hr = frontend_tlb_entries_barrier_4_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pw = frontend_tlb_entries_barrier_4_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_4_io_y_px = frontend_tlb_entries_barrier_4_io_x_px ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pr = frontend_tlb_entries_barrier_4_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_4_io_y_ppp = frontend_tlb_entries_barrier_4_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_4_io_y_pal = frontend_tlb_entries_barrier_4_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_4_io_y_paa = frontend_tlb_entries_barrier_4_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_4_io_y_eff = frontend_tlb_entries_barrier_4_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_4_io_y_c = frontend_tlb_entries_barrier_4_io_x_c ; 
  assign  frontend_tlb_entries_barrier_4_io_y_fragmented_superpage = frontend_tlb_entries_barrier_4_io_x_fragmented_superpage ;
     
    wire frontend_tlb__entries_WIRE_10_fragmented_superpage = frontend_tlb__entries_WIRE_11 [0]; 
    wire frontend_tlb__entries_WIRE_10_c = frontend_tlb__entries_WIRE_11 [1]; 
    wire frontend_tlb__entries_WIRE_10_eff = frontend_tlb__entries_WIRE_11 [2]; 
    wire frontend_tlb__entries_WIRE_10_paa = frontend_tlb__entries_WIRE_11 [3]; 
    wire frontend_tlb__entries_WIRE_10_pal = frontend_tlb__entries_WIRE_11 [4]; 
    wire frontend_tlb__entries_WIRE_10_ppp = frontend_tlb__entries_WIRE_11 [5]; 
    wire frontend_tlb__entries_WIRE_10_pr = frontend_tlb__entries_WIRE_11 [6]; 
    wire frontend_tlb__entries_WIRE_10_px = frontend_tlb__entries_WIRE_11 [7]; 
    wire frontend_tlb__entries_WIRE_10_pw = frontend_tlb__entries_WIRE_11 [8]; 
    wire frontend_tlb__entries_WIRE_10_hr = frontend_tlb__entries_WIRE_11 [9]; 
    wire frontend_tlb__entries_WIRE_10_hx = frontend_tlb__entries_WIRE_11 [10]; 
    wire frontend_tlb__entries_WIRE_10_hw = frontend_tlb__entries_WIRE_11 [11]; 
    wire frontend_tlb__entries_WIRE_10_sr = frontend_tlb__entries_WIRE_11 [12]; 
    wire frontend_tlb__entries_WIRE_10_sx = frontend_tlb__entries_WIRE_11 [13]; 
    wire frontend_tlb__entries_WIRE_10_sw = frontend_tlb__entries_WIRE_11 [14]; 
    wire frontend_tlb__entries_WIRE_10_gf = frontend_tlb__entries_WIRE_11 [15]; 
    wire frontend_tlb__entries_WIRE_10_pf = frontend_tlb__entries_WIRE_11 [16]; 
    wire frontend_tlb__entries_WIRE_10_ae_stage2 = frontend_tlb__entries_WIRE_11 [17]; 
    wire frontend_tlb__entries_WIRE_10_ae_final = frontend_tlb__entries_WIRE_11 [18]; 
    wire frontend_tlb__entries_WIRE_10_ae_ptw = frontend_tlb__entries_WIRE_11 [19]; 
    wire frontend_tlb__entries_WIRE_10_g = frontend_tlb__entries_WIRE_11 [20]; 
    wire frontend_tlb__entries_WIRE_10_u = frontend_tlb__entries_WIRE_11 [21]; 
    wire[19:0] frontend_tlb__entries_WIRE_10_ppn = frontend_tlb__entries_WIRE_11 [41:22];  
    
    assign  frontend_tlb_entries_barrier_5_io_y_ppn = frontend_tlb_entries_barrier_5_io_x_ppn ; 
  assign  frontend_tlb_entries_barrier_5_io_y_u = frontend_tlb_entries_barrier_5_io_x_u ; 
  assign  frontend_tlb_entries_barrier_5_io_y_g = frontend_tlb_entries_barrier_5_io_x_g ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_ptw = frontend_tlb_entries_barrier_5_io_x_ae_ptw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_final = frontend_tlb_entries_barrier_5_io_x_ae_final ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ae_stage2 = frontend_tlb_entries_barrier_5_io_x_ae_stage2 ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pf = frontend_tlb_entries_barrier_5_io_x_pf ; 
  assign  frontend_tlb_entries_barrier_5_io_y_gf = frontend_tlb_entries_barrier_5_io_x_gf ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sw = frontend_tlb_entries_barrier_5_io_x_sw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sx = frontend_tlb_entries_barrier_5_io_x_sx ; 
  assign  frontend_tlb_entries_barrier_5_io_y_sr = frontend_tlb_entries_barrier_5_io_x_sr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hw = frontend_tlb_entries_barrier_5_io_x_hw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hx = frontend_tlb_entries_barrier_5_io_x_hx ; 
  assign  frontend_tlb_entries_barrier_5_io_y_hr = frontend_tlb_entries_barrier_5_io_x_hr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pw = frontend_tlb_entries_barrier_5_io_x_pw ; 
  assign  frontend_tlb_entries_barrier_5_io_y_px = frontend_tlb_entries_barrier_5_io_x_px ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pr = frontend_tlb_entries_barrier_5_io_x_pr ; 
  assign  frontend_tlb_entries_barrier_5_io_y_ppp = frontend_tlb_entries_barrier_5_io_x_ppp ; 
  assign  frontend_tlb_entries_barrier_5_io_y_pal = frontend_tlb_entries_barrier_5_io_x_pal ; 
  assign  frontend_tlb_entries_barrier_5_io_y_paa = frontend_tlb_entries_barrier_5_io_x_paa ; 
  assign  frontend_tlb_entries_barrier_5_io_y_eff = frontend_tlb_entries_barrier_5_io_x_eff ; 
  assign  frontend_tlb_entries_barrier_5_io_y_c = frontend_tlb_entries_barrier_5_io_x_c ; 
  assign  frontend_tlb_entries_barrier_5_io_y_fragmented_superpage = frontend_tlb_entries_barrier_5_io_x_fragmented_superpage ;
    assign frontend_tlb_mpu_ppn_barrier_clock = frontend_tlb_clock;
    assign frontend_tlb_mpu_ppn_barrier_reset = frontend_tlb_reset;
    assign frontend_tlb_mpu_ppn_barrier_io_x_ppn = frontend_tlb__mpu_ppn_WIRE_ppn;
    assign frontend_tlb_mpu_ppn_barrier_io_x_u = frontend_tlb__mpu_ppn_WIRE_u;
    assign frontend_tlb_mpu_ppn_barrier_io_x_g = frontend_tlb__mpu_ppn_WIRE_g;
    assign frontend_tlb_mpu_ppn_barrier_io_x_ae_ptw = frontend_tlb__mpu_ppn_WIRE_ae_ptw;
    assign frontend_tlb_mpu_ppn_barrier_io_x_ae_final = frontend_tlb__mpu_ppn_WIRE_ae_final;
    assign frontend_tlb_mpu_ppn_barrier_io_x_ae_stage2 = frontend_tlb__mpu_ppn_WIRE_ae_stage2;
    assign frontend_tlb_mpu_ppn_barrier_io_x_pf = frontend_tlb__mpu_ppn_WIRE_pf;
    assign frontend_tlb_mpu_ppn_barrier_io_x_gf = frontend_tlb__mpu_ppn_WIRE_gf;
    assign frontend_tlb_mpu_ppn_barrier_io_x_sw = frontend_tlb__mpu_ppn_WIRE_sw;
    assign frontend_tlb_mpu_ppn_barrier_io_x_sx = frontend_tlb__mpu_ppn_WIRE_sx;
    assign frontend_tlb_mpu_ppn_barrier_io_x_sr = frontend_tlb__mpu_ppn_WIRE_sr;
    assign frontend_tlb_mpu_ppn_barrier_io_x_hw = frontend_tlb__mpu_ppn_WIRE_hw;
    assign frontend_tlb_mpu_ppn_barrier_io_x_hx = frontend_tlb__mpu_ppn_WIRE_hx;
    assign frontend_tlb_mpu_ppn_barrier_io_x_hr = frontend_tlb__mpu_ppn_WIRE_hr;
    assign frontend_tlb_mpu_ppn_barrier_io_x_pw = frontend_tlb__mpu_ppn_WIRE_pw;
    assign frontend_tlb_mpu_ppn_barrier_io_x_px = frontend_tlb__mpu_ppn_WIRE_px;
    assign frontend_tlb_mpu_ppn_barrier_io_x_pr = frontend_tlb__mpu_ppn_WIRE_pr;
    assign frontend_tlb_mpu_ppn_barrier_io_x_ppp = frontend_tlb__mpu_ppn_WIRE_ppp;
    assign frontend_tlb_mpu_ppn_barrier_io_x_pal = frontend_tlb__mpu_ppn_WIRE_pal;
    assign frontend_tlb_mpu_ppn_barrier_io_x_paa = frontend_tlb__mpu_ppn_WIRE_paa;
    assign frontend_tlb_mpu_ppn_barrier_io_x_eff = frontend_tlb__mpu_ppn_WIRE_eff;
    assign frontend_tlb_mpu_ppn_barrier_io_x_c = frontend_tlb__mpu_ppn_WIRE_c;
    assign frontend_tlb_mpu_ppn_barrier_io_x_fragmented_superpage = frontend_tlb__mpu_ppn_WIRE_fragmented_superpage;
    assign frontend_tlb__mpu_ppn_barrier_io_y_ppn = frontend_tlb_mpu_ppn_barrier_io_y_ppn;
    assign frontend_tlb_entries_barrier_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_io_x_ppn = frontend_tlb__entries_WIRE_ppn;
    assign frontend_tlb_entries_barrier_io_x_u = frontend_tlb__entries_WIRE_u;
    assign frontend_tlb_entries_barrier_io_x_g = frontend_tlb__entries_WIRE_g;
    assign frontend_tlb_entries_barrier_io_x_ae_ptw = frontend_tlb__entries_WIRE_ae_ptw;
    assign frontend_tlb_entries_barrier_io_x_ae_final = frontend_tlb__entries_WIRE_ae_final;
    assign frontend_tlb_entries_barrier_io_x_ae_stage2 = frontend_tlb__entries_WIRE_ae_stage2;
    assign frontend_tlb_entries_barrier_io_x_pf = frontend_tlb__entries_WIRE_pf;
    assign frontend_tlb_entries_barrier_io_x_gf = frontend_tlb__entries_WIRE_gf;
    assign frontend_tlb_entries_barrier_io_x_sw = frontend_tlb__entries_WIRE_sw;
    assign frontend_tlb_entries_barrier_io_x_sx = frontend_tlb__entries_WIRE_sx;
    assign frontend_tlb_entries_barrier_io_x_sr = frontend_tlb__entries_WIRE_sr;
    assign frontend_tlb_entries_barrier_io_x_hw = frontend_tlb__entries_WIRE_hw;
    assign frontend_tlb_entries_barrier_io_x_hx = frontend_tlb__entries_WIRE_hx;
    assign frontend_tlb_entries_barrier_io_x_hr = frontend_tlb__entries_WIRE_hr;
    assign frontend_tlb_entries_barrier_io_x_pw = frontend_tlb__entries_WIRE_pw;
    assign frontend_tlb_entries_barrier_io_x_px = frontend_tlb__entries_WIRE_px;
    assign frontend_tlb_entries_barrier_io_x_pr = frontend_tlb__entries_WIRE_pr;
    assign frontend_tlb_entries_barrier_io_x_ppp = frontend_tlb__entries_WIRE_ppp;
    assign frontend_tlb_entries_barrier_io_x_pal = frontend_tlb__entries_WIRE_pal;
    assign frontend_tlb_entries_barrier_io_x_paa = frontend_tlb__entries_WIRE_paa;
    assign frontend_tlb_entries_barrier_io_x_eff = frontend_tlb__entries_WIRE_eff;
    assign frontend_tlb_entries_barrier_io_x_c = frontend_tlb__entries_WIRE_c;
    assign frontend_tlb_entries_barrier_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_fragmented_superpage;
    assign frontend_tlb__entries_barrier_io_y_ppn = frontend_tlb_entries_barrier_io_y_ppn;
    assign frontend_tlb__entries_barrier_io_y_u = frontend_tlb_entries_barrier_io_y_u;
    assign frontend_tlb__entries_barrier_io_y_ae_ptw = frontend_tlb_entries_barrier_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_io_y_ae_final = frontend_tlb_entries_barrier_io_y_ae_final;
    assign frontend_tlb__entries_barrier_io_y_ae_stage2 = frontend_tlb_entries_barrier_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_io_y_pf = frontend_tlb_entries_barrier_io_y_pf;
    assign frontend_tlb__entries_barrier_io_y_gf = frontend_tlb_entries_barrier_io_y_gf;
    assign frontend_tlb__entries_barrier_io_y_sw = frontend_tlb_entries_barrier_io_y_sw;
    assign frontend_tlb__entries_barrier_io_y_sx = frontend_tlb_entries_barrier_io_y_sx;
    assign frontend_tlb__entries_barrier_io_y_sr = frontend_tlb_entries_barrier_io_y_sr;
    assign frontend_tlb__entries_barrier_io_y_hw = frontend_tlb_entries_barrier_io_y_hw;
    assign frontend_tlb__entries_barrier_io_y_hx = frontend_tlb_entries_barrier_io_y_hx;
    assign frontend_tlb__entries_barrier_io_y_hr = frontend_tlb_entries_barrier_io_y_hr;
    assign frontend_tlb__entries_barrier_io_y_pw = frontend_tlb_entries_barrier_io_y_pw;
    assign frontend_tlb__entries_barrier_io_y_px = frontend_tlb_entries_barrier_io_y_px;
    assign frontend_tlb__entries_barrier_io_y_pr = frontend_tlb_entries_barrier_io_y_pr;
    assign frontend_tlb__entries_barrier_io_y_ppp = frontend_tlb_entries_barrier_io_y_ppp;
    assign frontend_tlb__entries_barrier_io_y_pal = frontend_tlb_entries_barrier_io_y_pal;
    assign frontend_tlb__entries_barrier_io_y_paa = frontend_tlb_entries_barrier_io_y_paa;
    assign frontend_tlb__entries_barrier_io_y_eff = frontend_tlb_entries_barrier_io_y_eff;
    assign frontend_tlb__entries_barrier_io_y_c = frontend_tlb_entries_barrier_io_y_c;
    assign frontend_tlb_entries_barrier_1_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_1_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_1_io_x_ppn = frontend_tlb__entries_WIRE_2_ppn;
    assign frontend_tlb_entries_barrier_1_io_x_u = frontend_tlb__entries_WIRE_2_u;
    assign frontend_tlb_entries_barrier_1_io_x_g = frontend_tlb__entries_WIRE_2_g;
    assign frontend_tlb_entries_barrier_1_io_x_ae_ptw = frontend_tlb__entries_WIRE_2_ae_ptw;
    assign frontend_tlb_entries_barrier_1_io_x_ae_final = frontend_tlb__entries_WIRE_2_ae_final;
    assign frontend_tlb_entries_barrier_1_io_x_ae_stage2 = frontend_tlb__entries_WIRE_2_ae_stage2;
    assign frontend_tlb_entries_barrier_1_io_x_pf = frontend_tlb__entries_WIRE_2_pf;
    assign frontend_tlb_entries_barrier_1_io_x_gf = frontend_tlb__entries_WIRE_2_gf;
    assign frontend_tlb_entries_barrier_1_io_x_sw = frontend_tlb__entries_WIRE_2_sw;
    assign frontend_tlb_entries_barrier_1_io_x_sx = frontend_tlb__entries_WIRE_2_sx;
    assign frontend_tlb_entries_barrier_1_io_x_sr = frontend_tlb__entries_WIRE_2_sr;
    assign frontend_tlb_entries_barrier_1_io_x_hw = frontend_tlb__entries_WIRE_2_hw;
    assign frontend_tlb_entries_barrier_1_io_x_hx = frontend_tlb__entries_WIRE_2_hx;
    assign frontend_tlb_entries_barrier_1_io_x_hr = frontend_tlb__entries_WIRE_2_hr;
    assign frontend_tlb_entries_barrier_1_io_x_pw = frontend_tlb__entries_WIRE_2_pw;
    assign frontend_tlb_entries_barrier_1_io_x_px = frontend_tlb__entries_WIRE_2_px;
    assign frontend_tlb_entries_barrier_1_io_x_pr = frontend_tlb__entries_WIRE_2_pr;
    assign frontend_tlb_entries_barrier_1_io_x_ppp = frontend_tlb__entries_WIRE_2_ppp;
    assign frontend_tlb_entries_barrier_1_io_x_pal = frontend_tlb__entries_WIRE_2_pal;
    assign frontend_tlb_entries_barrier_1_io_x_paa = frontend_tlb__entries_WIRE_2_paa;
    assign frontend_tlb_entries_barrier_1_io_x_eff = frontend_tlb__entries_WIRE_2_eff;
    assign frontend_tlb_entries_barrier_1_io_x_c = frontend_tlb__entries_WIRE_2_c;
    assign frontend_tlb_entries_barrier_1_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_2_fragmented_superpage;
    assign frontend_tlb__entries_barrier_1_io_y_ppn = frontend_tlb_entries_barrier_1_io_y_ppn;
    assign frontend_tlb__entries_barrier_1_io_y_u = frontend_tlb_entries_barrier_1_io_y_u;
    assign frontend_tlb__entries_barrier_1_io_y_ae_ptw = frontend_tlb_entries_barrier_1_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_1_io_y_ae_final = frontend_tlb_entries_barrier_1_io_y_ae_final;
    assign frontend_tlb__entries_barrier_1_io_y_ae_stage2 = frontend_tlb_entries_barrier_1_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_1_io_y_pf = frontend_tlb_entries_barrier_1_io_y_pf;
    assign frontend_tlb__entries_barrier_1_io_y_gf = frontend_tlb_entries_barrier_1_io_y_gf;
    assign frontend_tlb__entries_barrier_1_io_y_sw = frontend_tlb_entries_barrier_1_io_y_sw;
    assign frontend_tlb__entries_barrier_1_io_y_sx = frontend_tlb_entries_barrier_1_io_y_sx;
    assign frontend_tlb__entries_barrier_1_io_y_sr = frontend_tlb_entries_barrier_1_io_y_sr;
    assign frontend_tlb__entries_barrier_1_io_y_hw = frontend_tlb_entries_barrier_1_io_y_hw;
    assign frontend_tlb__entries_barrier_1_io_y_hx = frontend_tlb_entries_barrier_1_io_y_hx;
    assign frontend_tlb__entries_barrier_1_io_y_hr = frontend_tlb_entries_barrier_1_io_y_hr;
    assign frontend_tlb__entries_barrier_1_io_y_pw = frontend_tlb_entries_barrier_1_io_y_pw;
    assign frontend_tlb__entries_barrier_1_io_y_px = frontend_tlb_entries_barrier_1_io_y_px;
    assign frontend_tlb__entries_barrier_1_io_y_pr = frontend_tlb_entries_barrier_1_io_y_pr;
    assign frontend_tlb__entries_barrier_1_io_y_ppp = frontend_tlb_entries_barrier_1_io_y_ppp;
    assign frontend_tlb__entries_barrier_1_io_y_pal = frontend_tlb_entries_barrier_1_io_y_pal;
    assign frontend_tlb__entries_barrier_1_io_y_paa = frontend_tlb_entries_barrier_1_io_y_paa;
    assign frontend_tlb__entries_barrier_1_io_y_eff = frontend_tlb_entries_barrier_1_io_y_eff;
    assign frontend_tlb__entries_barrier_1_io_y_c = frontend_tlb_entries_barrier_1_io_y_c;
    assign frontend_tlb_entries_barrier_2_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_2_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_2_io_x_ppn = frontend_tlb__entries_WIRE_4_ppn;
    assign frontend_tlb_entries_barrier_2_io_x_u = frontend_tlb__entries_WIRE_4_u;
    assign frontend_tlb_entries_barrier_2_io_x_g = frontend_tlb__entries_WIRE_4_g;
    assign frontend_tlb_entries_barrier_2_io_x_ae_ptw = frontend_tlb__entries_WIRE_4_ae_ptw;
    assign frontend_tlb_entries_barrier_2_io_x_ae_final = frontend_tlb__entries_WIRE_4_ae_final;
    assign frontend_tlb_entries_barrier_2_io_x_ae_stage2 = frontend_tlb__entries_WIRE_4_ae_stage2;
    assign frontend_tlb_entries_barrier_2_io_x_pf = frontend_tlb__entries_WIRE_4_pf;
    assign frontend_tlb_entries_barrier_2_io_x_gf = frontend_tlb__entries_WIRE_4_gf;
    assign frontend_tlb_entries_barrier_2_io_x_sw = frontend_tlb__entries_WIRE_4_sw;
    assign frontend_tlb_entries_barrier_2_io_x_sx = frontend_tlb__entries_WIRE_4_sx;
    assign frontend_tlb_entries_barrier_2_io_x_sr = frontend_tlb__entries_WIRE_4_sr;
    assign frontend_tlb_entries_barrier_2_io_x_hw = frontend_tlb__entries_WIRE_4_hw;
    assign frontend_tlb_entries_barrier_2_io_x_hx = frontend_tlb__entries_WIRE_4_hx;
    assign frontend_tlb_entries_barrier_2_io_x_hr = frontend_tlb__entries_WIRE_4_hr;
    assign frontend_tlb_entries_barrier_2_io_x_pw = frontend_tlb__entries_WIRE_4_pw;
    assign frontend_tlb_entries_barrier_2_io_x_px = frontend_tlb__entries_WIRE_4_px;
    assign frontend_tlb_entries_barrier_2_io_x_pr = frontend_tlb__entries_WIRE_4_pr;
    assign frontend_tlb_entries_barrier_2_io_x_ppp = frontend_tlb__entries_WIRE_4_ppp;
    assign frontend_tlb_entries_barrier_2_io_x_pal = frontend_tlb__entries_WIRE_4_pal;
    assign frontend_tlb_entries_barrier_2_io_x_paa = frontend_tlb__entries_WIRE_4_paa;
    assign frontend_tlb_entries_barrier_2_io_x_eff = frontend_tlb__entries_WIRE_4_eff;
    assign frontend_tlb_entries_barrier_2_io_x_c = frontend_tlb__entries_WIRE_4_c;
    assign frontend_tlb_entries_barrier_2_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_4_fragmented_superpage;
    assign frontend_tlb__entries_barrier_2_io_y_ppn = frontend_tlb_entries_barrier_2_io_y_ppn;
    assign frontend_tlb__entries_barrier_2_io_y_u = frontend_tlb_entries_barrier_2_io_y_u;
    assign frontend_tlb__entries_barrier_2_io_y_ae_ptw = frontend_tlb_entries_barrier_2_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_2_io_y_ae_final = frontend_tlb_entries_barrier_2_io_y_ae_final;
    assign frontend_tlb__entries_barrier_2_io_y_ae_stage2 = frontend_tlb_entries_barrier_2_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_2_io_y_pf = frontend_tlb_entries_barrier_2_io_y_pf;
    assign frontend_tlb__entries_barrier_2_io_y_gf = frontend_tlb_entries_barrier_2_io_y_gf;
    assign frontend_tlb__entries_barrier_2_io_y_sw = frontend_tlb_entries_barrier_2_io_y_sw;
    assign frontend_tlb__entries_barrier_2_io_y_sx = frontend_tlb_entries_barrier_2_io_y_sx;
    assign frontend_tlb__entries_barrier_2_io_y_sr = frontend_tlb_entries_barrier_2_io_y_sr;
    assign frontend_tlb__entries_barrier_2_io_y_hw = frontend_tlb_entries_barrier_2_io_y_hw;
    assign frontend_tlb__entries_barrier_2_io_y_hx = frontend_tlb_entries_barrier_2_io_y_hx;
    assign frontend_tlb__entries_barrier_2_io_y_hr = frontend_tlb_entries_barrier_2_io_y_hr;
    assign frontend_tlb__entries_barrier_2_io_y_pw = frontend_tlb_entries_barrier_2_io_y_pw;
    assign frontend_tlb__entries_barrier_2_io_y_px = frontend_tlb_entries_barrier_2_io_y_px;
    assign frontend_tlb__entries_barrier_2_io_y_pr = frontend_tlb_entries_barrier_2_io_y_pr;
    assign frontend_tlb__entries_barrier_2_io_y_ppp = frontend_tlb_entries_barrier_2_io_y_ppp;
    assign frontend_tlb__entries_barrier_2_io_y_pal = frontend_tlb_entries_barrier_2_io_y_pal;
    assign frontend_tlb__entries_barrier_2_io_y_paa = frontend_tlb_entries_barrier_2_io_y_paa;
    assign frontend_tlb__entries_barrier_2_io_y_eff = frontend_tlb_entries_barrier_2_io_y_eff;
    assign frontend_tlb__entries_barrier_2_io_y_c = frontend_tlb_entries_barrier_2_io_y_c;
    assign frontend_tlb_entries_barrier_3_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_3_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_3_io_x_ppn = frontend_tlb__entries_WIRE_6_ppn;
    assign frontend_tlb_entries_barrier_3_io_x_u = frontend_tlb__entries_WIRE_6_u;
    assign frontend_tlb_entries_barrier_3_io_x_g = frontend_tlb__entries_WIRE_6_g;
    assign frontend_tlb_entries_barrier_3_io_x_ae_ptw = frontend_tlb__entries_WIRE_6_ae_ptw;
    assign frontend_tlb_entries_barrier_3_io_x_ae_final = frontend_tlb__entries_WIRE_6_ae_final;
    assign frontend_tlb_entries_barrier_3_io_x_ae_stage2 = frontend_tlb__entries_WIRE_6_ae_stage2;
    assign frontend_tlb_entries_barrier_3_io_x_pf = frontend_tlb__entries_WIRE_6_pf;
    assign frontend_tlb_entries_barrier_3_io_x_gf = frontend_tlb__entries_WIRE_6_gf;
    assign frontend_tlb_entries_barrier_3_io_x_sw = frontend_tlb__entries_WIRE_6_sw;
    assign frontend_tlb_entries_barrier_3_io_x_sx = frontend_tlb__entries_WIRE_6_sx;
    assign frontend_tlb_entries_barrier_3_io_x_sr = frontend_tlb__entries_WIRE_6_sr;
    assign frontend_tlb_entries_barrier_3_io_x_hw = frontend_tlb__entries_WIRE_6_hw;
    assign frontend_tlb_entries_barrier_3_io_x_hx = frontend_tlb__entries_WIRE_6_hx;
    assign frontend_tlb_entries_barrier_3_io_x_hr = frontend_tlb__entries_WIRE_6_hr;
    assign frontend_tlb_entries_barrier_3_io_x_pw = frontend_tlb__entries_WIRE_6_pw;
    assign frontend_tlb_entries_barrier_3_io_x_px = frontend_tlb__entries_WIRE_6_px;
    assign frontend_tlb_entries_barrier_3_io_x_pr = frontend_tlb__entries_WIRE_6_pr;
    assign frontend_tlb_entries_barrier_3_io_x_ppp = frontend_tlb__entries_WIRE_6_ppp;
    assign frontend_tlb_entries_barrier_3_io_x_pal = frontend_tlb__entries_WIRE_6_pal;
    assign frontend_tlb_entries_barrier_3_io_x_paa = frontend_tlb__entries_WIRE_6_paa;
    assign frontend_tlb_entries_barrier_3_io_x_eff = frontend_tlb__entries_WIRE_6_eff;
    assign frontend_tlb_entries_barrier_3_io_x_c = frontend_tlb__entries_WIRE_6_c;
    assign frontend_tlb_entries_barrier_3_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_6_fragmented_superpage;
    assign frontend_tlb__entries_barrier_3_io_y_ppn = frontend_tlb_entries_barrier_3_io_y_ppn;
    assign frontend_tlb__entries_barrier_3_io_y_u = frontend_tlb_entries_barrier_3_io_y_u;
    assign frontend_tlb__entries_barrier_3_io_y_ae_ptw = frontend_tlb_entries_barrier_3_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_3_io_y_ae_final = frontend_tlb_entries_barrier_3_io_y_ae_final;
    assign frontend_tlb__entries_barrier_3_io_y_ae_stage2 = frontend_tlb_entries_barrier_3_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_3_io_y_pf = frontend_tlb_entries_barrier_3_io_y_pf;
    assign frontend_tlb__entries_barrier_3_io_y_gf = frontend_tlb_entries_barrier_3_io_y_gf;
    assign frontend_tlb__entries_barrier_3_io_y_sw = frontend_tlb_entries_barrier_3_io_y_sw;
    assign frontend_tlb__entries_barrier_3_io_y_sx = frontend_tlb_entries_barrier_3_io_y_sx;
    assign frontend_tlb__entries_barrier_3_io_y_sr = frontend_tlb_entries_barrier_3_io_y_sr;
    assign frontend_tlb__entries_barrier_3_io_y_hw = frontend_tlb_entries_barrier_3_io_y_hw;
    assign frontend_tlb__entries_barrier_3_io_y_hx = frontend_tlb_entries_barrier_3_io_y_hx;
    assign frontend_tlb__entries_barrier_3_io_y_hr = frontend_tlb_entries_barrier_3_io_y_hr;
    assign frontend_tlb__entries_barrier_3_io_y_pw = frontend_tlb_entries_barrier_3_io_y_pw;
    assign frontend_tlb__entries_barrier_3_io_y_px = frontend_tlb_entries_barrier_3_io_y_px;
    assign frontend_tlb__entries_barrier_3_io_y_pr = frontend_tlb_entries_barrier_3_io_y_pr;
    assign frontend_tlb__entries_barrier_3_io_y_ppp = frontend_tlb_entries_barrier_3_io_y_ppp;
    assign frontend_tlb__entries_barrier_3_io_y_pal = frontend_tlb_entries_barrier_3_io_y_pal;
    assign frontend_tlb__entries_barrier_3_io_y_paa = frontend_tlb_entries_barrier_3_io_y_paa;
    assign frontend_tlb__entries_barrier_3_io_y_eff = frontend_tlb_entries_barrier_3_io_y_eff;
    assign frontend_tlb__entries_barrier_3_io_y_c = frontend_tlb_entries_barrier_3_io_y_c;
    assign frontend_tlb_entries_barrier_4_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_4_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_4_io_x_ppn = frontend_tlb__entries_WIRE_8_ppn;
    assign frontend_tlb_entries_barrier_4_io_x_u = frontend_tlb__entries_WIRE_8_u;
    assign frontend_tlb_entries_barrier_4_io_x_g = frontend_tlb__entries_WIRE_8_g;
    assign frontend_tlb_entries_barrier_4_io_x_ae_ptw = frontend_tlb__entries_WIRE_8_ae_ptw;
    assign frontend_tlb_entries_barrier_4_io_x_ae_final = frontend_tlb__entries_WIRE_8_ae_final;
    assign frontend_tlb_entries_barrier_4_io_x_ae_stage2 = frontend_tlb__entries_WIRE_8_ae_stage2;
    assign frontend_tlb_entries_barrier_4_io_x_pf = frontend_tlb__entries_WIRE_8_pf;
    assign frontend_tlb_entries_barrier_4_io_x_gf = frontend_tlb__entries_WIRE_8_gf;
    assign frontend_tlb_entries_barrier_4_io_x_sw = frontend_tlb__entries_WIRE_8_sw;
    assign frontend_tlb_entries_barrier_4_io_x_sx = frontend_tlb__entries_WIRE_8_sx;
    assign frontend_tlb_entries_barrier_4_io_x_sr = frontend_tlb__entries_WIRE_8_sr;
    assign frontend_tlb_entries_barrier_4_io_x_hw = frontend_tlb__entries_WIRE_8_hw;
    assign frontend_tlb_entries_barrier_4_io_x_hx = frontend_tlb__entries_WIRE_8_hx;
    assign frontend_tlb_entries_barrier_4_io_x_hr = frontend_tlb__entries_WIRE_8_hr;
    assign frontend_tlb_entries_barrier_4_io_x_pw = frontend_tlb__entries_WIRE_8_pw;
    assign frontend_tlb_entries_barrier_4_io_x_px = frontend_tlb__entries_WIRE_8_px;
    assign frontend_tlb_entries_barrier_4_io_x_pr = frontend_tlb__entries_WIRE_8_pr;
    assign frontend_tlb_entries_barrier_4_io_x_ppp = frontend_tlb__entries_WIRE_8_ppp;
    assign frontend_tlb_entries_barrier_4_io_x_pal = frontend_tlb__entries_WIRE_8_pal;
    assign frontend_tlb_entries_barrier_4_io_x_paa = frontend_tlb__entries_WIRE_8_paa;
    assign frontend_tlb_entries_barrier_4_io_x_eff = frontend_tlb__entries_WIRE_8_eff;
    assign frontend_tlb_entries_barrier_4_io_x_c = frontend_tlb__entries_WIRE_8_c;
    assign frontend_tlb_entries_barrier_4_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_8_fragmented_superpage;
    assign frontend_tlb__entries_barrier_4_io_y_ppn = frontend_tlb_entries_barrier_4_io_y_ppn;
    assign frontend_tlb__entries_barrier_4_io_y_u = frontend_tlb_entries_barrier_4_io_y_u;
    assign frontend_tlb__entries_barrier_4_io_y_ae_ptw = frontend_tlb_entries_barrier_4_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_4_io_y_ae_final = frontend_tlb_entries_barrier_4_io_y_ae_final;
    assign frontend_tlb__entries_barrier_4_io_y_ae_stage2 = frontend_tlb_entries_barrier_4_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_4_io_y_pf = frontend_tlb_entries_barrier_4_io_y_pf;
    assign frontend_tlb__entries_barrier_4_io_y_gf = frontend_tlb_entries_barrier_4_io_y_gf;
    assign frontend_tlb__entries_barrier_4_io_y_sw = frontend_tlb_entries_barrier_4_io_y_sw;
    assign frontend_tlb__entries_barrier_4_io_y_sx = frontend_tlb_entries_barrier_4_io_y_sx;
    assign frontend_tlb__entries_barrier_4_io_y_sr = frontend_tlb_entries_barrier_4_io_y_sr;
    assign frontend_tlb__entries_barrier_4_io_y_hw = frontend_tlb_entries_barrier_4_io_y_hw;
    assign frontend_tlb__entries_barrier_4_io_y_hx = frontend_tlb_entries_barrier_4_io_y_hx;
    assign frontend_tlb__entries_barrier_4_io_y_hr = frontend_tlb_entries_barrier_4_io_y_hr;
    assign frontend_tlb__entries_barrier_4_io_y_pw = frontend_tlb_entries_barrier_4_io_y_pw;
    assign frontend_tlb__entries_barrier_4_io_y_px = frontend_tlb_entries_barrier_4_io_y_px;
    assign frontend_tlb__entries_barrier_4_io_y_pr = frontend_tlb_entries_barrier_4_io_y_pr;
    assign frontend_tlb__entries_barrier_4_io_y_ppp = frontend_tlb_entries_barrier_4_io_y_ppp;
    assign frontend_tlb__entries_barrier_4_io_y_pal = frontend_tlb_entries_barrier_4_io_y_pal;
    assign frontend_tlb__entries_barrier_4_io_y_paa = frontend_tlb_entries_barrier_4_io_y_paa;
    assign frontend_tlb__entries_barrier_4_io_y_eff = frontend_tlb_entries_barrier_4_io_y_eff;
    assign frontend_tlb__entries_barrier_4_io_y_c = frontend_tlb_entries_barrier_4_io_y_c;
    assign frontend_tlb_entries_barrier_5_clock = frontend_tlb_clock;
    assign frontend_tlb_entries_barrier_5_reset = frontend_tlb_reset;
    assign frontend_tlb_entries_barrier_5_io_x_ppn = frontend_tlb__entries_WIRE_10_ppn;
    assign frontend_tlb_entries_barrier_5_io_x_u = frontend_tlb__entries_WIRE_10_u;
    assign frontend_tlb_entries_barrier_5_io_x_g = frontend_tlb__entries_WIRE_10_g;
    assign frontend_tlb_entries_barrier_5_io_x_ae_ptw = frontend_tlb__entries_WIRE_10_ae_ptw;
    assign frontend_tlb_entries_barrier_5_io_x_ae_final = frontend_tlb__entries_WIRE_10_ae_final;
    assign frontend_tlb_entries_barrier_5_io_x_ae_stage2 = frontend_tlb__entries_WIRE_10_ae_stage2;
    assign frontend_tlb_entries_barrier_5_io_x_pf = frontend_tlb__entries_WIRE_10_pf;
    assign frontend_tlb_entries_barrier_5_io_x_gf = frontend_tlb__entries_WIRE_10_gf;
    assign frontend_tlb_entries_barrier_5_io_x_sw = frontend_tlb__entries_WIRE_10_sw;
    assign frontend_tlb_entries_barrier_5_io_x_sx = frontend_tlb__entries_WIRE_10_sx;
    assign frontend_tlb_entries_barrier_5_io_x_sr = frontend_tlb__entries_WIRE_10_sr;
    assign frontend_tlb_entries_barrier_5_io_x_hw = frontend_tlb__entries_WIRE_10_hw;
    assign frontend_tlb_entries_barrier_5_io_x_hx = frontend_tlb__entries_WIRE_10_hx;
    assign frontend_tlb_entries_barrier_5_io_x_hr = frontend_tlb__entries_WIRE_10_hr;
    assign frontend_tlb_entries_barrier_5_io_x_pw = frontend_tlb__entries_WIRE_10_pw;
    assign frontend_tlb_entries_barrier_5_io_x_px = frontend_tlb__entries_WIRE_10_px;
    assign frontend_tlb_entries_barrier_5_io_x_pr = frontend_tlb__entries_WIRE_10_pr;
    assign frontend_tlb_entries_barrier_5_io_x_ppp = frontend_tlb__entries_WIRE_10_ppp;
    assign frontend_tlb_entries_barrier_5_io_x_pal = frontend_tlb__entries_WIRE_10_pal;
    assign frontend_tlb_entries_barrier_5_io_x_paa = frontend_tlb__entries_WIRE_10_paa;
    assign frontend_tlb_entries_barrier_5_io_x_eff = frontend_tlb__entries_WIRE_10_eff;
    assign frontend_tlb_entries_barrier_5_io_x_c = frontend_tlb__entries_WIRE_10_c;
    assign frontend_tlb_entries_barrier_5_io_x_fragmented_superpage = frontend_tlb__entries_WIRE_10_fragmented_superpage;
    assign frontend_tlb__entries_barrier_5_io_y_ppn = frontend_tlb_entries_barrier_5_io_y_ppn;
    assign frontend_tlb__entries_barrier_5_io_y_u = frontend_tlb_entries_barrier_5_io_y_u;
    assign frontend_tlb__entries_barrier_5_io_y_ae_ptw = frontend_tlb_entries_barrier_5_io_y_ae_ptw;
    assign frontend_tlb__entries_barrier_5_io_y_ae_final = frontend_tlb_entries_barrier_5_io_y_ae_final;
    assign frontend_tlb__entries_barrier_5_io_y_ae_stage2 = frontend_tlb_entries_barrier_5_io_y_ae_stage2;
    assign frontend_tlb__entries_barrier_5_io_y_pf = frontend_tlb_entries_barrier_5_io_y_pf;
    assign frontend_tlb__entries_barrier_5_io_y_gf = frontend_tlb_entries_barrier_5_io_y_gf;
    assign frontend_tlb__entries_barrier_5_io_y_sw = frontend_tlb_entries_barrier_5_io_y_sw;
    assign frontend_tlb__entries_barrier_5_io_y_sx = frontend_tlb_entries_barrier_5_io_y_sx;
    assign frontend_tlb__entries_barrier_5_io_y_sr = frontend_tlb_entries_barrier_5_io_y_sr;
    assign frontend_tlb__entries_barrier_5_io_y_hw = frontend_tlb_entries_barrier_5_io_y_hw;
    assign frontend_tlb__entries_barrier_5_io_y_hx = frontend_tlb_entries_barrier_5_io_y_hx;
    assign frontend_tlb__entries_barrier_5_io_y_hr = frontend_tlb_entries_barrier_5_io_y_hr;
     
    wire[19:0] frontend_tlb_ppn =( frontend_tlb_hitsVec_0  ?  frontend_tlb__entries_barrier_io_y_ppn :20'h0)|( frontend_tlb_hitsVec_1  ?  frontend_tlb__entries_barrier_1_io_y_ppn :20'h0)|( frontend_tlb_hitsVec_2  ?  frontend_tlb__entries_barrier_2_io_y_ppn :20'h0)|( frontend_tlb_hitsVec_3  ?  frontend_tlb__entries_barrier_3_io_y_ppn :20'h0)|( frontend_tlb_hitsVec_4  ?  frontend_tlb__entries_barrier_4_io_y_ppn :20'h0)|( frontend_tlb_hitsVec_5  ?  frontend_tlb__entries_barrier_5_io_y_ppn :20'h0)|( frontend_tlb_vm_enabled ==1'h0 ?  frontend_tlb_vpn [19:0]:20'h0); 
    wire[1:0] frontend_tlb_ptw_ae_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_ptw , frontend_tlb__entries_barrier_1_io_y_ae_ptw }; 
    wire[2:0] frontend_tlb_ptw_ae_array_lo ={ frontend_tlb_ptw_ae_array_lo_hi , frontend_tlb__entries_barrier_io_y_ae_ptw }; 
    wire[1:0] frontend_tlb_ptw_ae_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_ptw , frontend_tlb__entries_barrier_4_io_y_ae_ptw }; 
    wire[2:0] frontend_tlb_ptw_ae_array_hi ={ frontend_tlb_ptw_ae_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_ptw }; 
    wire[6:0] frontend_tlb_ptw_ae_array ={1'h0,{ frontend_tlb_ptw_ae_array_hi , frontend_tlb_ptw_ae_array_lo }}; 
    wire[1:0] frontend_tlb_final_ae_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_final , frontend_tlb__entries_barrier_1_io_y_ae_final }; 
    wire[2:0] frontend_tlb_final_ae_array_lo ={ frontend_tlb_final_ae_array_lo_hi , frontend_tlb__entries_barrier_io_y_ae_final }; 
    wire[1:0] frontend_tlb_final_ae_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_final , frontend_tlb__entries_barrier_4_io_y_ae_final }; 
    wire[2:0] frontend_tlb_final_ae_array_hi ={ frontend_tlb_final_ae_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_final }; 
    wire[6:0] frontend_tlb_final_ae_array ={1'h0,{ frontend_tlb_final_ae_array_hi , frontend_tlb_final_ae_array_lo }}; 
    wire[1:0] frontend_tlb_ptw_pf_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_pf , frontend_tlb__entries_barrier_1_io_y_pf }; 
    wire[2:0] frontend_tlb_ptw_pf_array_lo ={ frontend_tlb_ptw_pf_array_lo_hi , frontend_tlb__entries_barrier_io_y_pf }; 
    wire[1:0] frontend_tlb_ptw_pf_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_pf , frontend_tlb__entries_barrier_4_io_y_pf }; 
    wire[2:0] frontend_tlb_ptw_pf_array_hi ={ frontend_tlb_ptw_pf_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_pf }; 
    wire[6:0] frontend_tlb_ptw_pf_array ={1'h0,{ frontend_tlb_ptw_pf_array_hi , frontend_tlb_ptw_pf_array_lo }}; 
    wire[1:0] frontend_tlb_ptw_gf_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_gf , frontend_tlb__entries_barrier_1_io_y_gf }; 
    wire[2:0] frontend_tlb_ptw_gf_array_lo ={ frontend_tlb_ptw_gf_array_lo_hi , frontend_tlb__entries_barrier_io_y_gf }; 
    wire[1:0] frontend_tlb_ptw_gf_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_gf , frontend_tlb__entries_barrier_4_io_y_gf }; 
    wire[2:0] frontend_tlb_ptw_gf_array_hi ={ frontend_tlb_ptw_gf_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_gf }; 
    wire[6:0] frontend_tlb_ptw_gf_array ={1'h0,{ frontend_tlb_ptw_gf_array_hi , frontend_tlb_ptw_gf_array_lo }}; 
    wire frontend_tlb_sum = frontend_tlb_priv_v  ?  frontend_tlb_io_ptw_gstatus_sum : frontend_tlb_io_ptw_status_sum ; 
    wire[1:0] frontend_tlb_priv_rw_ok_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_u , frontend_tlb__entries_barrier_1_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_lo ={ frontend_tlb_priv_rw_ok_lo_hi , frontend_tlb__entries_barrier_io_y_u }; 
    wire[1:0] frontend_tlb_priv_rw_ok_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_u , frontend_tlb__entries_barrier_4_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_hi ={ frontend_tlb_priv_rw_ok_hi_hi , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[1:0] frontend_tlb_priv_rw_ok_lo_hi_1 ={ frontend_tlb__entries_barrier_2_io_y_u , frontend_tlb__entries_barrier_1_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_lo_1 ={ frontend_tlb_priv_rw_ok_lo_hi_1 , frontend_tlb__entries_barrier_io_y_u }; 
    wire[1:0] frontend_tlb_priv_rw_ok_hi_hi_1 ={ frontend_tlb__entries_barrier_5_io_y_u , frontend_tlb__entries_barrier_4_io_y_u }; 
    wire[2:0] frontend_tlb_priv_rw_ok_hi_1 ={ frontend_tlb_priv_rw_ok_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[5:0] frontend_tlb_priv_rw_ok =( frontend_tlb_priv_s ==1'h0| frontend_tlb_sum  ? { frontend_tlb_priv_rw_ok_hi , frontend_tlb_priv_rw_ok_lo }:6'h0)|( frontend_tlb_priv_s  ? ~{ frontend_tlb_priv_rw_ok_hi_1 , frontend_tlb_priv_rw_ok_lo_1 }:6'h0); 
    wire[1:0] frontend_tlb_priv_x_ok_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_u , frontend_tlb__entries_barrier_1_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_lo ={ frontend_tlb_priv_x_ok_lo_hi , frontend_tlb__entries_barrier_io_y_u }; 
    wire[1:0] frontend_tlb_priv_x_ok_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_u , frontend_tlb__entries_barrier_4_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_hi ={ frontend_tlb_priv_x_ok_hi_hi , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[1:0] frontend_tlb_priv_x_ok_lo_hi_1 ={ frontend_tlb__entries_barrier_2_io_y_u , frontend_tlb__entries_barrier_1_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_lo_1 ={ frontend_tlb_priv_x_ok_lo_hi_1 , frontend_tlb__entries_barrier_io_y_u }; 
    wire[1:0] frontend_tlb_priv_x_ok_hi_hi_1 ={ frontend_tlb__entries_barrier_5_io_y_u , frontend_tlb__entries_barrier_4_io_y_u }; 
    wire[2:0] frontend_tlb_priv_x_ok_hi_1 ={ frontend_tlb_priv_x_ok_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_u }; 
    wire[5:0] frontend_tlb_priv_x_ok = frontend_tlb_priv_s  ? ~{ frontend_tlb_priv_x_ok_hi , frontend_tlb_priv_x_ok_lo }:{ frontend_tlb_priv_x_ok_hi_1 , frontend_tlb_priv_x_ok_lo_1 }; 
    wire[1:0] frontend_tlb_stage1_bypass_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_ae_stage2 , frontend_tlb__entries_barrier_1_io_y_ae_stage2 }; 
    wire[2:0] frontend_tlb_stage1_bypass_lo ={ frontend_tlb_stage1_bypass_lo_hi , frontend_tlb__entries_barrier_io_y_ae_stage2 }; 
    wire[1:0] frontend_tlb_stage1_bypass_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_ae_stage2 , frontend_tlb__entries_barrier_4_io_y_ae_stage2 }; 
    wire[2:0] frontend_tlb_stage1_bypass_hi ={ frontend_tlb_stage1_bypass_hi_hi , frontend_tlb__entries_barrier_3_io_y_ae_stage2 }; 
    wire frontend_tlb_mxr = frontend_tlb_io_ptw_status_mxr |( frontend_tlb_priv_v  ?  frontend_tlb_io_ptw_gstatus_mxr :1'h0); 
    wire[1:0] frontend_tlb_r_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_sr , frontend_tlb__entries_barrier_1_io_y_sr }; 
    wire[2:0] frontend_tlb_r_array_lo ={ frontend_tlb_r_array_lo_hi , frontend_tlb__entries_barrier_io_y_sr }; 
    wire[1:0] frontend_tlb_r_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_sr , frontend_tlb__entries_barrier_4_io_y_sr }; 
    wire[2:0] frontend_tlb_r_array_hi ={ frontend_tlb_r_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sr }; 
    wire[1:0] frontend_tlb_r_array_lo_hi_1 ={ frontend_tlb__entries_barrier_2_io_y_sx , frontend_tlb__entries_barrier_1_io_y_sx }; 
    wire[2:0] frontend_tlb_r_array_lo_1 ={ frontend_tlb_r_array_lo_hi_1 , frontend_tlb__entries_barrier_io_y_sx }; 
    wire[1:0] frontend_tlb_r_array_hi_hi_1 ={ frontend_tlb__entries_barrier_5_io_y_sx , frontend_tlb__entries_barrier_4_io_y_sx }; 
    wire[2:0] frontend_tlb_r_array_hi_1 ={ frontend_tlb_r_array_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_sx }; 
    wire[6:0] frontend_tlb_r_array ={1'h1, frontend_tlb_priv_rw_ok &({ frontend_tlb_r_array_hi , frontend_tlb_r_array_lo }|( frontend_tlb_mxr  ? { frontend_tlb_r_array_hi_1 , frontend_tlb_r_array_lo_1 }:6'h0))| frontend_tlb_stage1_bypass }; 
    wire[1:0] frontend_tlb_w_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_sw , frontend_tlb__entries_barrier_1_io_y_sw }; 
    wire[2:0] frontend_tlb_w_array_lo ={ frontend_tlb_w_array_lo_hi , frontend_tlb__entries_barrier_io_y_sw }; 
    wire[1:0] frontend_tlb_w_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_sw , frontend_tlb__entries_barrier_4_io_y_sw }; 
    wire[2:0] frontend_tlb_w_array_hi ={ frontend_tlb_w_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sw }; 
    wire[6:0] frontend_tlb_w_array ={1'h1, frontend_tlb_priv_rw_ok &{ frontend_tlb_w_array_hi , frontend_tlb_w_array_lo }| frontend_tlb_stage1_bypass }; 
    wire[1:0] frontend_tlb_x_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_sx , frontend_tlb__entries_barrier_1_io_y_sx }; 
    wire[2:0] frontend_tlb_x_array_lo ={ frontend_tlb_x_array_lo_hi , frontend_tlb__entries_barrier_io_y_sx }; 
    wire[1:0] frontend_tlb_x_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_sx , frontend_tlb__entries_barrier_4_io_y_sx }; 
    wire[2:0] frontend_tlb_x_array_hi ={ frontend_tlb_x_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_sx }; 
    wire[6:0] frontend_tlb_x_array ={1'h1, frontend_tlb_priv_x_ok &{ frontend_tlb_x_array_hi , frontend_tlb_x_array_lo }| frontend_tlb_stage1_bypass }; 
    wire[5:0] frontend_tlb_stage2_bypass = frontend_tlb_stage2_en ==1'h0 ? 6'h3F:6'h0; 
    wire[1:0] frontend_tlb_hr_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_hr , frontend_tlb__entries_barrier_1_io_y_hr }; 
    wire[2:0] frontend_tlb_hr_array_lo ={ frontend_tlb_hr_array_lo_hi , frontend_tlb__entries_barrier_io_y_hr }; 
    wire[1:0] frontend_tlb_hr_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_hr , frontend_tlb__entries_barrier_4_io_y_hr }; 
    wire[2:0] frontend_tlb_hr_array_hi ={ frontend_tlb_hr_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hr }; 
    wire[1:0] frontend_tlb_hr_array_lo_hi_1 ={ frontend_tlb__entries_barrier_2_io_y_hx , frontend_tlb__entries_barrier_1_io_y_hx }; 
    wire[2:0] frontend_tlb_hr_array_lo_1 ={ frontend_tlb_hr_array_lo_hi_1 , frontend_tlb__entries_barrier_io_y_hx }; 
    wire[1:0] frontend_tlb_hr_array_hi_hi_1 ={ frontend_tlb__entries_barrier_5_io_y_hx , frontend_tlb__entries_barrier_4_io_y_hx }; 
    wire[2:0] frontend_tlb_hr_array_hi_1 ={ frontend_tlb_hr_array_hi_hi_1 , frontend_tlb__entries_barrier_3_io_y_hx }; 
    wire[6:0] frontend_tlb_hr_array ={1'h1,{ frontend_tlb_hr_array_hi , frontend_tlb_hr_array_lo }|( frontend_tlb_io_ptw_status_mxr  ? { frontend_tlb_hr_array_hi_1 , frontend_tlb_hr_array_lo_1 }:6'h0)| frontend_tlb_stage2_bypass }; 
    wire[1:0] frontend_tlb_hw_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_hw , frontend_tlb__entries_barrier_1_io_y_hw }; 
    wire[2:0] frontend_tlb_hw_array_lo ={ frontend_tlb_hw_array_lo_hi , frontend_tlb__entries_barrier_io_y_hw }; 
    wire[1:0] frontend_tlb_hw_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_hw , frontend_tlb__entries_barrier_4_io_y_hw }; 
    wire[2:0] frontend_tlb_hw_array_hi ={ frontend_tlb_hw_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hw }; 
    wire[6:0] frontend_tlb_hw_array ={1'h1,{ frontend_tlb_hw_array_hi , frontend_tlb_hw_array_lo }| frontend_tlb_stage2_bypass }; 
    wire[1:0] frontend_tlb_hx_array_lo_hi ={ frontend_tlb__entries_barrier_2_io_y_hx , frontend_tlb__entries_barrier_1_io_y_hx }; 
    wire[2:0] frontend_tlb_hx_array_lo ={ frontend_tlb_hx_array_lo_hi , frontend_tlb__entries_barrier_io_y_hx }; 
    wire[1:0] frontend_tlb_hx_array_hi_hi ={ frontend_tlb__entries_barrier_5_io_y_hx , frontend_tlb__entries_barrier_4_io_y_hx }; 
    wire[2:0] frontend_tlb_hx_array_hi ={ frontend_tlb_hx_array_hi_hi , frontend_tlb__entries_barrier_3_io_y_hx }; 
    wire[6:0] frontend_tlb_hx_array ={1'h1,{ frontend_tlb_hx_array_hi , frontend_tlb_hx_array_lo }| frontend_tlb_stage2_bypass }; 
    wire[1:0] frontend_tlb_pr_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pr , frontend_tlb__entries_barrier_io_y_pr }; 
    wire[1:0] frontend_tlb_pr_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pr , frontend_tlb__entries_barrier_3_io_y_pr }; 
    wire[2:0] frontend_tlb_pr_array_hi ={ frontend_tlb_pr_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pr }; 
    wire[6:0] frontend_tlb_pr_array ={ frontend_tlb_prot_r  ? 2'h3:2'h0,{ frontend_tlb_pr_array_hi , frontend_tlb_pr_array_lo }}&~( frontend_tlb_ptw_ae_array | frontend_tlb_final_ae_array ); 
    wire[1:0] frontend_tlb_pw_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pw , frontend_tlb__entries_barrier_io_y_pw }; 
    wire[1:0] frontend_tlb_pw_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pw , frontend_tlb__entries_barrier_3_io_y_pw }; 
    wire[2:0] frontend_tlb_pw_array_hi ={ frontend_tlb_pw_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pw }; 
    wire[6:0] frontend_tlb_pw_array ={ frontend_tlb_prot_w  ? 2'h3:2'h0,{ frontend_tlb_pw_array_hi , frontend_tlb_pw_array_lo }}&~( frontend_tlb_ptw_ae_array | frontend_tlb_final_ae_array ); 
    wire[1:0] frontend_tlb_px_array_lo ={ frontend_tlb__entries_barrier_1_io_y_px , frontend_tlb__entries_barrier_io_y_px }; 
    wire[1:0] frontend_tlb_px_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_px , frontend_tlb__entries_barrier_3_io_y_px }; 
    wire[2:0] frontend_tlb_px_array_hi ={ frontend_tlb_px_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_px }; 
    wire[6:0] frontend_tlb_px_array ={ frontend_tlb_prot_x  ? 2'h3:2'h0,{ frontend_tlb_px_array_hi , frontend_tlb_px_array_lo }}&~( frontend_tlb_ptw_ae_array | frontend_tlb_final_ae_array ); 
    wire[1:0] frontend_tlb_eff_array_lo ={ frontend_tlb__entries_barrier_1_io_y_eff , frontend_tlb__entries_barrier_io_y_eff }; 
    wire[1:0] frontend_tlb_eff_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_eff , frontend_tlb__entries_barrier_3_io_y_eff }; 
    wire[2:0] frontend_tlb_eff_array_hi ={ frontend_tlb_eff_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_eff }; 
    wire[6:0] frontend_tlb_eff_array ={ frontend_tlb_prot_eff  ? 2'h3:2'h0,{ frontend_tlb_eff_array_hi , frontend_tlb_eff_array_lo }}; 
    wire[1:0] frontend_tlb_c_array_lo ={ frontend_tlb__entries_barrier_1_io_y_c , frontend_tlb__entries_barrier_io_y_c }; 
    wire[1:0] frontend_tlb_c_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_c , frontend_tlb__entries_barrier_3_io_y_c }; 
    wire[2:0] frontend_tlb_c_array_hi ={ frontend_tlb_c_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_c }; 
    wire[6:0] frontend_tlb_c_array ={ frontend_tlb_cacheable  ? 2'h3:2'h0,{ frontend_tlb_c_array_hi , frontend_tlb_c_array_lo }}; 
    wire[6:0] frontend_tlb_lrscAllowed = frontend_tlb_c_array ; 
    wire[1:0] frontend_tlb_ppp_array_lo ={ frontend_tlb__entries_barrier_1_io_y_ppp , frontend_tlb__entries_barrier_io_y_ppp }; 
    wire[1:0] frontend_tlb_ppp_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_ppp , frontend_tlb__entries_barrier_3_io_y_ppp }; 
    wire[2:0] frontend_tlb_ppp_array_hi ={ frontend_tlb_ppp_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_ppp }; 
    wire[6:0] frontend_tlb_ppp_array ={ frontend_tlb_prot_pp  ? 2'h3:2'h0,{ frontend_tlb_ppp_array_hi , frontend_tlb_ppp_array_lo }}; 
    wire[1:0] frontend_tlb_paa_array_lo ={ frontend_tlb__entries_barrier_1_io_y_paa , frontend_tlb__entries_barrier_io_y_paa }; 
    wire[1:0] frontend_tlb_paa_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_paa , frontend_tlb__entries_barrier_3_io_y_paa }; 
    wire[2:0] frontend_tlb_paa_array_hi ={ frontend_tlb_paa_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_paa }; 
    wire[6:0] frontend_tlb_paa_array ={ frontend_tlb_prot_aa  ? 2'h3:2'h0,{ frontend_tlb_paa_array_hi , frontend_tlb_paa_array_lo }}; 
    wire[1:0] frontend_tlb_pal_array_lo ={ frontend_tlb__entries_barrier_1_io_y_pal , frontend_tlb__entries_barrier_io_y_pal }; 
    wire[1:0] frontend_tlb_pal_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_pal , frontend_tlb__entries_barrier_3_io_y_pal }; 
    wire[2:0] frontend_tlb_pal_array_hi ={ frontend_tlb_pal_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_pal }; 
    wire[6:0] frontend_tlb_pal_array ={ frontend_tlb_prot_al  ? 2'h3:2'h0,{ frontend_tlb_pal_array_hi , frontend_tlb_pal_array_lo }}; 
    wire[6:0] frontend_tlb_ppp_array_if_cached = frontend_tlb_ppp_array | frontend_tlb_c_array ; 
    wire[6:0] frontend_tlb_paa_array_if_cached = frontend_tlb_paa_array | frontend_tlb_c_array ; 
    wire[6:0] frontend_tlb_pal_array_if_cached = frontend_tlb_pal_array | frontend_tlb_c_array ; 
    wire[1:0] frontend_tlb_prefetchable_array_lo ={ frontend_tlb__entries_barrier_1_io_y_c , frontend_tlb__entries_barrier_io_y_c }; 
    wire[1:0] frontend_tlb_prefetchable_array_hi_hi ={ frontend_tlb__entries_barrier_4_io_y_c , frontend_tlb__entries_barrier_3_io_y_c }; 
    wire[2:0] frontend_tlb_prefetchable_array_hi ={ frontend_tlb_prefetchable_array_hi_hi , frontend_tlb__entries_barrier_2_io_y_c }; 
    wire[6:0] frontend_tlb_prefetchable_array ={{ frontend_tlb_cacheable & frontend_tlb_homogeneous ,1'h0},{ frontend_tlb_prefetchable_array_hi , frontend_tlb_prefetchable_array_lo }}; 
    wire[4:0] frontend_tlb__GEN_33 ={1'h0,4'h1<< frontend_tlb_io_req_bits_size }-5'h1; 
    wire frontend_tlb_misaligned =|( frontend_tlb_io_req_bits_vaddr &{30'h0, frontend_tlb__GEN_33 [3:0]}); 
    wire frontend_tlb_cmd_lrsc =( frontend_tlb_io_req_bits_cmd ==5'h6| frontend_tlb_io_req_bits_cmd ==5'h7)&1'h1; 
    wire frontend_tlb_cmd_amo_logical =( frontend_tlb_io_req_bits_cmd ==5'h4| frontend_tlb_io_req_bits_cmd ==5'h9| frontend_tlb_io_req_bits_cmd ==5'hA| frontend_tlb_io_req_bits_cmd ==5'hB)&1'h1; 
    wire frontend_tlb_cmd_amo_arithmetic =( frontend_tlb_io_req_bits_cmd ==5'h8| frontend_tlb_io_req_bits_cmd ==5'hC| frontend_tlb_io_req_bits_cmd ==5'hD| frontend_tlb_io_req_bits_cmd ==5'hE| frontend_tlb_io_req_bits_cmd ==5'hF)&1'h1; 
    wire frontend_tlb_cmd_put_partial = frontend_tlb_io_req_bits_cmd ==5'h11; 
    wire frontend_tlb_cmd_read = frontend_tlb_io_req_bits_cmd ==5'h0| frontend_tlb_io_req_bits_cmd ==5'h10| frontend_tlb_io_req_bits_cmd ==5'h6| frontend_tlb_io_req_bits_cmd ==5'h7| frontend_tlb_io_req_bits_cmd ==5'h4| frontend_tlb_io_req_bits_cmd ==5'h9| frontend_tlb_io_req_bits_cmd ==5'hA| frontend_tlb_io_req_bits_cmd ==5'hB| frontend_tlb_io_req_bits_cmd ==5'h8| frontend_tlb_io_req_bits_cmd ==5'hC| frontend_tlb_io_req_bits_cmd ==5'hD| frontend_tlb_io_req_bits_cmd ==5'hE| frontend_tlb_io_req_bits_cmd ==5'hF; 
    wire frontend_tlb_cmd_write = frontend_tlb_io_req_bits_cmd ==5'h1| frontend_tlb_io_req_bits_cmd ==5'h11| frontend_tlb_io_req_bits_cmd ==5'h7| frontend_tlb_io_req_bits_cmd ==5'h4| frontend_tlb_io_req_bits_cmd ==5'h9| frontend_tlb_io_req_bits_cmd ==5'hA| frontend_tlb_io_req_bits_cmd ==5'hB| frontend_tlb_io_req_bits_cmd ==5'h8| frontend_tlb_io_req_bits_cmd ==5'hC| frontend_tlb_io_req_bits_cmd ==5'hD| frontend_tlb_io_req_bits_cmd ==5'hE| frontend_tlb_io_req_bits_cmd ==5'hF; 
    wire frontend_tlb_cmd_write_perms = frontend_tlb_cmd_write | frontend_tlb_io_req_bits_cmd ==5'h5| frontend_tlb_io_req_bits_cmd ==5'h17; 
    wire[6:0] frontend_tlb_ae_array =( frontend_tlb_misaligned  ?  frontend_tlb_eff_array :7'h0)|( frontend_tlb_cmd_lrsc  ? ~ frontend_tlb_lrscAllowed :7'h0); 
    wire[6:0] frontend_tlb_ae_ld_array = frontend_tlb_cmd_read  ?  frontend_tlb_ae_array |~ frontend_tlb_pr_array :7'h0; 
    wire[6:0] frontend_tlb_ae_st_array =( frontend_tlb_cmd_write_perms  ?  frontend_tlb_ae_array |~ frontend_tlb_pw_array :7'h0)|( frontend_tlb_cmd_put_partial  ? ~ frontend_tlb_ppp_array_if_cached :7'h0)|( frontend_tlb_cmd_amo_logical  ? ~ frontend_tlb_pal_array_if_cached :7'h0)|( frontend_tlb_cmd_amo_arithmetic  ? ~ frontend_tlb_paa_array_if_cached :7'h0); 
    wire[6:0] frontend_tlb_must_alloc_array =( frontend_tlb_cmd_put_partial  ? ~ frontend_tlb_ppp_array :7'h0)|( frontend_tlb_cmd_amo_logical  ? ~ frontend_tlb_pal_array :7'h0)|( frontend_tlb_cmd_amo_arithmetic  ? ~ frontend_tlb_paa_array :7'h0)|( frontend_tlb_cmd_lrsc  ? 7'h7F:7'h0); 
    wire[6:0] frontend_tlb_pf_ld_array = frontend_tlb_cmd_read  ? (~( frontend_tlb_cmd_readx  ?  frontend_tlb_x_array : frontend_tlb_r_array )&~ frontend_tlb_ptw_ae_array | frontend_tlb_ptw_pf_array )&~ frontend_tlb_ptw_gf_array :7'h0; 
    wire[6:0] frontend_tlb_pf_st_array = frontend_tlb_cmd_write_perms  ? (~ frontend_tlb_w_array &~ frontend_tlb_ptw_ae_array | frontend_tlb_ptw_pf_array )&~ frontend_tlb_ptw_gf_array :7'h0; 
    wire[6:0] frontend_tlb_pf_inst_array =(~ frontend_tlb_x_array &~ frontend_tlb_ptw_ae_array | frontend_tlb_ptw_pf_array )&~ frontend_tlb_ptw_gf_array ; 
    wire[6:0] frontend_tlb_gf_ld_array = frontend_tlb_priv_v & frontend_tlb_cmd_read  ? (~( frontend_tlb_cmd_readx  ?  frontend_tlb_hx_array : frontend_tlb_hr_array )| frontend_tlb_ptw_gf_array )&~ frontend_tlb_ptw_ae_array :7'h0; 
    wire[6:0] frontend_tlb_gf_st_array = frontend_tlb_priv_v & frontend_tlb_cmd_write_perms  ? (~ frontend_tlb_hw_array | frontend_tlb_ptw_gf_array )&~ frontend_tlb_ptw_ae_array :7'h0; 
    wire[6:0] frontend_tlb_gf_inst_array = frontend_tlb_priv_v  ? (~ frontend_tlb_hx_array | frontend_tlb_ptw_gf_array )&~ frontend_tlb_ptw_ae_array :7'h0; 
    wire[5:0] frontend_tlb_gpa_hits_hit_mask ={1'h0, frontend_tlb_r_gpa_valid & frontend_tlb_r_gpa_vpn == frontend_tlb_vpn  ? 5'h1F:5'h0}|( frontend_tlb_vstage1_en ==1'h0 ? 6'h3F:6'h0); 
    wire[5:0] frontend_tlb_gpa_hits = frontend_tlb_gpa_hits_hit_mask |~( frontend_tlb_gf_inst_array [5:0]); 
    wire frontend_tlb_tlb_hit_if_not_gpa_miss =| frontend_tlb_real_hits ; 
    wire frontend_tlb_tlb_hit =|( frontend_tlb_real_hits & frontend_tlb_gpa_hits ); 
    wire frontend_tlb_tlb_miss = frontend_tlb_vm_enabled & frontend_tlb_vsatp_mode_mismatch ==1'h0& frontend_tlb_tlb_hit ==1'h0; reg[2:0] frontend_tlb_state_reg_1 ; 
    wire frontend_tlb__GEN_34 = frontend_tlb_io_req_valid & frontend_tlb_vm_enabled ; 
    wire frontend_tlb__GEN_35 = frontend_tlb_superpage_hits_0 | frontend_tlb_superpage_hits_1 | frontend_tlb_superpage_hits_2 | frontend_tlb_superpage_hits_3 ; 
    wire[1:0] frontend_tlb_lo ={ frontend_tlb_superpage_hits_1 , frontend_tlb_superpage_hits_0 }; 
    wire[1:0] frontend_tlb_hi ={ frontend_tlb_superpage_hits_3 , frontend_tlb_superpage_hits_2 }; 
    wire[3:0] frontend_tlb__GEN_36 ={ frontend_tlb_hi , frontend_tlb_lo }; 
    wire[1:0] frontend_tlb_hi_1 = frontend_tlb__GEN_36 [3:2]; 
    wire[1:0] frontend_tlb_lo_1 = frontend_tlb__GEN_36 [1:0]; 
    wire[1:0] frontend_tlb__GEN_37 = frontend_tlb_hi_1 | frontend_tlb_lo_1 ; 
    wire[1:0] frontend_tlb_state_reg_touch_way_sized ={| frontend_tlb_hi_1 , frontend_tlb__GEN_37 [1]}; 
    wire frontend_tlb_state_reg_set_left_older = frontend_tlb_state_reg_touch_way_sized [1]==1'h0; 
    wire frontend_tlb_state_reg_left_subtree_state = frontend_tlb_state_reg_1 [1]; 
    wire frontend_tlb_state_reg_right_subtree_state = frontend_tlb_state_reg_1 [0]; 
    wire[1:0] frontend_tlb_state_reg_hi ={ frontend_tlb_state_reg_set_left_older , frontend_tlb_state_reg_set_left_older  ?  frontend_tlb_state_reg_left_subtree_state : frontend_tlb_state_reg_touch_way_sized [0]==1'h0}; 
    wire[2:0] frontend_tlb__GEN_38 ={ frontend_tlb_state_reg_hi , frontend_tlb_state_reg_set_left_older  ?  frontend_tlb_state_reg_touch_way_sized [0]==1'h0: frontend_tlb_state_reg_right_subtree_state }; 
    wire[2:0] frontend_tlb__real_hits_2to0 = frontend_tlb_real_hits [2:0]; 
    wire frontend_tlb_multipleHits_leftOne = frontend_tlb__real_hits_2to0 [0]; 
    wire[1:0] frontend_tlb__real_hits_2to0_2to1 = frontend_tlb__real_hits_2to0 [2:1]; 
    wire frontend_tlb_multipleHits_leftOne_1 = frontend_tlb__real_hits_2to0_2to1 [0]; 
    wire frontend_tlb_multipleHits_rightOne = frontend_tlb__real_hits_2to0_2to1 [1]; 
    wire frontend_tlb_multipleHits_rightOne_1 = frontend_tlb_multipleHits_leftOne_1 | frontend_tlb_multipleHits_rightOne ; 
    wire frontend_tlb_multipleHits_rightTwo = frontend_tlb_multipleHits_leftOne_1 & frontend_tlb_multipleHits_rightOne |1'h0; 
    wire frontend_tlb_multipleHits_leftOne_2 = frontend_tlb_multipleHits_leftOne | frontend_tlb_multipleHits_rightOne_1 ; 
    wire frontend_tlb_multipleHits_leftTwo = frontend_tlb_multipleHits_rightTwo |1'h0| frontend_tlb_multipleHits_leftOne & frontend_tlb_multipleHits_rightOne_1 ; 
    wire[2:0] frontend_tlb__real_hits_5to3 = frontend_tlb_real_hits [5:3]; 
    wire frontend_tlb_multipleHits_leftOne_3 = frontend_tlb__real_hits_5to3 [0]; 
    wire[1:0] frontend_tlb__real_hits_5to3_2to1 = frontend_tlb__real_hits_5to3 [2:1]; 
    wire frontend_tlb_multipleHits_leftOne_4 = frontend_tlb__real_hits_5to3_2to1 [0]; 
    wire frontend_tlb_multipleHits_rightOne_2 = frontend_tlb__real_hits_5to3_2to1 [1]; 
    wire frontend_tlb_multipleHits_rightOne_3 = frontend_tlb_multipleHits_leftOne_4 | frontend_tlb_multipleHits_rightOne_2 ; 
    wire frontend_tlb_multipleHits_rightTwo_1 = frontend_tlb_multipleHits_leftOne_4 & frontend_tlb_multipleHits_rightOne_2 |1'h0; 
    wire frontend_tlb_multipleHits_rightOne_4 = frontend_tlb_multipleHits_leftOne_3 | frontend_tlb_multipleHits_rightOne_3 ; 
    wire frontend_tlb_multipleHits_rightTwo_2 = frontend_tlb_multipleHits_rightTwo_1 |1'h0| frontend_tlb_multipleHits_leftOne_3 & frontend_tlb_multipleHits_rightOne_3 ; 
    wire frontend_tlb_multipleHits = frontend_tlb_multipleHits_leftTwo | frontend_tlb_multipleHits_rightTwo_2 | frontend_tlb_multipleHits_leftOne_2 & frontend_tlb_multipleHits_rightOne_4 ; 
    wire frontend_tlb__io_resp_gpa_is_pte_output = frontend_tlb_vstage1_en & frontend_tlb_r_gpa_is_pte ; 
    wire[21:0] frontend_tlb_io_resp_gpa_page = frontend_tlb_vstage1_en ==1'h0 ? {1'h0, frontend_tlb_vpn }:{1'h0, frontend_tlb_r_gpa [32:12]}; 
    wire[11:0] frontend_tlb_io_resp_gpa_offset = frontend_tlb__io_resp_gpa_is_pte_output  ?  frontend_tlb_r_gpa [11:0]: frontend_tlb_io_req_bits_vaddr [11:0]; 
  always @( posedge  frontend_tlb_clock )
         begin 
             if ( frontend_tlb_do_refill )
                 begin 
                     if ( frontend_tlb__GEN_1 )
                         begin  
                             frontend_tlb_special_entry_level  <= frontend_tlb_io_ptw_resp_bits_level ; 
                             frontend_tlb_special_entry_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                             frontend_tlb_special_entry_tag_v  <= frontend_tlb_refill_v ; 
                             frontend_tlb_special_entry_data_0  <= frontend_tlb__GEN_2 ; 
                             frontend_tlb_special_entry_valid_0  <=1'h1;
                         end 
                      else 
                         if ( frontend_tlb__GEN_4 )
                             begin 
                                 if ( frontend_tlb__GEN_6 )
                                     begin  
                                         frontend_tlb_superpage_entries_0_level  <= frontend_tlb__GEN_7 ; 
                                         frontend_tlb_superpage_entries_0_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                                         frontend_tlb_superpage_entries_0_tag_v  <= frontend_tlb_refill_v ; 
                                         frontend_tlb_superpage_entries_0_data_0  <= frontend_tlb__GEN_8 ; 
                                         frontend_tlb_superpage_entries_0_valid_0  <= frontend_tlb__GEN_9 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_10 )
                                     begin  
                                         frontend_tlb_superpage_entries_1_level  <= frontend_tlb__GEN_11 ; 
                                         frontend_tlb_superpage_entries_1_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                                         frontend_tlb_superpage_entries_1_tag_v  <= frontend_tlb_refill_v ; 
                                         frontend_tlb_superpage_entries_1_data_0  <= frontend_tlb__GEN_12 ; 
                                         frontend_tlb_superpage_entries_1_valid_0  <= frontend_tlb__GEN_13 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_14 )
                                     begin  
                                         frontend_tlb_superpage_entries_2_level  <= frontend_tlb__GEN_15 ; 
                                         frontend_tlb_superpage_entries_2_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                                         frontend_tlb_superpage_entries_2_tag_v  <= frontend_tlb_refill_v ; 
                                         frontend_tlb_superpage_entries_2_data_0  <= frontend_tlb__GEN_16 ; 
                                         frontend_tlb_superpage_entries_2_valid_0  <= frontend_tlb__GEN_17 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_18 )
                                     begin  
                                         frontend_tlb_superpage_entries_3_level  <= frontend_tlb__GEN_19 ; 
                                         frontend_tlb_superpage_entries_3_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                                         frontend_tlb_superpage_entries_3_tag_v  <= frontend_tlb_refill_v ; 
                                         frontend_tlb_superpage_entries_3_data_0  <= frontend_tlb__GEN_20 ; 
                                         frontend_tlb_superpage_entries_3_valid_0  <= frontend_tlb__GEN_21 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin  
                                 frontend_tlb_sectored_entries_0_0_level  <=2'h0; 
                                 frontend_tlb_sectored_entries_0_0_tag_vpn  <= frontend_tlb_r_refill_tag ; 
                                 frontend_tlb_sectored_entries_0_0_tag_v  <= frontend_tlb_refill_v ;
                                 if ( frontend_tlb__GEN_29 ) 
                                     frontend_tlb_sectored_entries_0_0_data_0  <= frontend_tlb__GEN_28 ;
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_30 ) 
                                     frontend_tlb_sectored_entries_0_0_data_1  <= frontend_tlb__GEN_28 ;
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_31 ) 
                                     frontend_tlb_sectored_entries_0_0_data_2  <= frontend_tlb__GEN_28 ;
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb__GEN_32 ) 
                                     frontend_tlb_sectored_entries_0_0_data_3  <= frontend_tlb__GEN_28 ;
                                  else 
                                     begin 
                                     end 
                                 if ( frontend_tlb_invalidate_refill )
                                     begin  
                                         frontend_tlb_sectored_entries_0_0_valid_0  <=1'h0; 
                                         frontend_tlb_sectored_entries_0_0_valid_1  <=1'h0; 
                                         frontend_tlb_sectored_entries_0_0_valid_2  <=1'h0; 
                                         frontend_tlb_sectored_entries_0_0_valid_3  <=1'h0;
                                     end 
                                  else 
                                     begin 
                                         if ( frontend_tlb__GEN_24 ) 
                                             frontend_tlb_sectored_entries_0_0_valid_0  <=1'h1;
                                          else 
                                             if ( frontend_tlb__GEN_23 ) 
                                                 frontend_tlb_sectored_entries_0_0_valid_0  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( frontend_tlb__GEN_25 ) 
                                             frontend_tlb_sectored_entries_0_0_valid_1  <=1'h1;
                                          else 
                                             if ( frontend_tlb__GEN_23 ) 
                                                 frontend_tlb_sectored_entries_0_0_valid_1  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( frontend_tlb__GEN_26 ) 
                                             frontend_tlb_sectored_entries_0_0_valid_2  <=1'h1;
                                          else 
                                             if ( frontend_tlb__GEN_23 ) 
                                                 frontend_tlb_sectored_entries_0_0_valid_2  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         if ( frontend_tlb__GEN_27 ) 
                                             frontend_tlb_sectored_entries_0_0_valid_3  <=1'h1;
                                          else 
                                             if ( frontend_tlb__GEN_23 ) 
                                                 frontend_tlb_sectored_entries_0_0_valid_3  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                     end 
                             end  
                     frontend_tlb_r_gpa_valid  <= frontend_tlb_io_ptw_resp_bits_gpa_valid ; 
                     frontend_tlb_r_gpa  <= frontend_tlb_io_ptw_resp_bits_gpa_bits ; 
                     frontend_tlb_r_gpa_is_pte  <= frontend_tlb_io_ptw_resp_bits_gpa_is_pte ;
                 end 
              else 
                 begin 
                 end 
         end
  always @( posedge  frontend_tlb_clock )
         begin 
             if ( frontend_tlb_reset )
                 begin  
                     frontend_tlb_state  <=2'h0; 
                     frontend_tlb_v_entries_use_stage1  <=1'h0; 
                     frontend_tlb_state_reg_1  <=3'h0;
                 end 
              else 
                 if ( frontend_tlb__GEN_34 )
                     begin 
                         if ( frontend_tlb__GEN_35 ) 
                             frontend_tlb_state_reg_1  <= frontend_tlb__GEN_38 ;
                          else 
                             begin 
                             end 
                     end 
                  else 
                     begin 
                     end 
         end
  assign  frontend_tlb_io_req_ready = frontend_tlb_state ==2'h0; 
  assign  frontend_tlb_io_resp_miss = frontend_tlb_do_refill | frontend_tlb_vsatp_mode_mismatch | frontend_tlb_tlb_miss | frontend_tlb_multipleHits ; 
  assign  frontend_tlb_io_resp_paddr ={ frontend_tlb_ppn , frontend_tlb_io_req_bits_vaddr [11:0]}; 
  assign  frontend_tlb_io_resp_gpa ={ frontend_tlb_io_resp_gpa_page , frontend_tlb_io_resp_gpa_offset }; 
  assign  frontend_tlb_io_resp_gpa_is_pte = frontend_tlb__io_resp_gpa_is_pte_output ; 
  assign  frontend_tlb_io_resp_pf_ld =(|( frontend_tlb_pf_ld_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_pf_st =(|( frontend_tlb_pf_st_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_pf_inst =(|( frontend_tlb_pf_inst_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_gf_ld =(|( frontend_tlb_gf_ld_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_gf_st =(|( frontend_tlb_gf_st_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_gf_inst =(|( frontend_tlb_gf_inst_array & frontend_tlb_hits ))|1'h0; 
  assign  frontend_tlb_io_resp_ae_ld =|( frontend_tlb_ae_ld_array & frontend_tlb_hits ); 
  assign  frontend_tlb_io_resp_ae_st =|( frontend_tlb_ae_st_array & frontend_tlb_hits ); 
  assign  frontend_tlb_io_resp_ae_inst =|(~ frontend_tlb_px_array & frontend_tlb_hits ); 
  assign  frontend_tlb_io_resp_ma_ld = frontend_tlb_misaligned & frontend_tlb_cmd_read ; 
  assign  frontend_tlb_io_resp_ma_st = frontend_tlb_misaligned & frontend_tlb_cmd_write ; 
  assign  frontend_tlb_io_resp_ma_inst =1'h0; 
  assign  frontend_tlb_io_resp_cacheable =|( frontend_tlb_c_array & frontend_tlb_hits ); 
  assign  frontend_tlb_io_resp_must_alloc =|( frontend_tlb_must_alloc_array & frontend_tlb_hits ); 
  assign  frontend_tlb_io_resp_prefetchable =1'h0; 
  assign  frontend_tlb_io_ptw_req_valid = frontend_tlb_state ==2'h1; 
  assign  frontend_tlb_io_ptw_req_bits_valid = frontend_tlb_io_kill ==1'h0; 
  assign  frontend_tlb_io_ptw_req_bits_bits_addr = frontend_tlb_r_refill_tag ; 
  assign  frontend_tlb_io_ptw_req_bits_bits_need_gpa = frontend_tlb_r_need_gpa ; 
  assign  frontend_tlb_io_ptw_req_bits_bits_vstage1 = frontend_tlb_r_vstage1_en ; 
  assign  frontend_tlb_io_ptw_req_bits_bits_stage2 = frontend_tlb_r_stage2_en ; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_0_stall =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_0_set =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_0_sdata =64'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_1_stall =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_1_set =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_1_sdata =64'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_2_stall =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_2_set =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_2_sdata =64'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_3_stall =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_3_set =1'h0; 
  assign  frontend_tlb_io_ptw_customCSRs_csrs_3_sdata =64'h0;
    assign frontend_tlb_clock = frontend_clock;
    assign frontend_tlb_reset = frontend_reset;
    assign frontend__tlb_io_req_ready = frontend_tlb_io_req_ready;
    assign frontend_tlb_io_req_valid = frontend__GEN_7;
    assign frontend_tlb_io_req_bits_vaddr = frontend_s1_pc;
    assign frontend_tlb_io_req_bits_passthrough = 1'h0;
    assign frontend_tlb_io_req_bits_size = 2'h2;
    assign frontend_tlb_io_req_bits_cmd = 5'h0;
    assign frontend_tlb_io_req_bits_prv = frontend_io_ptw_status_prv;
    assign frontend_tlb_io_req_bits_v = frontend_io_ptw_status_v;
    assign frontend__tlb_io_resp_miss = frontend_tlb_io_resp_miss;
    assign frontend__tlb_io_resp_paddr = frontend_tlb_io_resp_paddr;
    assign frontend__tlb_io_resp_gpa = frontend_tlb_io_resp_gpa;
    assign frontend__tlb_io_resp_gpa_is_pte = frontend_tlb_io_resp_gpa_is_pte;
    assign frontend__tlb_io_resp_pf_ld = frontend_tlb_io_resp_pf_ld;
    assign frontend__tlb_io_resp_pf_st = frontend_tlb_io_resp_pf_st;
    assign frontend__tlb_io_resp_pf_inst = frontend_tlb_io_resp_pf_inst;
    assign frontend__tlb_io_resp_gf_ld = frontend_tlb_io_resp_gf_ld;
    assign frontend__tlb_io_resp_gf_st = frontend_tlb_io_resp_gf_st;
    assign frontend__tlb_io_resp_gf_inst = frontend_tlb_io_resp_gf_inst;
    assign frontend__tlb_io_resp_ae_ld = frontend_tlb_io_resp_ae_ld;
    assign frontend__tlb_io_resp_ae_st = frontend_tlb_io_resp_ae_st;
    assign frontend__tlb_io_resp_ae_inst = frontend_tlb_io_resp_ae_inst;
    assign frontend__tlb_io_resp_ma_ld = frontend_tlb_io_resp_ma_ld;
    assign frontend__tlb_io_resp_ma_st = frontend_tlb_io_resp_ma_st;
    assign frontend__tlb_io_resp_ma_inst = frontend_tlb_io_resp_ma_inst;
    assign frontend__tlb_io_resp_cacheable = frontend_tlb_io_resp_cacheable;
    assign frontend__tlb_io_resp_must_alloc = frontend_tlb_io_resp_must_alloc;
    assign frontend__tlb_io_resp_prefetchable = frontend_tlb_io_resp_prefetchable;
    assign frontend_tlb_io_sfence_valid = frontend_io_cpu_sfence_valid;
    assign frontend_tlb_io_sfence_bits_rs1 = frontend_io_cpu_sfence_bits_rs1;
    assign frontend_tlb_io_sfence_bits_rs2 = frontend_io_cpu_sfence_bits_rs2;
    assign frontend_tlb_io_sfence_bits_addr = frontend_io_cpu_sfence_bits_addr;
    assign frontend_tlb_io_sfence_bits_asid = frontend_io_cpu_sfence_bits_asid;
    assign frontend_tlb_io_sfence_bits_hv = frontend_io_cpu_sfence_bits_hv;
    assign frontend_tlb_io_sfence_bits_hg = frontend_io_cpu_sfence_bits_hg;
    assign frontend_tlb_io_ptw_req_ready = frontend_io_ptw_req_ready;
    assign frontend__io_ptw_req_valid_output = frontend_tlb_io_ptw_req_valid;
    assign frontend_io_ptw_req_bits_valid = frontend_tlb_io_ptw_req_bits_valid;
    assign frontend_io_ptw_req_bits_bits_addr = frontend_tlb_io_ptw_req_bits_bits_addr;
    assign frontend_io_ptw_req_bits_bits_need_gpa = frontend_tlb_io_ptw_req_bits_bits_need_gpa;
    assign frontend_io_ptw_req_bits_bits_vstage1 = frontend_tlb_io_ptw_req_bits_bits_vstage1;
    assign frontend_io_ptw_req_bits_bits_stage2 = frontend_tlb_io_ptw_req_bits_bits_stage2;
    assign frontend_tlb_io_ptw_resp_valid = frontend_io_ptw_resp_valid;
    assign frontend_tlb_io_ptw_resp_bits_ae_ptw = frontend_io_ptw_resp_bits_ae_ptw;
    assign frontend_tlb_io_ptw_resp_bits_ae_final = frontend_io_ptw_resp_bits_ae_final;
    assign frontend_tlb_io_ptw_resp_bits_pf = frontend_io_ptw_resp_bits_pf;
    assign frontend_tlb_io_ptw_resp_bits_gf = frontend_io_ptw_resp_bits_gf;
    assign frontend_tlb_io_ptw_resp_bits_hr = frontend_io_ptw_resp_bits_hr;
    assign frontend_tlb_io_ptw_resp_bits_hw = frontend_io_ptw_resp_bits_hw;
    assign frontend_tlb_io_ptw_resp_bits_hx = frontend_io_ptw_resp_bits_hx;
    assign frontend_tlb_io_ptw_resp_bits_pte_reserved_for_future = frontend_io_ptw_resp_bits_pte_reserved_for_future;
    assign frontend_tlb_io_ptw_resp_bits_pte_ppn = frontend_io_ptw_resp_bits_pte_ppn;
    assign frontend_tlb_io_ptw_resp_bits_pte_reserved_for_software = frontend_io_ptw_resp_bits_pte_reserved_for_software;
    assign frontend_tlb_io_ptw_resp_bits_pte_d = frontend_io_ptw_resp_bits_pte_d;
    assign frontend_tlb_io_ptw_resp_bits_pte_a = frontend_io_ptw_resp_bits_pte_a;
    assign frontend_tlb_io_ptw_resp_bits_pte_g = frontend_io_ptw_resp_bits_pte_g;
    assign frontend_tlb_io_ptw_resp_bits_pte_u = frontend_io_ptw_resp_bits_pte_u;
    assign frontend_tlb_io_ptw_resp_bits_pte_x = frontend_io_ptw_resp_bits_pte_x;
    assign frontend_tlb_io_ptw_resp_bits_pte_w = frontend_io_ptw_resp_bits_pte_w;
    assign frontend_tlb_io_ptw_resp_bits_pte_r = frontend_io_ptw_resp_bits_pte_r;
    assign frontend_tlb_io_ptw_resp_bits_pte_v = frontend_io_ptw_resp_bits_pte_v;
    assign frontend_tlb_io_ptw_resp_bits_level = frontend_io_ptw_resp_bits_level;
    assign frontend_tlb_io_ptw_resp_bits_fragmented_superpage = frontend_io_ptw_resp_bits_fragmented_superpage;
    assign frontend_tlb_io_ptw_resp_bits_homogeneous = frontend_io_ptw_resp_bits_homogeneous;
    assign frontend_tlb_io_ptw_resp_bits_gpa_valid = frontend_io_ptw_resp_bits_gpa_valid;
    assign frontend_tlb_io_ptw_resp_bits_gpa_bits = frontend_io_ptw_resp_bits_gpa_bits;
    assign frontend_tlb_io_ptw_resp_bits_gpa_is_pte = frontend_io_ptw_resp_bits_gpa_is_pte;
    assign frontend_tlb_io_ptw_ptbr_mode = frontend_io_ptw_ptbr_mode;
    assign frontend_tlb_io_ptw_ptbr_asid = frontend_io_ptw_ptbr_asid;
    assign frontend_tlb_io_ptw_ptbr_ppn = frontend_io_ptw_ptbr_ppn;
    assign frontend_tlb_io_ptw_hgatp_mode = frontend_io_ptw_hgatp_mode;
    assign frontend_tlb_io_ptw_hgatp_asid = frontend_io_ptw_hgatp_asid;
    assign frontend_tlb_io_ptw_hgatp_ppn = frontend_io_ptw_hgatp_ppn;
    assign frontend_tlb_io_ptw_vsatp_mode = frontend_io_ptw_vsatp_mode;
    assign frontend_tlb_io_ptw_vsatp_asid = frontend_io_ptw_vsatp_asid;
    assign frontend_tlb_io_ptw_vsatp_ppn = frontend_io_ptw_vsatp_ppn;
    assign frontend_tlb_io_ptw_status_debug = frontend_io_ptw_status_debug;
    assign frontend_tlb_io_ptw_status_cease = frontend_io_ptw_status_cease;
    assign frontend_tlb_io_ptw_status_wfi = frontend_io_ptw_status_wfi;
    assign frontend_tlb_io_ptw_status_isa = frontend_io_ptw_status_isa;
    assign frontend_tlb_io_ptw_status_dprv = frontend_io_ptw_status_dprv;
    assign frontend_tlb_io_ptw_status_dv = frontend_io_ptw_status_dv;
    assign frontend_tlb_io_ptw_status_prv = frontend_io_ptw_status_prv;
    assign frontend_tlb_io_ptw_status_v = frontend_io_ptw_status_v;
    assign frontend_tlb_io_ptw_status_sd = frontend_io_ptw_status_sd;
    assign frontend_tlb_io_ptw_status_zero2 = frontend_io_ptw_status_zero2;
    assign frontend_tlb_io_ptw_status_mpv = frontend_io_ptw_status_mpv;
    assign frontend_tlb_io_ptw_status_gva = frontend_io_ptw_status_gva;
    assign frontend_tlb_io_ptw_status_mbe = frontend_io_ptw_status_mbe;
    assign frontend_tlb_io_ptw_status_sbe = frontend_io_ptw_status_sbe;
    assign frontend_tlb_io_ptw_status_sxl = frontend_io_ptw_status_sxl;
    assign frontend_tlb_io_ptw_status_uxl = frontend_io_ptw_status_uxl;
    assign frontend_tlb_io_ptw_status_sd_rv32 = frontend_io_ptw_status_sd_rv32;
    assign frontend_tlb_io_ptw_status_zero1 = frontend_io_ptw_status_zero1;
    assign frontend_tlb_io_ptw_status_tsr = frontend_io_ptw_status_tsr;
    assign frontend_tlb_io_ptw_status_tw = frontend_io_ptw_status_tw;
    assign frontend_tlb_io_ptw_status_tvm = frontend_io_ptw_status_tvm;
    assign frontend_tlb_io_ptw_status_mxr = frontend_io_ptw_status_mxr;
    assign frontend_tlb_io_ptw_status_sum = frontend_io_ptw_status_sum;
    assign frontend_tlb_io_ptw_status_mprv = frontend_io_ptw_status_mprv;
    assign frontend_tlb_io_ptw_status_xs = frontend_io_ptw_status_xs;
    assign frontend_tlb_io_ptw_status_fs = frontend_io_ptw_status_fs;
    assign frontend_tlb_io_ptw_status_mpp = frontend_io_ptw_status_mpp;
    assign frontend_tlb_io_ptw_status_vs = frontend_io_ptw_status_vs;
    assign frontend_tlb_io_ptw_status_spp = frontend_io_ptw_status_spp;
    assign frontend_tlb_io_ptw_status_mpie = frontend_io_ptw_status_mpie;
    assign frontend_tlb_io_ptw_status_ube = frontend_io_ptw_status_ube;
    assign frontend_tlb_io_ptw_status_spie = frontend_io_ptw_status_spie;
    assign frontend_tlb_io_ptw_status_upie = frontend_io_ptw_status_upie;
    assign frontend_tlb_io_ptw_status_mie = frontend_io_ptw_status_mie;
    assign frontend_tlb_io_ptw_status_hie = frontend_io_ptw_status_hie;
    assign frontend_tlb_io_ptw_status_sie = frontend_io_ptw_status_sie;
    assign frontend_tlb_io_ptw_status_uie = frontend_io_ptw_status_uie;
    assign frontend_tlb_io_ptw_hstatus_zero6 = frontend_io_ptw_hstatus_zero6;
    assign frontend_tlb_io_ptw_hstatus_vsxl = frontend_io_ptw_hstatus_vsxl;
    assign frontend_tlb_io_ptw_hstatus_zero5 = frontend_io_ptw_hstatus_zero5;
    assign frontend_tlb_io_ptw_hstatus_vtsr = frontend_io_ptw_hstatus_vtsr;
    assign frontend_tlb_io_ptw_hstatus_vtw = frontend_io_ptw_hstatus_vtw;
    assign frontend_tlb_io_ptw_hstatus_vtvm = frontend_io_ptw_hstatus_vtvm;
    assign frontend_tlb_io_ptw_hstatus_zero3 = frontend_io_ptw_hstatus_zero3;
    assign frontend_tlb_io_ptw_hstatus_vgein = frontend_io_ptw_hstatus_vgein;
    assign frontend_tlb_io_ptw_hstatus_zero2 = frontend_io_ptw_hstatus_zero2;
    assign frontend_tlb_io_ptw_hstatus_hu = frontend_io_ptw_hstatus_hu;
    assign frontend_tlb_io_ptw_hstatus_spvp = frontend_io_ptw_hstatus_spvp;
    assign frontend_tlb_io_ptw_hstatus_spv = frontend_io_ptw_hstatus_spv;
    assign frontend_tlb_io_ptw_hstatus_gva = frontend_io_ptw_hstatus_gva;
    assign frontend_tlb_io_ptw_hstatus_vsbe = frontend_io_ptw_hstatus_vsbe;
    assign frontend_tlb_io_ptw_hstatus_zero1 = frontend_io_ptw_hstatus_zero1;
    assign frontend_tlb_io_ptw_gstatus_debug = frontend_io_ptw_gstatus_debug;
    assign frontend_tlb_io_ptw_gstatus_cease = frontend_io_ptw_gstatus_cease;
    assign frontend_tlb_io_ptw_gstatus_wfi = frontend_io_ptw_gstatus_wfi;
    assign frontend_tlb_io_ptw_gstatus_isa = frontend_io_ptw_gstatus_isa;
    assign frontend_tlb_io_ptw_gstatus_dprv = frontend_io_ptw_gstatus_dprv;
    assign frontend_tlb_io_ptw_gstatus_dv = frontend_io_ptw_gstatus_dv;
    assign frontend_tlb_io_ptw_gstatus_prv = frontend_io_ptw_gstatus_prv;
    assign frontend_tlb_io_ptw_gstatus_v = frontend_io_ptw_gstatus_v;
    assign frontend_tlb_io_ptw_gstatus_sd = frontend_io_ptw_gstatus_sd;
    assign frontend_tlb_io_ptw_gstatus_zero2 = frontend_io_ptw_gstatus_zero2;
    assign frontend_tlb_io_ptw_gstatus_mpv = frontend_io_ptw_gstatus_mpv;
    assign frontend_tlb_io_ptw_gstatus_gva = frontend_io_ptw_gstatus_gva;
    assign frontend_tlb_io_ptw_gstatus_mbe = frontend_io_ptw_gstatus_mbe;
    assign frontend_tlb_io_ptw_gstatus_sbe = frontend_io_ptw_gstatus_sbe;
    assign frontend_tlb_io_ptw_gstatus_sxl = frontend_io_ptw_gstatus_sxl;
    assign frontend_tlb_io_ptw_gstatus_uxl = frontend_io_ptw_gstatus_uxl;
    assign frontend_tlb_io_ptw_gstatus_sd_rv32 = frontend_io_ptw_gstatus_sd_rv32;
    assign frontend_tlb_io_ptw_gstatus_zero1 = frontend_io_ptw_gstatus_zero1;
    assign frontend_tlb_io_ptw_gstatus_tsr = frontend_io_ptw_gstatus_tsr;
    assign frontend_tlb_io_ptw_gstatus_tw = frontend_io_ptw_gstatus_tw;
    assign frontend_tlb_io_ptw_gstatus_tvm = frontend_io_ptw_gstatus_tvm;
    assign frontend_tlb_io_ptw_gstatus_mxr = frontend_io_ptw_gstatus_mxr;
    assign frontend_tlb_io_ptw_gstatus_sum = frontend_io_ptw_gstatus_sum;
    assign frontend_tlb_io_ptw_gstatus_mprv = frontend_io_ptw_gstatus_mprv;
    assign frontend_tlb_io_ptw_gstatus_xs = frontend_io_ptw_gstatus_xs;
    assign frontend_tlb_io_ptw_gstatus_fs = frontend_io_ptw_gstatus_fs;
    assign frontend_tlb_io_ptw_gstatus_mpp = frontend_io_ptw_gstatus_mpp;
    assign frontend_tlb_io_ptw_gstatus_vs = frontend_io_ptw_gstatus_vs;
    assign frontend_tlb_io_ptw_gstatus_spp = frontend_io_ptw_gstatus_spp;
    assign frontend_tlb_io_ptw_gstatus_mpie = frontend_io_ptw_gstatus_mpie;
    assign frontend_tlb_io_ptw_gstatus_ube = frontend_io_ptw_gstatus_ube;
    assign frontend_tlb_io_ptw_gstatus_spie = frontend_io_ptw_gstatus_spie;
    assign frontend_tlb_io_ptw_gstatus_upie = frontend_io_ptw_gstatus_upie;
    assign frontend_tlb_io_ptw_gstatus_mie = frontend_io_ptw_gstatus_mie;
    assign frontend_tlb_io_ptw_gstatus_hie = frontend_io_ptw_gstatus_hie;
    assign frontend_tlb_io_ptw_gstatus_sie = frontend_io_ptw_gstatus_sie;
    assign frontend_tlb_io_ptw_gstatus_uie = frontend_io_ptw_gstatus_uie;
    assign frontend_tlb_io_ptw_pmp_0_cfg_l = frontend_io_ptw_pmp_0_cfg_l;
    assign frontend_tlb_io_ptw_pmp_0_cfg_res = frontend_io_ptw_pmp_0_cfg_res;
    assign frontend_tlb_io_ptw_pmp_0_cfg_a = frontend_io_ptw_pmp_0_cfg_a;
    assign frontend_tlb_io_ptw_pmp_0_cfg_x = frontend_io_ptw_pmp_0_cfg_x;
    assign frontend_tlb_io_ptw_pmp_0_cfg_w = frontend_io_ptw_pmp_0_cfg_w;
    assign frontend_tlb_io_ptw_pmp_0_cfg_r = frontend_io_ptw_pmp_0_cfg_r;
    assign frontend_tlb_io_ptw_pmp_0_addr = frontend_io_ptw_pmp_0_addr;
    assign frontend_tlb_io_ptw_pmp_0_mask = frontend_io_ptw_pmp_0_mask;
    assign frontend_tlb_io_ptw_pmp_1_cfg_l = frontend_io_ptw_pmp_1_cfg_l;
    assign frontend_tlb_io_ptw_pmp_1_cfg_res = frontend_io_ptw_pmp_1_cfg_res;
    assign frontend_tlb_io_ptw_pmp_1_cfg_a = frontend_io_ptw_pmp_1_cfg_a;
    assign frontend_tlb_io_ptw_pmp_1_cfg_x = frontend_io_ptw_pmp_1_cfg_x;
    assign frontend_tlb_io_ptw_pmp_1_cfg_w = frontend_io_ptw_pmp_1_cfg_w;
    assign frontend_tlb_io_ptw_pmp_1_cfg_r = frontend_io_ptw_pmp_1_cfg_r;
    assign frontend_tlb_io_ptw_pmp_1_addr = frontend_io_ptw_pmp_1_addr;
    assign frontend_tlb_io_ptw_pmp_1_mask = frontend_io_ptw_pmp_1_mask;
    assign frontend_tlb_io_ptw_pmp_2_cfg_l = frontend_io_ptw_pmp_2_cfg_l;
    assign frontend_tlb_io_ptw_pmp_2_cfg_res = frontend_io_ptw_pmp_2_cfg_res;
    assign frontend_tlb_io_ptw_pmp_2_cfg_a = frontend_io_ptw_pmp_2_cfg_a;
    assign frontend_tlb_io_ptw_pmp_2_cfg_x = frontend_io_ptw_pmp_2_cfg_x;
    assign frontend_tlb_io_ptw_pmp_2_cfg_w = frontend_io_ptw_pmp_2_cfg_w;
    assign frontend_tlb_io_ptw_pmp_2_cfg_r = frontend_io_ptw_pmp_2_cfg_r;
    assign frontend_tlb_io_ptw_pmp_2_addr = frontend_io_ptw_pmp_2_addr;
    assign frontend_tlb_io_ptw_pmp_2_mask = frontend_io_ptw_pmp_2_mask;
    assign frontend_tlb_io_ptw_pmp_3_cfg_l = frontend_io_ptw_pmp_3_cfg_l;
    assign frontend_tlb_io_ptw_pmp_3_cfg_res = frontend_io_ptw_pmp_3_cfg_res;
    assign frontend_tlb_io_ptw_pmp_3_cfg_a = frontend_io_ptw_pmp_3_cfg_a;
    assign frontend_tlb_io_ptw_pmp_3_cfg_x = frontend_io_ptw_pmp_3_cfg_x;
    assign frontend_tlb_io_ptw_pmp_3_cfg_w = frontend_io_ptw_pmp_3_cfg_w;
    assign frontend_tlb_io_ptw_pmp_3_cfg_r = frontend_io_ptw_pmp_3_cfg_r;
    assign frontend_tlb_io_ptw_pmp_3_addr = frontend_io_ptw_pmp_3_addr;
    assign frontend_tlb_io_ptw_pmp_3_mask = frontend_io_ptw_pmp_3_mask;
    assign frontend_tlb_io_ptw_pmp_4_cfg_l = frontend_io_ptw_pmp_4_cfg_l;
    assign frontend_tlb_io_ptw_pmp_4_cfg_res = frontend_io_ptw_pmp_4_cfg_res;
    assign frontend_tlb_io_ptw_pmp_4_cfg_a = frontend_io_ptw_pmp_4_cfg_a;
    assign frontend_tlb_io_ptw_pmp_4_cfg_x = frontend_io_ptw_pmp_4_cfg_x;
    assign frontend_tlb_io_ptw_pmp_4_cfg_w = frontend_io_ptw_pmp_4_cfg_w;
    assign frontend_tlb_io_ptw_pmp_4_cfg_r = frontend_io_ptw_pmp_4_cfg_r;
    assign frontend_tlb_io_ptw_pmp_4_addr = frontend_io_ptw_pmp_4_addr;
    assign frontend_tlb_io_ptw_pmp_4_mask = frontend_io_ptw_pmp_4_mask;
    assign frontend_tlb_io_ptw_pmp_5_cfg_l = frontend_io_ptw_pmp_5_cfg_l;
    assign frontend_tlb_io_ptw_pmp_5_cfg_res = frontend_io_ptw_pmp_5_cfg_res;
    assign frontend_tlb_io_ptw_pmp_5_cfg_a = frontend_io_ptw_pmp_5_cfg_a;
    assign frontend_tlb_io_ptw_pmp_5_cfg_x = frontend_io_ptw_pmp_5_cfg_x;
    assign frontend_tlb_io_ptw_pmp_5_cfg_w = frontend_io_ptw_pmp_5_cfg_w;
    assign frontend_tlb_io_ptw_pmp_5_cfg_r = frontend_io_ptw_pmp_5_cfg_r;
    assign frontend_tlb_io_ptw_pmp_5_addr = frontend_io_ptw_pmp_5_addr;
    assign frontend_tlb_io_ptw_pmp_5_mask = frontend_io_ptw_pmp_5_mask;
    assign frontend_tlb_io_ptw_pmp_6_cfg_l = frontend_io_ptw_pmp_6_cfg_l;
    assign frontend_tlb_io_ptw_pmp_6_cfg_res = frontend_io_ptw_pmp_6_cfg_res;
    assign frontend_tlb_io_ptw_pmp_6_cfg_a = frontend_io_ptw_pmp_6_cfg_a;
    assign frontend_tlb_io_ptw_pmp_6_cfg_x = frontend_io_ptw_pmp_6_cfg_x;
    assign frontend_tlb_io_ptw_pmp_6_cfg_w = frontend_io_ptw_pmp_6_cfg_w;
    assign frontend_tlb_io_ptw_pmp_6_cfg_r = frontend_io_ptw_pmp_6_cfg_r;
    assign frontend_tlb_io_ptw_pmp_6_addr = frontend_io_ptw_pmp_6_addr;
    assign frontend_tlb_io_ptw_pmp_6_mask = frontend_io_ptw_pmp_6_mask;
    assign frontend_tlb_io_ptw_pmp_7_cfg_l = frontend_io_ptw_pmp_7_cfg_l;
    assign frontend_tlb_io_ptw_pmp_7_cfg_res = frontend_io_ptw_pmp_7_cfg_res;
    assign frontend_tlb_io_ptw_pmp_7_cfg_a = frontend_io_ptw_pmp_7_cfg_a;
    assign frontend_tlb_io_ptw_pmp_7_cfg_x = frontend_io_ptw_pmp_7_cfg_x;
    assign frontend_tlb_io_ptw_pmp_7_cfg_w = frontend_io_ptw_pmp_7_cfg_w;
    assign frontend_tlb_io_ptw_pmp_7_cfg_r = frontend_io_ptw_pmp_7_cfg_r;
    assign frontend_tlb_io_ptw_pmp_7_addr = frontend_io_ptw_pmp_7_addr;
    assign frontend_tlb_io_ptw_pmp_7_mask = frontend_io_ptw_pmp_7_mask;
    assign frontend_tlb_io_ptw_customCSRs_csrs_0_ren = frontend_io_ptw_customCSRs_csrs_0_ren;
    assign frontend_tlb_io_ptw_customCSRs_csrs_0_wen = frontend_io_ptw_customCSRs_csrs_0_wen;
    assign frontend_tlb_io_ptw_customCSRs_csrs_0_wdata = frontend_io_ptw_customCSRs_csrs_0_wdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_0_value = frontend_io_ptw_customCSRs_csrs_0_value;
    assign frontend_io_ptw_customCSRs_csrs_0_stall = frontend_tlb_io_ptw_customCSRs_csrs_0_stall;
    assign frontend_io_ptw_customCSRs_csrs_0_set = frontend_tlb_io_ptw_customCSRs_csrs_0_set;
    assign frontend_io_ptw_customCSRs_csrs_0_sdata = frontend_tlb_io_ptw_customCSRs_csrs_0_sdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_1_ren = frontend_io_ptw_customCSRs_csrs_1_ren;
    assign frontend_tlb_io_ptw_customCSRs_csrs_1_wen = frontend_io_ptw_customCSRs_csrs_1_wen;
    assign frontend_tlb_io_ptw_customCSRs_csrs_1_wdata = frontend_io_ptw_customCSRs_csrs_1_wdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_1_value = frontend_io_ptw_customCSRs_csrs_1_value;
    assign frontend_io_ptw_customCSRs_csrs_1_stall = frontend_tlb_io_ptw_customCSRs_csrs_1_stall;
    assign frontend_io_ptw_customCSRs_csrs_1_set = frontend_tlb_io_ptw_customCSRs_csrs_1_set;
    assign frontend_io_ptw_customCSRs_csrs_1_sdata = frontend_tlb_io_ptw_customCSRs_csrs_1_sdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_2_ren = frontend_io_ptw_customCSRs_csrs_2_ren;
    assign frontend_tlb_io_ptw_customCSRs_csrs_2_wen = frontend_io_ptw_customCSRs_csrs_2_wen;
    assign frontend_tlb_io_ptw_customCSRs_csrs_2_wdata = frontend_io_ptw_customCSRs_csrs_2_wdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_2_value = frontend_io_ptw_customCSRs_csrs_2_value;
    assign frontend_io_ptw_customCSRs_csrs_2_stall = frontend_tlb_io_ptw_customCSRs_csrs_2_stall;
    assign frontend_io_ptw_customCSRs_csrs_2_set = frontend_tlb_io_ptw_customCSRs_csrs_2_set;
    assign frontend_io_ptw_customCSRs_csrs_2_sdata = frontend_tlb_io_ptw_customCSRs_csrs_2_sdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_3_ren = frontend_io_ptw_customCSRs_csrs_3_ren;
    assign frontend_tlb_io_ptw_customCSRs_csrs_3_wen = frontend_io_ptw_customCSRs_csrs_3_wen;
    assign frontend_tlb_io_ptw_customCSRs_csrs_3_wdata = frontend_io_ptw_customCSRs_csrs_3_wdata;
    assign frontend_tlb_io_ptw_customCSRs_csrs_3_value = frontend_io_ptw_customCSRs_csrs_3_value;
    assign frontend_io_ptw_customCSRs_csrs_3_stall = frontend_tlb_io_ptw_customCSRs_csrs_3_stall;
    assign frontend_io_ptw_customCSRs_csrs_3_set = frontend_tlb_io_ptw_customCSRs_csrs_3_set;
    assign frontend_io_ptw_customCSRs_csrs_3_sdata = frontend_tlb_io_ptw_customCSRs_csrs_3_sdata;
    assign frontend_tlb_io_kill = frontend__GEN_6;
     
    reg frontend_s1_valid ; 
    reg frontend_s2_valid ; 
    wire frontend_s0_fq_has_space = frontend__fq_io_mask [2]==1'h0| frontend__fq_io_mask [3]==1'h0&( frontend_s1_valid ==1'h0| frontend_s2_valid ==1'h0)| frontend__fq_io_mask [4]==1'h0& frontend_s1_valid ==1'h0& frontend_s2_valid ==1'h0; 
  assign  frontend_s0_valid = frontend_io_cpu_req_valid | frontend_s0_fq_has_space ; 
    reg frontend_s1_speculative ; 
    reg frontend_s2_btb_resp_bits_taken ; 
    reg frontend_s2_tlb_resp_miss ; reg[31:0] frontend_s2_tlb_resp_paddr ; reg[33:0] frontend_s2_tlb_resp_gpa ; 
    reg frontend_s2_tlb_resp_gpa_is_pte ; 
    reg frontend_s2_tlb_resp_pf_ld ; 
    reg frontend_s2_tlb_resp_pf_st ; 
    reg frontend_s2_tlb_resp_gf_ld ; 
    reg frontend_s2_tlb_resp_gf_st ; 
    reg frontend_s2_tlb_resp_ae_ld ; 
    reg frontend_s2_tlb_resp_ae_st ; 
    reg frontend_s2_tlb_resp_ae_inst ; 
    reg frontend_s2_tlb_resp_ma_ld ; 
    reg frontend_s2_tlb_resp_ma_st ; 
    reg frontend_s2_tlb_resp_ma_inst ; 
    reg frontend_s2_tlb_resp_must_alloc ; 
    reg frontend_s2_tlb_resp_prefetchable ; 
    wire frontend_s2_xcpt = frontend_s2_tlb_resp_ae_inst | frontend_s2_tlb_resp_pf_inst | frontend_s2_tlb_resp_gf_inst ; 
    reg frontend_s2_speculative ; 
    reg frontend_s2_partial_insn_valid ; reg[15:0] frontend_s2_partial_insn ; 
    reg frontend_wrong_path ; 
    wire[33:0] frontend_s1_base_pc =~(~ frontend_s1_pc |34'h3); 
    wire[34:0] frontend__GEN_9 ={1'h0, frontend_s1_base_pc }+35'h4; 
    wire[33:0] frontend_ntpc = frontend__GEN_9 [33:0]; 
    wire[33:0] frontend_predicted_npc = frontend_ntpc ; 
    wire frontend_s2_replay ; 
    reg frontend_s2_replay_REG ; 
  assign  frontend_s2_replay = frontend_s2_valid &( frontend__fq_io_enq_ready & frontend__GEN_2 )==1'h0| frontend_s2_replay_REG ; 
    wire[33:0] frontend_npc = frontend_s2_replay  ?  frontend_s2_pc : frontend_predicted_npc ; 
    wire frontend_s0_speculative = frontend_s1_speculative | frontend_s2_valid & frontend_s2_speculative ==1'h0| frontend_predicted_taken ; 
    wire frontend__GEN_10 = frontend_s2_replay ==1'h0; 
    wire frontend__GEN_11 = frontend_s2_redirect ==1'h0; reg[1:0] frontend_recent_progress_counter ; 
    wire frontend_recent_progress = frontend_recent_progress_counter >2'h0; 
    wire frontend__GEN_12 = frontend_io_ptw_req_ready & frontend__io_ptw_req_valid_output & frontend_recent_progress ; 
    wire[2:0] frontend__GEN_13 ={1'h0, frontend_recent_progress_counter }-3'h1; 
    wire frontend_s2_kill_speculative_tlb_refill = frontend_s2_speculative & frontend_recent_progress ==1'h0; 
  assign  frontend__GEN_7 = frontend_s1_valid & frontend_s2_replay ==1'h0; 
  assign  frontend__GEN_6 = frontend_s2_valid ==1'h0| frontend_s2_kill_speculative_tlb_refill ; 
    wire[33:0] frontend__io_cpu_npc_output ; 
  assign  frontend___io_cpu_npc_output_32to0 = frontend__io_cpu_npc_output [32:0]; 
  assign  frontend__s2_pc_32to0 = frontend_s2_pc [32:0]; 
  assign  frontend__GEN_5 = frontend_s2_redirect | frontend__tlb_io_resp_miss | frontend_s2_replay ; 
    wire frontend_s2_can_speculatively_refill = frontend_s2_tlb_resp_cacheable & frontend_io_ptw_customCSRs_csrs_0_value [3]==1'h0; 
  assign  frontend__GEN_4 = frontend_s2_speculative & frontend_s2_can_speculatively_refill ==1'h0| frontend_s2_xcpt ; 
  assign  frontend__GEN_3 = frontend_s2_tlb_resp_prefetchable & frontend_io_ptw_customCSRs_csrs_0_value [17]==1'h0; 
    reg frontend_fq_io_enq_valid_REG ; 
  assign  frontend__GEN_2 = frontend_fq_io_enq_valid_REG & frontend_s2_valid &( frontend__icache_io_resp_valid | frontend_s2_kill_speculative_tlb_refill & frontend_s2_tlb_resp_miss | frontend_s2_tlb_resp_miss ==1'h0& frontend__GEN_4 ); 
  assign  frontend__io_cpu_npc_output =~(~( frontend_io_cpu_req_valid  ?  frontend_io_cpu_req_bits_pc : frontend_npc )|34'h1); 
    wire[2:0] frontend__GEN_14 =3'h3<< frontend_s2_pc [1]; 
  assign  frontend__GEN_1 = frontend__GEN_14 [1:0]; 
  assign  frontend__GEN_0 = frontend__icache_io_resp_bits_replay | frontend__GEN_4 & frontend__icache_io_resp_valid ==1'h0& frontend_s2_xcpt ==1'h0| frontend_s2_kill_speculative_tlb_refill & frontend_s2_tlb_resp_miss ; 
    wire frontend__GEN_15 =( frontend_s2_speculative & frontend_io_ptw_customCSRs_csrs_0_value [3]& frontend__GEN_4 ==1'h0)==1'h0==1'h0; 
  always @( posedge  frontend_clock )
         begin 
             if ( frontend_reset ==1'h0& frontend__GEN_8 )
                 begin 
                     if (1)$error("Assertion failed\n    at Frontend.scala:92 assert(!(io.cpu.req.valid || io.cpu.sfence.valid || io.cpu.flush_icache || io.cpu.bht_update.valid || io.cpu.btb_update.valid) || io.cpu.might_request)\n");
                     if (1)$fatal;
                 end 
             if ( frontend_reset ==1'h0& frontend__GEN_15 )
                 begin 
                     if (1)$error("Assertion failed\n    at Frontend.scala:190 assert(!(s2_speculative && io.ptw.customCSRs.asInstanceOf[RocketCustomCSRs].disableSpeculativeICacheRefill && !icache.io.s2_kill))\n");
                     if (1)$fatal;
                 end 
         end
  assign  frontend__GEN = frontend__icache_io_resp_valid & frontend__icache_io_resp_bits_ae  ? 1'h1: frontend_s2_tlb_resp_ae_inst ; 
    reg frontend_gpa_valid ; reg[33:0] frontend_gpa ; 
    wire frontend__GEN_16 = frontend__fq_io_enq_ready & frontend__GEN_2 & frontend_s2_tlb_resp_gf_inst ; 
    wire frontend__GEN_17 = frontend_gpa_valid ==1'h0; 
  always @( posedge  frontend_clock )
         begin  
             frontend_clock_en_reg  <=1'h1; 
             frontend_s1_valid  <= frontend_s0_valid ; 
             frontend_s1_pc  <= frontend__io_cpu_npc_output ;
             if ( frontend_io_cpu_req_valid )
                 begin  
                     frontend_s1_speculative  <= frontend_io_cpu_req_bits_speculative ; 
                     frontend_gpa_valid  <=1'h0;
                 end 
              else 
                 begin 
                     if ( frontend_s2_replay ) 
                         frontend_s1_speculative  <= frontend_s2_speculative ;
                      else  
                         frontend_s1_speculative  <= frontend_s0_speculative ;
                     if ( frontend__GEN_16 ) 
                         frontend_gpa_valid  <=1'h1;
                      else 
                         begin 
                         end 
                 end 
             if ( frontend__GEN_10 )
                 begin  
                     frontend_s2_tlb_resp_miss  <= frontend__tlb_io_resp_miss ; 
                     frontend_s2_tlb_resp_paddr  <= frontend__tlb_io_resp_paddr ; 
                     frontend_s2_tlb_resp_gpa  <= frontend__tlb_io_resp_gpa ; 
                     frontend_s2_tlb_resp_gpa_is_pte  <= frontend__tlb_io_resp_gpa_is_pte ; 
                     frontend_s2_tlb_resp_pf_ld  <= frontend__tlb_io_resp_pf_ld ; 
                     frontend_s2_tlb_resp_pf_st  <= frontend__tlb_io_resp_pf_st ; 
                     frontend_s2_tlb_resp_pf_inst  <= frontend__tlb_io_resp_pf_inst ; 
                     frontend_s2_tlb_resp_gf_ld  <= frontend__tlb_io_resp_gf_ld ; 
                     frontend_s2_tlb_resp_gf_st  <= frontend__tlb_io_resp_gf_st ; 
                     frontend_s2_tlb_resp_gf_inst  <= frontend__tlb_io_resp_gf_inst ; 
                     frontend_s2_tlb_resp_ae_ld  <= frontend__tlb_io_resp_ae_ld ; 
                     frontend_s2_tlb_resp_ae_st  <= frontend__tlb_io_resp_ae_st ; 
                     frontend_s2_tlb_resp_ae_inst  <= frontend__tlb_io_resp_ae_inst ; 
                     frontend_s2_tlb_resp_ma_ld  <= frontend__tlb_io_resp_ma_ld ; 
                     frontend_s2_tlb_resp_ma_st  <= frontend__tlb_io_resp_ma_st ; 
                     frontend_s2_tlb_resp_ma_inst  <= frontend__tlb_io_resp_ma_inst ; 
                     frontend_s2_tlb_resp_cacheable  <= frontend__tlb_io_resp_cacheable ; 
                     frontend_s2_tlb_resp_must_alloc  <= frontend__tlb_io_resp_must_alloc ; 
                     frontend_s2_tlb_resp_prefetchable  <= frontend__tlb_io_resp_prefetchable ;
                 end 
              else 
                 begin 
                 end  
             frontend_fq_io_enq_valid_REG  <= frontend_s1_valid ;
             if ( frontend__GEN_16 )
                 begin 
                     if ( frontend__GEN_17 ) 
                         frontend_gpa  <= frontend_s2_tlb_resp_gpa ;
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end 
         end
  always @( posedge  frontend_clock )
         begin 
             if ( frontend_reset )
                 begin  
                     frontend_s2_valid  <=1'h0; 
                     frontend_s2_pc  <={2'h0,~(~ frontend_resetVectorSinkNodeIn |32'h1)}; 
                     frontend_s2_speculative  <=1'h0; 
                     frontend_s2_partial_insn_valid  <=1'h0; 
                     frontend_wrong_path  <=1'h0; 
                     frontend_s2_replay_REG  <=1'h1; 
                     frontend_recent_progress_counter  <=2'h3;
                 end 
              else 
                 begin 
                     if ( frontend__GEN_10 )
                         begin  
                             frontend_s2_valid  <= frontend__GEN_11 ; 
                             frontend_s2_pc  <= frontend_s1_pc ; 
                             frontend_s2_speculative  <= frontend_s1_speculative ;
                         end 
                      else  
                         frontend_s2_valid  <=1'h0; 
                     frontend_s2_replay_REG  <= frontend_s2_replay & frontend_s0_valid ==1'h0;
                     if ( frontend_io_cpu_progress ) 
                         frontend_recent_progress_counter  <=2'h3;
                      else 
                         if ( frontend__GEN_12 ) 
                             frontend_recent_progress_counter  <= frontend__GEN_13 [1:0];
                          else 
                             begin 
                             end 
                 end 
         end
  assign  frontend_io_cpu_clock_enabled = frontend_clock_en ; 
  assign  frontend_io_cpu_gpa_valid = frontend_gpa_valid ; 
  assign  frontend_io_cpu_gpa_bits = frontend_gpa ; 
  assign  frontend_io_cpu_npc = frontend__io_cpu_npc_output ; 
  assign  frontend_io_cpu_perf_tlbMiss = frontend_io_ptw_req_ready & frontend__io_ptw_req_valid_output ; 
  assign  frontend_io_ptw_req_valid = frontend__io_ptw_req_valid_output ;
    assign frontend_clock = clock;
    assign frontend_reset = reset;
    assign frontend_auto_icache_master_out_a_ready = widget_1_auto_in_a_ready;
    assign widget_1_auto_in_a_valid = frontend_auto_icache_master_out_a_valid;
    assign widget_1_auto_in_a_bits_opcode = frontend_auto_icache_master_out_a_bits_opcode;
    assign widget_1_auto_in_a_bits_param = frontend_auto_icache_master_out_a_bits_param;
    assign widget_1_auto_in_a_bits_size = frontend_auto_icache_master_out_a_bits_size;
    assign widget_1_auto_in_a_bits_source = frontend_auto_icache_master_out_a_bits_source;
    assign widget_1_auto_in_a_bits_address = frontend_auto_icache_master_out_a_bits_address;
    assign widget_1_auto_in_a_bits_user_amba_prot_bufferable = frontend_auto_icache_master_out_a_bits_user_amba_prot_bufferable;
    assign widget_1_auto_in_a_bits_user_amba_prot_modifiable = frontend_auto_icache_master_out_a_bits_user_amba_prot_modifiable;
    assign widget_1_auto_in_a_bits_user_amba_prot_readalloc = frontend_auto_icache_master_out_a_bits_user_amba_prot_readalloc;
    assign widget_1_auto_in_a_bits_user_amba_prot_writealloc = frontend_auto_icache_master_out_a_bits_user_amba_prot_writealloc;
    assign widget_1_auto_in_a_bits_user_amba_prot_privileged = frontend_auto_icache_master_out_a_bits_user_amba_prot_privileged;
    assign widget_1_auto_in_a_bits_user_amba_prot_secure = frontend_auto_icache_master_out_a_bits_user_amba_prot_secure;
    assign widget_1_auto_in_a_bits_user_amba_prot_fetch = frontend_auto_icache_master_out_a_bits_user_amba_prot_fetch;
    assign widget_1_auto_in_a_bits_mask = frontend_auto_icache_master_out_a_bits_mask;
    assign widget_1_auto_in_a_bits_data = frontend_auto_icache_master_out_a_bits_data;
    assign widget_1_auto_in_a_bits_corrupt = frontend_auto_icache_master_out_a_bits_corrupt;
    assign widget_1_auto_in_d_ready = frontend_auto_icache_master_out_d_ready;
    assign frontend_auto_icache_master_out_d_valid = widget_1_auto_in_d_valid;
    assign frontend_auto_icache_master_out_d_bits_opcode = widget_1_auto_in_d_bits_opcode;
    assign frontend_auto_icache_master_out_d_bits_param = widget_1_auto_in_d_bits_param;
    assign frontend_auto_icache_master_out_d_bits_size = widget_1_auto_in_d_bits_size;
    assign frontend_auto_icache_master_out_d_bits_source = widget_1_auto_in_d_bits_source;
    assign frontend_auto_icache_master_out_d_bits_sink = widget_1_auto_in_d_bits_sink;
    assign frontend_auto_icache_master_out_d_bits_denied = widget_1_auto_in_d_bits_denied;
    assign frontend_auto_icache_master_out_d_bits_data = widget_1_auto_in_d_bits_data;
    assign frontend_auto_icache_master_out_d_bits_corrupt = widget_1_auto_in_d_bits_corrupt;
    assign frontend_auto_reset_vector_sink_in = broadcast_1_auto_out_1;
    assign frontend_io_cpu_might_request = _core_io_imem_might_request;
    assign _frontend_io_cpu_clock_enabled = frontend_io_cpu_clock_enabled;
    assign frontend_io_cpu_req_valid = _core_io_imem_req_valid;
    assign frontend_io_cpu_req_bits_pc = _core_io_imem_req_bits_pc;
    assign frontend_io_cpu_req_bits_speculative = _core_io_imem_req_bits_speculative;
    assign frontend_io_cpu_sfence_valid = _core_io_imem_sfence_valid;
    assign frontend_io_cpu_sfence_bits_rs1 = _core_io_imem_sfence_bits_rs1;
    assign frontend_io_cpu_sfence_bits_rs2 = _core_io_imem_sfence_bits_rs2;
    assign frontend_io_cpu_sfence_bits_addr = _core_io_imem_sfence_bits_addr;
    assign frontend_io_cpu_sfence_bits_asid = _core_io_imem_sfence_bits_asid;
    assign frontend_io_cpu_sfence_bits_hv = _core_io_imem_sfence_bits_hv;
    assign frontend_io_cpu_sfence_bits_hg = _core_io_imem_sfence_bits_hg;
    assign frontend_io_cpu_resp_ready = _core_io_imem_resp_ready;
    assign _frontend_io_cpu_resp_valid = frontend_io_cpu_resp_valid;
    assign _frontend_io_cpu_resp_bits_btb_cfiType = frontend_io_cpu_resp_bits_btb_cfiType;
    assign _frontend_io_cpu_resp_bits_btb_taken = frontend_io_cpu_resp_bits_btb_taken;
    assign _frontend_io_cpu_resp_bits_btb_mask = frontend_io_cpu_resp_bits_btb_mask;
    assign _frontend_io_cpu_resp_bits_btb_bridx = frontend_io_cpu_resp_bits_btb_bridx;
    assign _frontend_io_cpu_resp_bits_btb_target = frontend_io_cpu_resp_bits_btb_target;
    assign _frontend_io_cpu_resp_bits_btb_entry = frontend_io_cpu_resp_bits_btb_entry;
    assign _frontend_io_cpu_resp_bits_btb_bht_history = frontend_io_cpu_resp_bits_btb_bht_history;
    assign _frontend_io_cpu_resp_bits_btb_bht_value = frontend_io_cpu_resp_bits_btb_bht_value;
    assign _frontend_io_cpu_resp_bits_pc = frontend_io_cpu_resp_bits_pc;
    assign _frontend_io_cpu_resp_bits_data = frontend_io_cpu_resp_bits_data;
    assign _frontend_io_cpu_resp_bits_mask = frontend_io_cpu_resp_bits_mask;
    assign _frontend_io_cpu_resp_bits_xcpt_pf_inst = frontend_io_cpu_resp_bits_xcpt_pf_inst;
    assign _frontend_io_cpu_resp_bits_xcpt_gf_inst = frontend_io_cpu_resp_bits_xcpt_gf_inst;
    assign _frontend_io_cpu_resp_bits_xcpt_ae_inst = frontend_io_cpu_resp_bits_xcpt_ae_inst;
    assign _frontend_io_cpu_resp_bits_replay = frontend_io_cpu_resp_bits_replay;
    assign _frontend_io_cpu_gpa_valid = frontend_io_cpu_gpa_valid;
    assign _frontend_io_cpu_gpa_bits = frontend_io_cpu_gpa_bits;
    assign frontend_io_cpu_btb_update_valid = _core_io_imem_btb_update_valid;
    assign frontend_io_cpu_btb_update_bits_prediction_cfiType = _core_io_imem_btb_update_bits_prediction_cfiType;
    assign frontend_io_cpu_btb_update_bits_prediction_taken = _core_io_imem_btb_update_bits_prediction_taken;
    assign frontend_io_cpu_btb_update_bits_prediction_mask = _core_io_imem_btb_update_bits_prediction_mask;
    assign frontend_io_cpu_btb_update_bits_prediction_bridx = _core_io_imem_btb_update_bits_prediction_bridx;
    assign frontend_io_cpu_btb_update_bits_prediction_target = _core_io_imem_btb_update_bits_prediction_target;
    assign frontend_io_cpu_btb_update_bits_prediction_entry = _core_io_imem_btb_update_bits_prediction_entry;
    assign frontend_io_cpu_btb_update_bits_prediction_bht_history = _core_io_imem_btb_update_bits_prediction_bht_history;
    assign frontend_io_cpu_btb_update_bits_prediction_bht_value = _core_io_imem_btb_update_bits_prediction_bht_value;
    assign frontend_io_cpu_btb_update_bits_pc = _core_io_imem_btb_update_bits_pc;
    assign frontend_io_cpu_btb_update_bits_target = _core_io_imem_btb_update_bits_target;
    assign frontend_io_cpu_btb_update_bits_taken = _core_io_imem_btb_update_bits_taken;
    assign frontend_io_cpu_btb_update_bits_isValid = _core_io_imem_btb_update_bits_isValid;
    assign frontend_io_cpu_btb_update_bits_br_pc = _core_io_imem_btb_update_bits_br_pc;
    assign frontend_io_cpu_btb_update_bits_cfiType = _core_io_imem_btb_update_bits_cfiType;
    assign frontend_io_cpu_bht_update_valid = _core_io_imem_bht_update_valid;
    assign frontend_io_cpu_bht_update_bits_prediction_history = _core_io_imem_bht_update_bits_prediction_history;
    assign frontend_io_cpu_bht_update_bits_prediction_value = _core_io_imem_bht_update_bits_prediction_value;
    assign frontend_io_cpu_bht_update_bits_pc = _core_io_imem_bht_update_bits_pc;
    assign frontend_io_cpu_bht_update_bits_branch = _core_io_imem_bht_update_bits_branch;
    assign frontend_io_cpu_bht_update_bits_taken = _core_io_imem_bht_update_bits_taken;
    assign frontend_io_cpu_bht_update_bits_mispredict = _core_io_imem_bht_update_bits_mispredict;
    assign frontend_io_cpu_ras_update_valid = _core_io_imem_ras_update_valid;
    assign frontend_io_cpu_ras_update_bits_cfiType = _core_io_imem_ras_update_bits_cfiType;
    assign frontend_io_cpu_ras_update_bits_returnAddr = _core_io_imem_ras_update_bits_returnAddr;
    assign frontend_io_cpu_flush_icache = _core_io_imem_flush_icache;
    assign _frontend_io_cpu_npc = frontend_io_cpu_npc;
    assign _frontend_io_cpu_perf_acquire = frontend_io_cpu_perf_acquire;
    assign _frontend_io_cpu_perf_tlbMiss = frontend_io_cpu_perf_tlbMiss;
    assign frontend_io_cpu_progress = _core_io_imem_progress;
    assign frontend_io_ptw_req_ready = _ptw_io_requestor_1_req_ready;
    assign _frontend_io_ptw_req_valid = frontend_io_ptw_req_valid;
    assign _frontend_io_ptw_req_bits_valid = frontend_io_ptw_req_bits_valid;
    assign _frontend_io_ptw_req_bits_bits_addr = frontend_io_ptw_req_bits_bits_addr;
    assign _frontend_io_ptw_req_bits_bits_need_gpa = frontend_io_ptw_req_bits_bits_need_gpa;
    assign _frontend_io_ptw_req_bits_bits_vstage1 = frontend_io_ptw_req_bits_bits_vstage1;
    assign _frontend_io_ptw_req_bits_bits_stage2 = frontend_io_ptw_req_bits_bits_stage2;
    assign frontend_io_ptw_resp_valid = _ptw_io_requestor_1_resp_valid;
    assign frontend_io_ptw_resp_bits_ae_ptw = _ptw_io_requestor_1_resp_bits_ae_ptw;
    assign frontend_io_ptw_resp_bits_ae_final = _ptw_io_requestor_1_resp_bits_ae_final;
    assign frontend_io_ptw_resp_bits_pf = _ptw_io_requestor_1_resp_bits_pf;
    assign frontend_io_ptw_resp_bits_gf = _ptw_io_requestor_1_resp_bits_gf;
    assign frontend_io_ptw_resp_bits_hr = _ptw_io_requestor_1_resp_bits_hr;
    assign frontend_io_ptw_resp_bits_hw = _ptw_io_requestor_1_resp_bits_hw;
    assign frontend_io_ptw_resp_bits_hx = _ptw_io_requestor_1_resp_bits_hx;
    assign frontend_io_ptw_resp_bits_pte_reserved_for_future = _ptw_io_requestor_1_resp_bits_pte_reserved_for_future;
    assign frontend_io_ptw_resp_bits_pte_ppn = _ptw_io_requestor_1_resp_bits_pte_ppn;
    assign frontend_io_ptw_resp_bits_pte_reserved_for_software = _ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
    assign frontend_io_ptw_resp_bits_pte_d = _ptw_io_requestor_1_resp_bits_pte_d;
    assign frontend_io_ptw_resp_bits_pte_a = _ptw_io_requestor_1_resp_bits_pte_a;
    assign frontend_io_ptw_resp_bits_pte_g = _ptw_io_requestor_1_resp_bits_pte_g;
    assign frontend_io_ptw_resp_bits_pte_u = _ptw_io_requestor_1_resp_bits_pte_u;
    assign frontend_io_ptw_resp_bits_pte_x = _ptw_io_requestor_1_resp_bits_pte_x;
    assign frontend_io_ptw_resp_bits_pte_w = _ptw_io_requestor_1_resp_bits_pte_w;
    assign frontend_io_ptw_resp_bits_pte_r = _ptw_io_requestor_1_resp_bits_pte_r;
    assign frontend_io_ptw_resp_bits_pte_v = _ptw_io_requestor_1_resp_bits_pte_v;
    assign frontend_io_ptw_resp_bits_level = _ptw_io_requestor_1_resp_bits_level;
    assign frontend_io_ptw_resp_bits_fragmented_superpage = _ptw_io_requestor_1_resp_bits_fragmented_superpage;
    assign frontend_io_ptw_resp_bits_homogeneous = _ptw_io_requestor_1_resp_bits_homogeneous;
    assign frontend_io_ptw_resp_bits_gpa_valid = _ptw_io_requestor_1_resp_bits_gpa_valid;
    assign frontend_io_ptw_resp_bits_gpa_bits = _ptw_io_requestor_1_resp_bits_gpa_bits;
    assign frontend_io_ptw_resp_bits_gpa_is_pte = _ptw_io_requestor_1_resp_bits_gpa_is_pte;
    assign frontend_io_ptw_ptbr_mode = _ptw_io_requestor_1_ptbr_mode;
    assign frontend_io_ptw_ptbr_asid = _ptw_io_requestor_1_ptbr_asid;
    assign frontend_io_ptw_ptbr_ppn = _ptw_io_requestor_1_ptbr_ppn;
    assign frontend_io_ptw_hgatp_mode = _ptw_io_requestor_1_hgatp_mode;
    assign frontend_io_ptw_hgatp_asid = _ptw_io_requestor_1_hgatp_asid;
    assign frontend_io_ptw_hgatp_ppn = _ptw_io_requestor_1_hgatp_ppn;
    assign frontend_io_ptw_vsatp_mode = _ptw_io_requestor_1_vsatp_mode;
    assign frontend_io_ptw_vsatp_asid = _ptw_io_requestor_1_vsatp_asid;
    assign frontend_io_ptw_vsatp_ppn = _ptw_io_requestor_1_vsatp_ppn;
    assign frontend_io_ptw_status_debug = _ptw_io_requestor_1_status_debug;
    assign frontend_io_ptw_status_cease = _ptw_io_requestor_1_status_cease;
    assign frontend_io_ptw_status_wfi = _ptw_io_requestor_1_status_wfi;
    assign frontend_io_ptw_status_isa = _ptw_io_requestor_1_status_isa;
    assign frontend_io_ptw_status_dprv = _ptw_io_requestor_1_status_dprv;
    assign frontend_io_ptw_status_dv = _ptw_io_requestor_1_status_dv;
    assign frontend_io_ptw_status_prv = _ptw_io_requestor_1_status_prv;
    assign frontend_io_ptw_status_v = _ptw_io_requestor_1_status_v;
    assign frontend_io_ptw_status_sd = _ptw_io_requestor_1_status_sd;
    assign frontend_io_ptw_status_zero2 = _ptw_io_requestor_1_status_zero2;
    assign frontend_io_ptw_status_mpv = _ptw_io_requestor_1_status_mpv;
    assign frontend_io_ptw_status_gva = _ptw_io_requestor_1_status_gva;
    assign frontend_io_ptw_status_mbe = _ptw_io_requestor_1_status_mbe;
    assign frontend_io_ptw_status_sbe = _ptw_io_requestor_1_status_sbe;
    assign frontend_io_ptw_status_sxl = _ptw_io_requestor_1_status_sxl;
    assign frontend_io_ptw_status_uxl = _ptw_io_requestor_1_status_uxl;
    assign frontend_io_ptw_status_sd_rv32 = _ptw_io_requestor_1_status_sd_rv32;
    assign frontend_io_ptw_status_zero1 = _ptw_io_requestor_1_status_zero1;
    assign frontend_io_ptw_status_tsr = _ptw_io_requestor_1_status_tsr;
    assign frontend_io_ptw_status_tw = _ptw_io_requestor_1_status_tw;
    assign frontend_io_ptw_status_tvm = _ptw_io_requestor_1_status_tvm;
    assign frontend_io_ptw_status_mxr = _ptw_io_requestor_1_status_mxr;
    assign frontend_io_ptw_status_sum = _ptw_io_requestor_1_status_sum;
    assign frontend_io_ptw_status_mprv = _ptw_io_requestor_1_status_mprv;
    assign frontend_io_ptw_status_xs = _ptw_io_requestor_1_status_xs;
    assign frontend_io_ptw_status_fs = _ptw_io_requestor_1_status_fs;
    assign frontend_io_ptw_status_mpp = _ptw_io_requestor_1_status_mpp;
    assign frontend_io_ptw_status_vs = _ptw_io_requestor_1_status_vs;
    assign frontend_io_ptw_status_spp = _ptw_io_requestor_1_status_spp;
    assign frontend_io_ptw_status_mpie = _ptw_io_requestor_1_status_mpie;
    assign frontend_io_ptw_status_ube = _ptw_io_requestor_1_status_ube;
    assign frontend_io_ptw_status_spie = _ptw_io_requestor_1_status_spie;
    assign frontend_io_ptw_status_upie = _ptw_io_requestor_1_status_upie;
    assign frontend_io_ptw_status_mie = _ptw_io_requestor_1_status_mie;
    assign frontend_io_ptw_status_hie = _ptw_io_requestor_1_status_hie;
    assign frontend_io_ptw_status_sie = _ptw_io_requestor_1_status_sie;
    assign frontend_io_ptw_status_uie = _ptw_io_requestor_1_status_uie;
    assign frontend_io_ptw_hstatus_zero6 = _ptw_io_requestor_1_hstatus_zero6;
    assign frontend_io_ptw_hstatus_vsxl = _ptw_io_requestor_1_hstatus_vsxl;
    assign frontend_io_ptw_hstatus_zero5 = _ptw_io_requestor_1_hstatus_zero5;
    assign frontend_io_ptw_hstatus_vtsr = _ptw_io_requestor_1_hstatus_vtsr;
    assign frontend_io_ptw_hstatus_vtw = _ptw_io_requestor_1_hstatus_vtw;
    assign frontend_io_ptw_hstatus_vtvm = _ptw_io_requestor_1_hstatus_vtvm;
    assign frontend_io_ptw_hstatus_zero3 = _ptw_io_requestor_1_hstatus_zero3;
    assign frontend_io_ptw_hstatus_vgein = _ptw_io_requestor_1_hstatus_vgein;
    assign frontend_io_ptw_hstatus_zero2 = _ptw_io_requestor_1_hstatus_zero2;
    assign frontend_io_ptw_hstatus_hu = _ptw_io_requestor_1_hstatus_hu;
    assign frontend_io_ptw_hstatus_spvp = _ptw_io_requestor_1_hstatus_spvp;
    assign frontend_io_ptw_hstatus_spv = _ptw_io_requestor_1_hstatus_spv;
    assign frontend_io_ptw_hstatus_gva = _ptw_io_requestor_1_hstatus_gva;
    assign frontend_io_ptw_hstatus_vsbe = _ptw_io_requestor_1_hstatus_vsbe;
    assign frontend_io_ptw_hstatus_zero1 = _ptw_io_requestor_1_hstatus_zero1;
    assign frontend_io_ptw_gstatus_debug = _ptw_io_requestor_1_gstatus_debug;
    assign frontend_io_ptw_gstatus_cease = _ptw_io_requestor_1_gstatus_cease;
    assign frontend_io_ptw_gstatus_wfi = _ptw_io_requestor_1_gstatus_wfi;
    assign frontend_io_ptw_gstatus_isa = _ptw_io_requestor_1_gstatus_isa;
    assign frontend_io_ptw_gstatus_dprv = _ptw_io_requestor_1_gstatus_dprv;
    assign frontend_io_ptw_gstatus_dv = _ptw_io_requestor_1_gstatus_dv;
    assign frontend_io_ptw_gstatus_prv = _ptw_io_requestor_1_gstatus_prv;
    assign frontend_io_ptw_gstatus_v = _ptw_io_requestor_1_gstatus_v;
    assign frontend_io_ptw_gstatus_sd = _ptw_io_requestor_1_gstatus_sd;
    assign frontend_io_ptw_gstatus_zero2 = _ptw_io_requestor_1_gstatus_zero2;
    assign frontend_io_ptw_gstatus_mpv = _ptw_io_requestor_1_gstatus_mpv;
    assign frontend_io_ptw_gstatus_gva = _ptw_io_requestor_1_gstatus_gva;
    assign frontend_io_ptw_gstatus_mbe = _ptw_io_requestor_1_gstatus_mbe;
    assign frontend_io_ptw_gstatus_sbe = _ptw_io_requestor_1_gstatus_sbe;
    assign frontend_io_ptw_gstatus_sxl = _ptw_io_requestor_1_gstatus_sxl;
    assign frontend_io_ptw_gstatus_uxl = _ptw_io_requestor_1_gstatus_uxl;
    assign frontend_io_ptw_gstatus_sd_rv32 = _ptw_io_requestor_1_gstatus_sd_rv32;
    assign frontend_io_ptw_gstatus_zero1 = _ptw_io_requestor_1_gstatus_zero1;
    assign frontend_io_ptw_gstatus_tsr = _ptw_io_requestor_1_gstatus_tsr;
    assign frontend_io_ptw_gstatus_tw = _ptw_io_requestor_1_gstatus_tw;
    assign frontend_io_ptw_gstatus_tvm = _ptw_io_requestor_1_gstatus_tvm;
    assign frontend_io_ptw_gstatus_mxr = _ptw_io_requestor_1_gstatus_mxr;
    assign frontend_io_ptw_gstatus_sum = _ptw_io_requestor_1_gstatus_sum;
    assign frontend_io_ptw_gstatus_mprv = _ptw_io_requestor_1_gstatus_mprv;
    assign frontend_io_ptw_gstatus_xs = _ptw_io_requestor_1_gstatus_xs;
    assign frontend_io_ptw_gstatus_fs = _ptw_io_requestor_1_gstatus_fs;
    assign frontend_io_ptw_gstatus_mpp = _ptw_io_requestor_1_gstatus_mpp;
    assign frontend_io_ptw_gstatus_vs = _ptw_io_requestor_1_gstatus_vs;
    assign frontend_io_ptw_gstatus_spp = _ptw_io_requestor_1_gstatus_spp;
    assign frontend_io_ptw_gstatus_mpie = _ptw_io_requestor_1_gstatus_mpie;
    assign frontend_io_ptw_gstatus_ube = _ptw_io_requestor_1_gstatus_ube;
    assign frontend_io_ptw_gstatus_spie = _ptw_io_requestor_1_gstatus_spie;
    assign frontend_io_ptw_gstatus_upie = _ptw_io_requestor_1_gstatus_upie;
    assign frontend_io_ptw_gstatus_mie = _ptw_io_requestor_1_gstatus_mie;
    assign frontend_io_ptw_gstatus_hie = _ptw_io_requestor_1_gstatus_hie;
    assign frontend_io_ptw_gstatus_sie = _ptw_io_requestor_1_gstatus_sie;
    assign frontend_io_ptw_gstatus_uie = _ptw_io_requestor_1_gstatus_uie;
    assign frontend_io_ptw_pmp_0_cfg_l = _ptw_io_requestor_1_pmp_0_cfg_l;
    assign frontend_io_ptw_pmp_0_cfg_res = _ptw_io_requestor_1_pmp_0_cfg_res;
    assign frontend_io_ptw_pmp_0_cfg_a = _ptw_io_requestor_1_pmp_0_cfg_a;
    assign frontend_io_ptw_pmp_0_cfg_x = _ptw_io_requestor_1_pmp_0_cfg_x;
    assign frontend_io_ptw_pmp_0_cfg_w = _ptw_io_requestor_1_pmp_0_cfg_w;
    assign frontend_io_ptw_pmp_0_cfg_r = _ptw_io_requestor_1_pmp_0_cfg_r;
    assign frontend_io_ptw_pmp_0_addr = _ptw_io_requestor_1_pmp_0_addr;
    assign frontend_io_ptw_pmp_0_mask = _ptw_io_requestor_1_pmp_0_mask;
    assign frontend_io_ptw_pmp_1_cfg_l = _ptw_io_requestor_1_pmp_1_cfg_l;
    assign frontend_io_ptw_pmp_1_cfg_res = _ptw_io_requestor_1_pmp_1_cfg_res;
    assign frontend_io_ptw_pmp_1_cfg_a = _ptw_io_requestor_1_pmp_1_cfg_a;
    assign frontend_io_ptw_pmp_1_cfg_x = _ptw_io_requestor_1_pmp_1_cfg_x;
    assign frontend_io_ptw_pmp_1_cfg_w = _ptw_io_requestor_1_pmp_1_cfg_w;
    assign frontend_io_ptw_pmp_1_cfg_r = _ptw_io_requestor_1_pmp_1_cfg_r;
    assign frontend_io_ptw_pmp_1_addr = _ptw_io_requestor_1_pmp_1_addr;
    assign frontend_io_ptw_pmp_1_mask = _ptw_io_requestor_1_pmp_1_mask;
    assign frontend_io_ptw_pmp_2_cfg_l = _ptw_io_requestor_1_pmp_2_cfg_l;
    assign frontend_io_ptw_pmp_2_cfg_res = _ptw_io_requestor_1_pmp_2_cfg_res;
    assign frontend_io_ptw_pmp_2_cfg_a = _ptw_io_requestor_1_pmp_2_cfg_a;
    assign frontend_io_ptw_pmp_2_cfg_x = _ptw_io_requestor_1_pmp_2_cfg_x;
    assign frontend_io_ptw_pmp_2_cfg_w = _ptw_io_requestor_1_pmp_2_cfg_w;
    assign frontend_io_ptw_pmp_2_cfg_r = _ptw_io_requestor_1_pmp_2_cfg_r;
    assign frontend_io_ptw_pmp_2_addr = _ptw_io_requestor_1_pmp_2_addr;
    assign frontend_io_ptw_pmp_2_mask = _ptw_io_requestor_1_pmp_2_mask;
    assign frontend_io_ptw_pmp_3_cfg_l = _ptw_io_requestor_1_pmp_3_cfg_l;
    assign frontend_io_ptw_pmp_3_cfg_res = _ptw_io_requestor_1_pmp_3_cfg_res;
    assign frontend_io_ptw_pmp_3_cfg_a = _ptw_io_requestor_1_pmp_3_cfg_a;
    assign frontend_io_ptw_pmp_3_cfg_x = _ptw_io_requestor_1_pmp_3_cfg_x;
    assign frontend_io_ptw_pmp_3_cfg_w = _ptw_io_requestor_1_pmp_3_cfg_w;
    assign frontend_io_ptw_pmp_3_cfg_r = _ptw_io_requestor_1_pmp_3_cfg_r;
    assign frontend_io_ptw_pmp_3_addr = _ptw_io_requestor_1_pmp_3_addr;
    assign frontend_io_ptw_pmp_3_mask = _ptw_io_requestor_1_pmp_3_mask;
    assign frontend_io_ptw_pmp_4_cfg_l = _ptw_io_requestor_1_pmp_4_cfg_l;
    assign frontend_io_ptw_pmp_4_cfg_res = _ptw_io_requestor_1_pmp_4_cfg_res;
    assign frontend_io_ptw_pmp_4_cfg_a = _ptw_io_requestor_1_pmp_4_cfg_a;
    assign frontend_io_ptw_pmp_4_cfg_x = _ptw_io_requestor_1_pmp_4_cfg_x;
    assign frontend_io_ptw_pmp_4_cfg_w = _ptw_io_requestor_1_pmp_4_cfg_w;
    assign frontend_io_ptw_pmp_4_cfg_r = _ptw_io_requestor_1_pmp_4_cfg_r;
    assign frontend_io_ptw_pmp_4_addr = _ptw_io_requestor_1_pmp_4_addr;
    assign frontend_io_ptw_pmp_4_mask = _ptw_io_requestor_1_pmp_4_mask;
    assign frontend_io_ptw_pmp_5_cfg_l = _ptw_io_requestor_1_pmp_5_cfg_l;
    assign frontend_io_ptw_pmp_5_cfg_res = _ptw_io_requestor_1_pmp_5_cfg_res;
    assign frontend_io_ptw_pmp_5_cfg_a = _ptw_io_requestor_1_pmp_5_cfg_a;
    assign frontend_io_ptw_pmp_5_cfg_x = _ptw_io_requestor_1_pmp_5_cfg_x;
    assign frontend_io_ptw_pmp_5_cfg_w = _ptw_io_requestor_1_pmp_5_cfg_w;
    assign frontend_io_ptw_pmp_5_cfg_r = _ptw_io_requestor_1_pmp_5_cfg_r;
    assign frontend_io_ptw_pmp_5_addr = _ptw_io_requestor_1_pmp_5_addr;
    assign frontend_io_ptw_pmp_5_mask = _ptw_io_requestor_1_pmp_5_mask;
    assign frontend_io_ptw_pmp_6_cfg_l = _ptw_io_requestor_1_pmp_6_cfg_l;
    assign frontend_io_ptw_pmp_6_cfg_res = _ptw_io_requestor_1_pmp_6_cfg_res;
    assign frontend_io_ptw_pmp_6_cfg_a = _ptw_io_requestor_1_pmp_6_cfg_a;
    assign frontend_io_ptw_pmp_6_cfg_x = _ptw_io_requestor_1_pmp_6_cfg_x;
    assign frontend_io_ptw_pmp_6_cfg_w = _ptw_io_requestor_1_pmp_6_cfg_w;
    assign frontend_io_ptw_pmp_6_cfg_r = _ptw_io_requestor_1_pmp_6_cfg_r;
    assign frontend_io_ptw_pmp_6_addr = _ptw_io_requestor_1_pmp_6_addr;
    assign frontend_io_ptw_pmp_6_mask = _ptw_io_requestor_1_pmp_6_mask;
    assign frontend_io_ptw_pmp_7_cfg_l = _ptw_io_requestor_1_pmp_7_cfg_l;
    assign frontend_io_ptw_pmp_7_cfg_res = _ptw_io_requestor_1_pmp_7_cfg_res;
    assign frontend_io_ptw_pmp_7_cfg_a = _ptw_io_requestor_1_pmp_7_cfg_a;
    assign frontend_io_ptw_pmp_7_cfg_x = _ptw_io_requestor_1_pmp_7_cfg_x;
    assign frontend_io_ptw_pmp_7_cfg_w = _ptw_io_requestor_1_pmp_7_cfg_w;
    assign frontend_io_ptw_pmp_7_cfg_r = _ptw_io_requestor_1_pmp_7_cfg_r;
    assign frontend_io_ptw_pmp_7_addr = _ptw_io_requestor_1_pmp_7_addr;
    assign frontend_io_ptw_pmp_7_mask = _ptw_io_requestor_1_pmp_7_mask;
    assign frontend_io_ptw_customCSRs_csrs_0_ren = _ptw_io_requestor_1_customCSRs_csrs_0_ren;
    assign frontend_io_ptw_customCSRs_csrs_0_wen = _ptw_io_requestor_1_customCSRs_csrs_0_wen;
    assign frontend_io_ptw_customCSRs_csrs_0_wdata = _ptw_io_requestor_1_customCSRs_csrs_0_wdata;
    assign frontend_io_ptw_customCSRs_csrs_0_value = _ptw_io_requestor_1_customCSRs_csrs_0_value;
    assign _frontend_io_ptw_customCSRs_csrs_0_stall = frontend_io_ptw_customCSRs_csrs_0_stall;
    assign _frontend_io_ptw_customCSRs_csrs_0_set = frontend_io_ptw_customCSRs_csrs_0_set;
    assign _frontend_io_ptw_customCSRs_csrs_0_sdata = frontend_io_ptw_customCSRs_csrs_0_sdata;
    assign frontend_io_ptw_customCSRs_csrs_1_ren = _ptw_io_requestor_1_customCSRs_csrs_1_ren;
    assign frontend_io_ptw_customCSRs_csrs_1_wen = _ptw_io_requestor_1_customCSRs_csrs_1_wen;
    assign frontend_io_ptw_customCSRs_csrs_1_wdata = _ptw_io_requestor_1_customCSRs_csrs_1_wdata;
    assign frontend_io_ptw_customCSRs_csrs_1_value = _ptw_io_requestor_1_customCSRs_csrs_1_value;
    assign _frontend_io_ptw_customCSRs_csrs_1_stall = frontend_io_ptw_customCSRs_csrs_1_stall;
    assign _frontend_io_ptw_customCSRs_csrs_1_set = frontend_io_ptw_customCSRs_csrs_1_set;
    assign _frontend_io_ptw_customCSRs_csrs_1_sdata = frontend_io_ptw_customCSRs_csrs_1_sdata;
    assign frontend_io_ptw_customCSRs_csrs_2_ren = _ptw_io_requestor_1_customCSRs_csrs_2_ren;
    assign frontend_io_ptw_customCSRs_csrs_2_wen = _ptw_io_requestor_1_customCSRs_csrs_2_wen;
    assign frontend_io_ptw_customCSRs_csrs_2_wdata = _ptw_io_requestor_1_customCSRs_csrs_2_wdata;
    assign frontend_io_ptw_customCSRs_csrs_2_value = _ptw_io_requestor_1_customCSRs_csrs_2_value;
    assign _frontend_io_ptw_customCSRs_csrs_2_stall = frontend_io_ptw_customCSRs_csrs_2_stall;
    assign _frontend_io_ptw_customCSRs_csrs_2_set = frontend_io_ptw_customCSRs_csrs_2_set;
    assign _frontend_io_ptw_customCSRs_csrs_2_sdata = frontend_io_ptw_customCSRs_csrs_2_sdata;
    assign frontend_io_ptw_customCSRs_csrs_3_ren = _ptw_io_requestor_1_customCSRs_csrs_3_ren;
    assign frontend_io_ptw_customCSRs_csrs_3_wen = _ptw_io_requestor_1_customCSRs_csrs_3_wen;
    assign frontend_io_ptw_customCSRs_csrs_3_wdata = _ptw_io_requestor_1_customCSRs_csrs_3_wdata;
    assign frontend_io_ptw_customCSRs_csrs_3_value = _ptw_io_requestor_1_customCSRs_csrs_3_value;
    assign _frontend_io_ptw_customCSRs_csrs_3_stall = frontend_io_ptw_customCSRs_csrs_3_stall;
    assign _frontend_io_ptw_customCSRs_csrs_3_set = frontend_io_ptw_customCSRs_csrs_3_set;
    assign _frontend_io_ptw_customCSRs_csrs_3_sdata = frontend_io_ptw_customCSRs_csrs_3_sdata;
    
  wire        widget_1_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_valid = widget_1_auto_in_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_1_nodeIn_a_bits_opcode = widget_1_auto_in_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_1_nodeIn_a_bits_param = widget_1_auto_in_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_1_nodeIn_a_bits_size = widget_1_auto_in_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_source = widget_1_auto_in_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] widget_1_nodeIn_a_bits_address = widget_1_auto_in_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_bufferable =
    widget_1_auto_in_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_modifiable =
    widget_1_auto_in_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_readalloc =
    widget_1_auto_in_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_writealloc =
    widget_1_auto_in_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_privileged =
    widget_1_auto_in_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_secure =
    widget_1_auto_in_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_user_amba_prot_fetch =
    widget_1_auto_in_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  widget_1_nodeIn_a_bits_mask = widget_1_auto_in_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_1_nodeIn_a_bits_data = widget_1_auto_in_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_a_bits_corrupt = widget_1_auto_in_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_ready = widget_1_auto_in_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  widget_1_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_1_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  widget_1_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  widget_1_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] widget_1_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1_nodeOut_a_ready = widget_1_auto_out_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_1_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_1_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_1_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] widget_1_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  widget_1_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_1_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_valid = widget_1_auto_out_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  widget_1_nodeOut_d_bits_opcode = widget_1_auto_out_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_1_nodeOut_d_bits_param = widget_1_auto_out_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  widget_1_nodeOut_d_bits_size = widget_1_auto_out_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_source = widget_1_auto_out_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  widget_1_nodeOut_d_bits_sink = widget_1_auto_out_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_denied = widget_1_auto_out_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] widget_1_nodeOut_d_bits_data = widget_1_auto_out_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        widget_1_nodeOut_d_bits_corrupt = widget_1_auto_out_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_nodeIn_a_ready = widget_1_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_auto_out_a_valid = widget_1_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_opcode = widget_1_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_param = widget_1_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_size = widget_1_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_source = widget_1_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_address = widget_1_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_bufferable =
    widget_1_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_modifiable =
    widget_1_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_readalloc =
    widget_1_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_writealloc =
    widget_1_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_privileged =
    widget_1_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_secure =
    widget_1_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_user_amba_prot_fetch =
    widget_1_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_mask = widget_1_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_data = widget_1_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_a_bits_corrupt = widget_1_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_auto_out_d_ready = widget_1_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign widget_1_nodeIn_d_valid = widget_1_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_opcode = widget_1_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_param = widget_1_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_size = widget_1_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_source = widget_1_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_sink = widget_1_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_denied = widget_1_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_data = widget_1_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeIn_d_bits_corrupt = widget_1_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_auto_in_a_ready = widget_1_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_nodeOut_a_valid = widget_1_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_opcode = widget_1_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_param = widget_1_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_size = widget_1_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_source = widget_1_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_address = widget_1_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_bufferable =
    widget_1_nodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_modifiable =
    widget_1_nodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_readalloc =
    widget_1_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_writealloc =
    widget_1_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_privileged =
    widget_1_nodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_secure =
    widget_1_nodeIn_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_user_amba_prot_fetch =
    widget_1_nodeIn_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_mask = widget_1_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_data = widget_1_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_a_bits_corrupt = widget_1_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_nodeOut_d_ready = widget_1_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign widget_1_auto_in_d_valid = widget_1_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_opcode = widget_1_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_param = widget_1_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_size = widget_1_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_source = widget_1_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_sink = widget_1_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_denied = widget_1_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_data = widget_1_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign widget_1_auto_in_d_bits_corrupt = widget_1_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        widget_1__63 = widget_1__26;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [2:0]  widget_1__64 = widget_1__2;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [1:0]  widget_1__65 = widget_1__8;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [3:0]  widget_1__66 = widget_1__12;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__67 = widget_1__28;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [31:0] widget_1__68 = widget_1__16;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [7:0]  widget_1__69 = widget_1__20;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [63:0] widget_1__70 = widget_1__22;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__71 = widget_1__29;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__72 = widget_1__32;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [2:0]  widget_1__73 = widget_1__3;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [2:0]  widget_1__74 = widget_1__4;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [3:0]  widget_1__75 = widget_1__13;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__76 = widget_1__33;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [31:0] widget_1__77 = widget_1__17;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__78 = widget_1__34;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__79 = widget_1__35;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__80 = widget_1__36;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__81 = widget_1__37;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__82 = widget_1__38;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__83 = widget_1__39;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__84 = widget_1__40;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [63:0] widget_1__85 = widget_1__23;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__86 = widget_1__41;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__87 = widget_1__43;	// src/main/scala/tilelink/Bundles.scala:262:{61,74}
  wire [1:0]  widget_1__88 = widget_1__9;	// src/main/scala/tilelink/Bundles.scala:262:{61,74}
  wire        widget_1__89 = widget_1__45;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [2:0]  widget_1__90 = widget_1__5;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [1:0]  widget_1__91 = widget_1__10;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [3:0]  widget_1__92 = widget_1__14;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__93 = widget_1__46;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [31:0] widget_1__94 = widget_1__18;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [7:0]  widget_1__95 = widget_1__21;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire [63:0] widget_1__96 = widget_1__24;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__97 = widget_1__47;	// src/main/scala/tilelink/Bundles.scala:259:{61,74}
  wire        widget_1__98 = widget_1__48;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [2:0]  widget_1__99 = widget_1__6;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [2:0]  widget_1__100 = widget_1__7;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [3:0]  widget_1__101 = widget_1__15;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__102 = widget_1__50;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [31:0] widget_1__103 = widget_1__19;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__104 = widget_1__51;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__105 = widget_1__52;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__106 = widget_1__53;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__107 = widget_1__54;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__108 = widget_1__55;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__109 = widget_1__56;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__110 = widget_1__57;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire [63:0] widget_1__111 = widget_1__25;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__112 = widget_1__58;	// src/main/scala/tilelink/Bundles.scala:260:{61,74}
  wire        widget_1__113 = widget_1__60;	// src/main/scala/tilelink/Bundles.scala:262:{61,74}
  wire [1:0]  widget_1__114 = widget_1__11;	// src/main/scala/tilelink/Bundles.scala:262:{61,74}
  wire        buffer_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_ready = buffer_auto_in_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlOtherMastersNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_valid = buffer_auto_in_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeIn_a_bits_opcode = buffer_auto_in_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeIn_a_bits_param = buffer_auto_in_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeIn_a_bits_size = buffer_auto_in_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_a_bits_source = buffer_auto_in_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeIn_a_bits_address = buffer_auto_in_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_bufferable =
    buffer_auto_in_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_modifiable =
    buffer_auto_in_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_readalloc =
    buffer_auto_in_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_writealloc =
    buffer_auto_in_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_privileged =
    buffer_auto_in_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_secure =
    buffer_auto_in_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_user_amba_prot_fetch =
    buffer_auto_in_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  tlOtherMastersNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  buffer_nodeIn_a_bits_mask = buffer_auto_in_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeIn_a_bits_data = buffer_auto_in_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_a_bits_corrupt = buffer_auto_in_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_b_ready = buffer_auto_in_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeIn_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_nodeIn_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_b_valid = buffer_auto_in_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_b_bits_opcode = buffer_auto_in_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeIn_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_b_bits_param = buffer_auto_in_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeOut_b_bits_size = buffer_auto_in_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeIn_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_b_bits_source = buffer_auto_in_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  buffer_nodeIn_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeOut_b_bits_address = buffer_auto_in_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeIn_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [7:0]  tlOtherMastersNodeOut_b_bits_mask = buffer_auto_in_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeOut_b_bits_data = buffer_auto_in_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_b_bits_corrupt = buffer_auto_in_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlOtherMastersNodeOut_c_ready = buffer_auto_in_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlOtherMastersNodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_valid = buffer_auto_in_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeIn_c_bits_opcode = buffer_auto_in_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeIn_c_bits_param = buffer_auto_in_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeIn_c_bits_size = buffer_auto_in_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_c_bits_source = buffer_auto_in_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [31:0] tlOtherMastersNodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeIn_c_bits_address = buffer_auto_in_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_bufferable =
    buffer_auto_in_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_modifiable =
    buffer_auto_in_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_readalloc =
    buffer_auto_in_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_writealloc =
    buffer_auto_in_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_privileged =
    buffer_auto_in_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_secure =
    buffer_auto_in_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_user_amba_prot_fetch =
    buffer_auto_in_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeIn_c_bits_data = buffer_auto_in_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_c_bits_corrupt = buffer_auto_in_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_d_ready = buffer_auto_in_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  buffer_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_d_valid = buffer_auto_in_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [2:0]  tlOtherMastersNodeOut_d_bits_opcode = buffer_auto_in_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_d_bits_param = buffer_auto_in_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [3:0]  tlOtherMastersNodeOut_d_bits_size = buffer_auto_in_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_d_bits_source = buffer_auto_in_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_d_bits_sink = buffer_auto_in_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_d_bits_denied = buffer_auto_in_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [63:0] tlOtherMastersNodeOut_d_bits_data = buffer_auto_in_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        tlOtherMastersNodeOut_d_bits_corrupt = buffer_auto_in_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlOtherMastersNodeOut_e_ready = buffer_auto_in_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        tlOtherMastersNodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeIn_e_valid = buffer_auto_in_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire [1:0]  tlOtherMastersNodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeIn_e_bits_sink = buffer_auto_in_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  wire        buffer_nodeOut_a_ready = buffer_auto_out_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  buffer_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_b_valid = buffer_auto_out_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_b_bits_opcode = buffer_auto_out_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_b_bits_param = buffer_auto_out_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_b_bits_size = buffer_auto_out_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_b_bits_source = buffer_auto_out_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_b_bits_address = buffer_auto_out_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  buffer_nodeOut_b_bits_mask = buffer_auto_out_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeOut_b_bits_data = buffer_auto_out_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_b_bits_corrupt = buffer_auto_out_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_ready = buffer_auto_out_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_nodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_valid = buffer_auto_out_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_nodeOut_d_bits_opcode = buffer_auto_out_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_d_bits_param = buffer_auto_out_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_nodeOut_d_bits_size = buffer_auto_out_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_d_bits_source = buffer_auto_out_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_d_bits_sink = buffer_auto_out_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_denied = buffer_auto_out_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_nodeOut_d_bits_data = buffer_auto_out_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_d_bits_corrupt = buffer_auto_out_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_e_ready = buffer_auto_out_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_nodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_nodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_nodeIn_a_ready = buffer_nodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_auto_out_a_valid = buffer_nodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_auto_out_a_bits_opcode = buffer_nodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_auto_out_a_bits_param = buffer_nodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_auto_out_a_bits_size = buffer_nodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_auto_out_a_bits_source = buffer_nodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_auto_out_a_bits_address = buffer_nodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_bufferable =
    buffer_nodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_modifiable =
    buffer_nodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_readalloc =
    buffer_nodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_writealloc =
    buffer_nodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_privileged =
    buffer_nodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_secure =
    buffer_nodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_user_amba_prot_fetch =
    buffer_nodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [7:0]  buffer_auto_out_a_bits_mask = buffer_nodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_auto_out_a_bits_data = buffer_nodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_a_bits_corrupt = buffer_nodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_b_ready = buffer_nodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_nodeIn_b_valid = buffer_nodeOut_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_opcode = buffer_nodeOut_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_param = buffer_nodeOut_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_size = buffer_nodeOut_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_source = buffer_nodeOut_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_address = buffer_nodeOut_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_mask = buffer_nodeOut_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_data = buffer_nodeOut_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_b_bits_corrupt = buffer_nodeOut_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_c_ready = buffer_nodeOut_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_auto_out_c_valid = buffer_nodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_auto_out_c_bits_opcode = buffer_nodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [2:0]  buffer_auto_out_c_bits_param = buffer_nodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [3:0]  buffer_auto_out_c_bits_size = buffer_nodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_auto_out_c_bits_source = buffer_nodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [31:0] buffer_auto_out_c_bits_address = buffer_nodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_bufferable =
    buffer_nodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_modifiable =
    buffer_nodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_readalloc =
    buffer_nodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_writealloc =
    buffer_nodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_privileged =
    buffer_nodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_secure =
    buffer_nodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_user_amba_prot_fetch =
    buffer_nodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [63:0] buffer_auto_out_c_bits_data = buffer_nodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_c_bits_corrupt = buffer_nodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire        buffer_auto_out_d_ready = buffer_nodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_nodeIn_d_valid = buffer_nodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_opcode = buffer_nodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_param = buffer_nodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_size = buffer_nodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_source = buffer_nodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_sink = buffer_nodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_denied = buffer_nodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_data = buffer_nodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_d_bits_corrupt = buffer_nodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeIn_e_ready = buffer_nodeOut_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire        buffer_auto_out_e_valid = buffer_nodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  wire [1:0]  buffer_auto_out_e_bits_sink = buffer_nodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_ready = buffer_nodeIn_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeOut_a_valid = buffer_nodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_opcode = buffer_nodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_param = buffer_nodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_size = buffer_nodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_source = buffer_nodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_address = buffer_nodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_bufferable =
    buffer_nodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_modifiable =
    buffer_nodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_readalloc =
    buffer_nodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_writealloc =
    buffer_nodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_privileged =
    buffer_nodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_secure =
    buffer_nodeIn_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_user_amba_prot_fetch =
    buffer_nodeIn_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_mask = buffer_nodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_data = buffer_nodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_a_bits_corrupt = buffer_nodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_b_ready = buffer_nodeIn_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_auto_in_b_valid = buffer_nodeIn_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_opcode = buffer_nodeIn_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_param = buffer_nodeIn_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_size = buffer_nodeIn_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_source = buffer_nodeIn_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_address = buffer_nodeIn_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_mask = buffer_nodeIn_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_data = buffer_nodeIn_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_b_bits_corrupt = buffer_nodeIn_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_c_ready = buffer_nodeIn_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeOut_c_valid = buffer_nodeIn_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_opcode = buffer_nodeIn_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_param = buffer_nodeIn_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_size = buffer_nodeIn_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_source = buffer_nodeIn_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_address = buffer_nodeIn_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_bufferable =
    buffer_nodeIn_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_modifiable =
    buffer_nodeIn_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_readalloc =
    buffer_nodeIn_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_writealloc =
    buffer_nodeIn_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_privileged =
    buffer_nodeIn_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_secure =
    buffer_nodeIn_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_user_amba_prot_fetch =
    buffer_nodeIn_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_data = buffer_nodeIn_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_c_bits_corrupt = buffer_nodeIn_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_d_ready = buffer_nodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_auto_in_d_valid = buffer_nodeIn_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_opcode = buffer_nodeIn_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_param = buffer_nodeIn_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_size = buffer_nodeIn_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_source = buffer_nodeIn_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_sink = buffer_nodeIn_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_denied = buffer_nodeIn_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_data = buffer_nodeIn_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_d_bits_corrupt = buffer_nodeIn_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_auto_in_e_ready = buffer_nodeIn_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1214:17
  assign buffer_nodeOut_e_valid = buffer_nodeIn_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_nodeOut_e_bits_sink = buffer_nodeIn_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_a_ready = tlOtherMastersNodeOut_a_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_auto_in_a_valid = tlOtherMastersNodeOut_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_opcode = tlOtherMastersNodeOut_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_param = tlOtherMastersNodeOut_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_size = tlOtherMastersNodeOut_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_source = tlOtherMastersNodeOut_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_address = tlOtherMastersNodeOut_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_bufferable =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_modifiable =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_readalloc =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_writealloc =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_privileged =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_secure =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_user_amba_prot_fetch =
    tlOtherMastersNodeOut_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_mask = tlOtherMastersNodeOut_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_data = tlOtherMastersNodeOut_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_a_bits_corrupt = tlOtherMastersNodeOut_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_b_ready = tlOtherMastersNodeOut_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign tlOtherMastersNodeIn_b_valid = tlOtherMastersNodeOut_b_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_opcode = tlOtherMastersNodeOut_b_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_param = tlOtherMastersNodeOut_b_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_size = tlOtherMastersNodeOut_b_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_source = tlOtherMastersNodeOut_b_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_address = tlOtherMastersNodeOut_b_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_mask = tlOtherMastersNodeOut_b_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_data = tlOtherMastersNodeOut_b_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_b_bits_corrupt = tlOtherMastersNodeOut_b_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_c_ready = tlOtherMastersNodeOut_c_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_auto_in_c_valid = tlOtherMastersNodeOut_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_opcode = tlOtherMastersNodeOut_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_param = tlOtherMastersNodeOut_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_size = tlOtherMastersNodeOut_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_source = tlOtherMastersNodeOut_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_address = tlOtherMastersNodeOut_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_bufferable =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_modifiable =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_readalloc =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_writealloc =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_privileged =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_secure =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_user_amba_prot_fetch =
    tlOtherMastersNodeOut_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_data = tlOtherMastersNodeOut_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_c_bits_corrupt = tlOtherMastersNodeOut_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_d_ready = tlOtherMastersNodeOut_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign tlOtherMastersNodeIn_d_valid = tlOtherMastersNodeOut_d_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_opcode = tlOtherMastersNodeOut_d_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_param = tlOtherMastersNodeOut_d_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_size = tlOtherMastersNodeOut_d_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_source = tlOtherMastersNodeOut_d_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_sink = tlOtherMastersNodeOut_d_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_denied = tlOtherMastersNodeOut_d_bits_denied;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_data = tlOtherMastersNodeOut_d_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_d_bits_corrupt = tlOtherMastersNodeOut_d_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeIn_e_ready = tlOtherMastersNodeOut_e_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign buffer_auto_in_e_valid = tlOtherMastersNodeOut_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign buffer_auto_in_e_bits_sink = tlOtherMastersNodeOut_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign tlOtherMastersNodeOut_a_valid = tlOtherMastersNodeIn_a_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_opcode = tlOtherMastersNodeIn_a_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_param = tlOtherMastersNodeIn_a_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_size = tlOtherMastersNodeIn_a_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_source = tlOtherMastersNodeIn_a_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_address = tlOtherMastersNodeIn_a_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_bufferable =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_modifiable =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_readalloc =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_writealloc =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_privileged =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_secure =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_user_amba_prot_fetch =
    tlOtherMastersNodeIn_a_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_mask = tlOtherMastersNodeIn_a_bits_mask;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_data = tlOtherMastersNodeIn_a_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_a_bits_corrupt = tlOtherMastersNodeIn_a_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_b_ready = tlOtherMastersNodeIn_b_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_valid = tlOtherMastersNodeIn_c_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_opcode = tlOtherMastersNodeIn_c_bits_opcode;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_param = tlOtherMastersNodeIn_c_bits_param;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_size = tlOtherMastersNodeIn_c_bits_size;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_source = tlOtherMastersNodeIn_c_bits_source;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_address = tlOtherMastersNodeIn_c_bits_address;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_bufferable =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_bufferable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_modifiable =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_modifiable;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_readalloc =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_readalloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_writealloc =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_writealloc;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_privileged =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_privileged;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_secure =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_secure;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_user_amba_prot_fetch =
    tlOtherMastersNodeIn_c_bits_user_amba_prot_fetch;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_data = tlOtherMastersNodeIn_c_bits_data;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_c_bits_corrupt = tlOtherMastersNodeIn_c_bits_corrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_d_ready = tlOtherMastersNodeIn_d_ready;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_e_valid = tlOtherMastersNodeIn_e_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign tlOtherMastersNodeOut_e_bits_sink = tlOtherMastersNodeIn_e_bits_sink;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_auto_in = hartidOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign hartidOut = hartidIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_1_auto_in = reset_vectorOut;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign reset_vectorOut = reset_vectorIn;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_2_auto_in_rnmi = nmiOut_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_2_auto_in_rnmi_interrupt_vector = nmiOut_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_2_auto_in_rnmi_exception_vector = nmiOut_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign nmiOut_rnmi = nmiIn_rnmi;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign nmiOut_rnmi_interrupt_vector = nmiIn_rnmi_interrupt_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign nmiOut_rnmi_exception_vector = nmiIn_rnmi_exception_vector;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign broadcast_3_auto_in_insns_0_valid = traceSourceNodeOut_insns_0_valid;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_iaddr = traceSourceNodeOut_insns_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_insn = traceSourceNodeOut_insns_0_insn;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_priv = traceSourceNodeOut_insns_0_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_exception = traceSourceNodeOut_insns_0_exception;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_interrupt = traceSourceNodeOut_insns_0_interrupt;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_cause = traceSourceNodeOut_insns_0_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_insns_0_tval = traceSourceNodeOut_insns_0_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_3_auto_in_time = traceSourceNodeOut_time;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_4_auto_in_0_valid_0 = bpwatchSourceNodeOut_0_valid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_4_auto_in_0_rvalid_0 = bpwatchSourceNodeOut_0_rvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_4_auto_in_0_wvalid_0 = bpwatchSourceNodeOut_0_wvalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_4_auto_in_0_ivalid_0 = bpwatchSourceNodeOut_0_ivalid_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign broadcast_4_auto_in_0_action = bpwatchSourceNodeOut_0_action;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign int_localOut_0 = int_localIn_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign x1_int_localOut_0 = x1_int_localIn_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign x1_int_localOut_1 = x1_int_localIn_1;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  assign x1_int_localOut_1_0 = x1_int_localIn_1_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17, :1214:17
  wire dcacheArb_clock;
    wire dcacheArb_reset;
    wire dcacheArb_io_requestor_0_req_ready;
    wire dcacheArb_io_requestor_0_req_valid;
    wire[33:0] dcacheArb_io_requestor_0_req_bits_addr;
    wire[5:0] dcacheArb_io_requestor_0_req_bits_tag;
    wire[4:0] dcacheArb_io_requestor_0_req_bits_cmd;
    wire[1:0] dcacheArb_io_requestor_0_req_bits_size;
    wire dcacheArb_io_requestor_0_req_bits_signed;
    wire[1:0] dcacheArb_io_requestor_0_req_bits_dprv;
    wire dcacheArb_io_requestor_0_req_bits_dv;
    wire dcacheArb_io_requestor_0_req_bits_phys;
    wire dcacheArb_io_requestor_0_req_bits_no_alloc;
    wire dcacheArb_io_requestor_0_req_bits_no_xcpt;
    wire[63:0] dcacheArb_io_requestor_0_req_bits_data;
    wire[7:0] dcacheArb_io_requestor_0_req_bits_mask;
    wire dcacheArb_io_requestor_0_s1_kill;
    wire[63:0] dcacheArb_io_requestor_0_s1_data_data;
    wire[7:0] dcacheArb_io_requestor_0_s1_data_mask;
    wire dcacheArb_io_requestor_0_s2_nack;
    wire dcacheArb_io_requestor_0_s2_nack_cause_raw;
    wire dcacheArb_io_requestor_0_s2_kill;
    wire dcacheArb_io_requestor_0_s2_uncached;
    wire[31:0] dcacheArb_io_requestor_0_s2_paddr;
    wire dcacheArb_io_requestor_0_resp_valid;
    wire[33:0] dcacheArb_io_requestor_0_resp_bits_addr;
    wire[5:0] dcacheArb_io_requestor_0_resp_bits_tag;
    wire[4:0] dcacheArb_io_requestor_0_resp_bits_cmd;
    wire[1:0] dcacheArb_io_requestor_0_resp_bits_size;
    wire dcacheArb_io_requestor_0_resp_bits_signed;
    wire[1:0] dcacheArb_io_requestor_0_resp_bits_dprv;
    wire dcacheArb_io_requestor_0_resp_bits_dv;
    wire[63:0] dcacheArb_io_requestor_0_resp_bits_data;
    wire[7:0] dcacheArb_io_requestor_0_resp_bits_mask;
    wire dcacheArb_io_requestor_0_resp_bits_replay;
    wire dcacheArb_io_requestor_0_resp_bits_has_data;
    wire[63:0] dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    wire[63:0] dcacheArb_io_requestor_0_resp_bits_data_raw;
    wire[63:0] dcacheArb_io_requestor_0_resp_bits_store_data;
    wire dcacheArb_io_requestor_0_replay_next;
    wire dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    wire dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    wire dcacheArb_io_requestor_0_s2_xcpt_gf_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_gf_st;
    wire dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    wire dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    wire[33:0] dcacheArb_io_requestor_0_s2_gpa;
    wire dcacheArb_io_requestor_0_s2_gpa_is_pte;
    wire dcacheArb_io_requestor_0_ordered;
    wire dcacheArb_io_requestor_0_perf_acquire;
    wire dcacheArb_io_requestor_0_perf_release;
    wire dcacheArb_io_requestor_0_perf_grant;
    wire dcacheArb_io_requestor_0_perf_tlbMiss;
    wire dcacheArb_io_requestor_0_perf_blocked;
    wire dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad;
    wire dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW;
    wire dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad;
    wire dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad;
    wire dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore;
    wire dcacheArb_io_requestor_0_keep_clock_enabled;
    wire dcacheArb_io_requestor_0_clock_enabled;
    wire dcacheArb_io_mem_req_ready;
    wire dcacheArb_io_mem_req_valid;
    wire[33:0] dcacheArb_io_mem_req_bits_addr;
    wire[5:0] dcacheArb_io_mem_req_bits_tag;
    wire[4:0] dcacheArb_io_mem_req_bits_cmd;
    wire[1:0] dcacheArb_io_mem_req_bits_size;
    wire dcacheArb_io_mem_req_bits_signed;
    wire[1:0] dcacheArb_io_mem_req_bits_dprv;
    wire dcacheArb_io_mem_req_bits_dv;
    wire dcacheArb_io_mem_req_bits_phys;
    wire dcacheArb_io_mem_req_bits_no_alloc;
    wire dcacheArb_io_mem_req_bits_no_xcpt;
    wire[63:0] dcacheArb_io_mem_req_bits_data;
    wire[7:0] dcacheArb_io_mem_req_bits_mask;
    wire dcacheArb_io_mem_s1_kill;
    wire[63:0] dcacheArb_io_mem_s1_data_data;
    wire[7:0] dcacheArb_io_mem_s1_data_mask;
    wire dcacheArb_io_mem_s2_nack;
    wire dcacheArb_io_mem_s2_nack_cause_raw;
    wire dcacheArb_io_mem_s2_kill;
    wire dcacheArb_io_mem_s2_uncached;
    wire[31:0] dcacheArb_io_mem_s2_paddr;
    wire dcacheArb_io_mem_resp_valid;
    wire[33:0] dcacheArb_io_mem_resp_bits_addr;
    wire[5:0] dcacheArb_io_mem_resp_bits_tag;
    wire[4:0] dcacheArb_io_mem_resp_bits_cmd;
    wire[1:0] dcacheArb_io_mem_resp_bits_size;
    wire dcacheArb_io_mem_resp_bits_signed;
    wire[1:0] dcacheArb_io_mem_resp_bits_dprv;
    wire dcacheArb_io_mem_resp_bits_dv;
    wire[63:0] dcacheArb_io_mem_resp_bits_data;
    wire[7:0] dcacheArb_io_mem_resp_bits_mask;
    wire dcacheArb_io_mem_resp_bits_replay;
    wire dcacheArb_io_mem_resp_bits_has_data;
    wire[63:0] dcacheArb_io_mem_resp_bits_data_word_bypass;
    wire[63:0] dcacheArb_io_mem_resp_bits_data_raw;
    wire[63:0] dcacheArb_io_mem_resp_bits_store_data;
    wire dcacheArb_io_mem_replay_next;
    wire dcacheArb_io_mem_s2_xcpt_ma_ld;
    wire dcacheArb_io_mem_s2_xcpt_ma_st;
    wire dcacheArb_io_mem_s2_xcpt_pf_ld;
    wire dcacheArb_io_mem_s2_xcpt_pf_st;
    wire dcacheArb_io_mem_s2_xcpt_gf_ld;
    wire dcacheArb_io_mem_s2_xcpt_gf_st;
    wire dcacheArb_io_mem_s2_xcpt_ae_ld;
    wire dcacheArb_io_mem_s2_xcpt_ae_st;
    wire[33:0] dcacheArb_io_mem_s2_gpa;
    wire dcacheArb_io_mem_s2_gpa_is_pte;
    wire dcacheArb_io_mem_ordered;
    wire dcacheArb_io_mem_perf_acquire;
    wire dcacheArb_io_mem_perf_release;
    wire dcacheArb_io_mem_perf_grant;
    wire dcacheArb_io_mem_perf_tlbMiss;
    wire dcacheArb_io_mem_perf_blocked;
    wire dcacheArb_io_mem_perf_canAcceptStoreThenLoad;
    wire dcacheArb_io_mem_perf_canAcceptStoreThenRMW;
    wire dcacheArb_io_mem_perf_canAcceptLoadThenLoad;
    wire dcacheArb_io_mem_perf_storeBufferEmptyAfterLoad;
    wire dcacheArb_io_mem_perf_storeBufferEmptyAfterStore;
    wire dcacheArb_io_mem_keep_clock_enabled;
    wire dcacheArb_io_mem_clock_enabled;

    assign  dcacheArb_io_requestor_0_req_ready = dcacheArb_io_mem_req_ready ; 
  assign  dcacheArb_io_requestor_0_s2_nack = dcacheArb_io_mem_s2_nack ; 
  assign  dcacheArb_io_requestor_0_s2_nack_cause_raw = dcacheArb_io_mem_s2_nack_cause_raw ; 
  assign  dcacheArb_io_requestor_0_s2_uncached = dcacheArb_io_mem_s2_uncached ; 
  assign  dcacheArb_io_requestor_0_s2_paddr = dcacheArb_io_mem_s2_paddr ; 
  assign  dcacheArb_io_requestor_0_resp_valid = dcacheArb_io_mem_resp_valid ; 
  assign  dcacheArb_io_requestor_0_resp_bits_addr = dcacheArb_io_mem_resp_bits_addr ; 
  assign  dcacheArb_io_requestor_0_resp_bits_tag = dcacheArb_io_mem_resp_bits_tag ; 
  assign  dcacheArb_io_requestor_0_resp_bits_cmd = dcacheArb_io_mem_resp_bits_cmd ; 
  assign  dcacheArb_io_requestor_0_resp_bits_size = dcacheArb_io_mem_resp_bits_size ; 
  assign  dcacheArb_io_requestor_0_resp_bits_signed = dcacheArb_io_mem_resp_bits_signed ; 
  assign  dcacheArb_io_requestor_0_resp_bits_dprv = dcacheArb_io_mem_resp_bits_dprv ; 
  assign  dcacheArb_io_requestor_0_resp_bits_dv = dcacheArb_io_mem_resp_bits_dv ; 
  assign  dcacheArb_io_requestor_0_resp_bits_data = dcacheArb_io_mem_resp_bits_data ; 
  assign  dcacheArb_io_requestor_0_resp_bits_mask = dcacheArb_io_mem_resp_bits_mask ; 
  assign  dcacheArb_io_requestor_0_resp_bits_replay = dcacheArb_io_mem_resp_bits_replay ; 
  assign  dcacheArb_io_requestor_0_resp_bits_has_data = dcacheArb_io_mem_resp_bits_has_data ; 
  assign  dcacheArb_io_requestor_0_resp_bits_data_word_bypass = dcacheArb_io_mem_resp_bits_data_word_bypass ; 
  assign  dcacheArb_io_requestor_0_resp_bits_data_raw = dcacheArb_io_mem_resp_bits_data_raw ; 
  assign  dcacheArb_io_requestor_0_resp_bits_store_data = dcacheArb_io_mem_resp_bits_store_data ; 
  assign  dcacheArb_io_requestor_0_replay_next = dcacheArb_io_mem_replay_next ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ma_ld = dcacheArb_io_mem_s2_xcpt_ma_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ma_st = dcacheArb_io_mem_s2_xcpt_ma_st ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_pf_ld = dcacheArb_io_mem_s2_xcpt_pf_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_pf_st = dcacheArb_io_mem_s2_xcpt_pf_st ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_gf_ld = dcacheArb_io_mem_s2_xcpt_gf_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_gf_st = dcacheArb_io_mem_s2_xcpt_gf_st ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ae_ld = dcacheArb_io_mem_s2_xcpt_ae_ld ; 
  assign  dcacheArb_io_requestor_0_s2_xcpt_ae_st = dcacheArb_io_mem_s2_xcpt_ae_st ; 
  assign  dcacheArb_io_requestor_0_s2_gpa = dcacheArb_io_mem_s2_gpa ; 
  assign  dcacheArb_io_requestor_0_s2_gpa_is_pte = dcacheArb_io_mem_s2_gpa_is_pte ; 
  assign  dcacheArb_io_requestor_0_ordered = dcacheArb_io_mem_ordered ; 
  assign  dcacheArb_io_requestor_0_perf_acquire = dcacheArb_io_mem_perf_acquire ; 
  assign  dcacheArb_io_requestor_0_perf_release = dcacheArb_io_mem_perf_release ; 
  assign  dcacheArb_io_requestor_0_perf_grant = dcacheArb_io_mem_perf_grant ; 
  assign  dcacheArb_io_requestor_0_perf_tlbMiss = dcacheArb_io_mem_perf_tlbMiss ; 
  assign  dcacheArb_io_requestor_0_perf_blocked = dcacheArb_io_mem_perf_blocked ; 
  assign  dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad = dcacheArb_io_mem_perf_canAcceptStoreThenLoad ; 
  assign  dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW = dcacheArb_io_mem_perf_canAcceptStoreThenRMW ; 
  assign  dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad = dcacheArb_io_mem_perf_canAcceptLoadThenLoad ; 
  assign  dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad = dcacheArb_io_mem_perf_storeBufferEmptyAfterLoad ; 
  assign  dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore = dcacheArb_io_mem_perf_storeBufferEmptyAfterStore ; 
  assign  dcacheArb_io_requestor_0_clock_enabled = dcacheArb_io_mem_clock_enabled ; 
  assign  dcacheArb_io_mem_req_valid = dcacheArb_io_requestor_0_req_valid ; 
  assign  dcacheArb_io_mem_req_bits_addr = dcacheArb_io_requestor_0_req_bits_addr ; 
  assign  dcacheArb_io_mem_req_bits_tag = dcacheArb_io_requestor_0_req_bits_tag ; 
  assign  dcacheArb_io_mem_req_bits_cmd = dcacheArb_io_requestor_0_req_bits_cmd ; 
  assign  dcacheArb_io_mem_req_bits_size = dcacheArb_io_requestor_0_req_bits_size ; 
  assign  dcacheArb_io_mem_req_bits_signed = dcacheArb_io_requestor_0_req_bits_signed ; 
  assign  dcacheArb_io_mem_req_bits_dprv = dcacheArb_io_requestor_0_req_bits_dprv ; 
  assign  dcacheArb_io_mem_req_bits_dv = dcacheArb_io_requestor_0_req_bits_dv ; 
  assign  dcacheArb_io_mem_req_bits_phys = dcacheArb_io_requestor_0_req_bits_phys ; 
  assign  dcacheArb_io_mem_req_bits_no_alloc = dcacheArb_io_requestor_0_req_bits_no_alloc ; 
  assign  dcacheArb_io_mem_req_bits_no_xcpt = dcacheArb_io_requestor_0_req_bits_no_xcpt ; 
  assign  dcacheArb_io_mem_req_bits_data = dcacheArb_io_requestor_0_req_bits_data ; 
  assign  dcacheArb_io_mem_req_bits_mask = dcacheArb_io_requestor_0_req_bits_mask ; 
  assign  dcacheArb_io_mem_s1_kill = dcacheArb_io_requestor_0_s1_kill ; 
  assign  dcacheArb_io_mem_s1_data_data = dcacheArb_io_requestor_0_s1_data_data ; 
  assign  dcacheArb_io_mem_s1_data_mask = dcacheArb_io_requestor_0_s1_data_mask ; 
  assign  dcacheArb_io_mem_s2_kill = dcacheArb_io_requestor_0_s2_kill ; 
  assign  dcacheArb_io_mem_keep_clock_enabled = dcacheArb_io_requestor_0_keep_clock_enabled ;
    assign dcacheArb_clock = clock;
    assign dcacheArb_reset = reset;
    assign _dcacheArb_io_requestor_0_req_ready = dcacheArb_io_requestor_0_req_ready;
    assign dcacheArb_io_requestor_0_req_valid = _core_io_dmem_req_valid;
    assign dcacheArb_io_requestor_0_req_bits_addr = _core_io_dmem_req_bits_addr;
    assign dcacheArb_io_requestor_0_req_bits_tag = _core_io_dmem_req_bits_tag;
    assign dcacheArb_io_requestor_0_req_bits_cmd = _core_io_dmem_req_bits_cmd;
    assign dcacheArb_io_requestor_0_req_bits_size = _core_io_dmem_req_bits_size;
    assign dcacheArb_io_requestor_0_req_bits_signed = _core_io_dmem_req_bits_signed;
    assign dcacheArb_io_requestor_0_req_bits_dprv = _core_io_dmem_req_bits_dprv;
    assign dcacheArb_io_requestor_0_req_bits_dv = _core_io_dmem_req_bits_dv;
    assign dcacheArb_io_requestor_0_req_bits_phys = _core_io_dmem_req_bits_phys;
    assign dcacheArb_io_requestor_0_req_bits_no_alloc = _core_io_dmem_req_bits_no_alloc;
    assign dcacheArb_io_requestor_0_req_bits_no_xcpt = _core_io_dmem_req_bits_no_xcpt;
    assign dcacheArb_io_requestor_0_req_bits_data = _core_io_dmem_req_bits_data;
    assign dcacheArb_io_requestor_0_req_bits_mask = _core_io_dmem_req_bits_mask;
    assign dcacheArb_io_requestor_0_s1_kill = _core_io_dmem_s1_kill;
    assign dcacheArb_io_requestor_0_s1_data_data = _core_io_dmem_s1_data_data;
    assign dcacheArb_io_requestor_0_s1_data_mask = _core_io_dmem_s1_data_mask;
    assign _dcacheArb_io_requestor_0_s2_nack = dcacheArb_io_requestor_0_s2_nack;
    assign _dcacheArb_io_requestor_0_s2_nack_cause_raw = dcacheArb_io_requestor_0_s2_nack_cause_raw;
    assign dcacheArb_io_requestor_0_s2_kill = _core_io_dmem_s2_kill;
    assign _dcacheArb_io_requestor_0_s2_uncached = dcacheArb_io_requestor_0_s2_uncached;
    assign _dcacheArb_io_requestor_0_s2_paddr = dcacheArb_io_requestor_0_s2_paddr;
    assign _dcacheArb_io_requestor_0_resp_valid = dcacheArb_io_requestor_0_resp_valid;
    assign _dcacheArb_io_requestor_0_resp_bits_addr = dcacheArb_io_requestor_0_resp_bits_addr;
    assign _dcacheArb_io_requestor_0_resp_bits_tag = dcacheArb_io_requestor_0_resp_bits_tag;
    assign _dcacheArb_io_requestor_0_resp_bits_cmd = dcacheArb_io_requestor_0_resp_bits_cmd;
    assign _dcacheArb_io_requestor_0_resp_bits_size = dcacheArb_io_requestor_0_resp_bits_size;
    assign _dcacheArb_io_requestor_0_resp_bits_signed = dcacheArb_io_requestor_0_resp_bits_signed;
    assign _dcacheArb_io_requestor_0_resp_bits_dprv = dcacheArb_io_requestor_0_resp_bits_dprv;
    assign _dcacheArb_io_requestor_0_resp_bits_dv = dcacheArb_io_requestor_0_resp_bits_dv;
    assign _dcacheArb_io_requestor_0_resp_bits_data = dcacheArb_io_requestor_0_resp_bits_data;
    assign _dcacheArb_io_requestor_0_resp_bits_mask = dcacheArb_io_requestor_0_resp_bits_mask;
    assign _dcacheArb_io_requestor_0_resp_bits_replay = dcacheArb_io_requestor_0_resp_bits_replay;
    assign _dcacheArb_io_requestor_0_resp_bits_has_data = dcacheArb_io_requestor_0_resp_bits_has_data;
    assign _dcacheArb_io_requestor_0_resp_bits_data_word_bypass = dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    assign _dcacheArb_io_requestor_0_resp_bits_data_raw = dcacheArb_io_requestor_0_resp_bits_data_raw;
    assign _dcacheArb_io_requestor_0_resp_bits_store_data = dcacheArb_io_requestor_0_resp_bits_store_data;
    assign _dcacheArb_io_requestor_0_replay_next = dcacheArb_io_requestor_0_replay_next;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ma_ld = dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ma_st = dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    assign _dcacheArb_io_requestor_0_s2_xcpt_pf_ld = dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_pf_st = dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    assign _dcacheArb_io_requestor_0_s2_xcpt_gf_ld = dcacheArb_io_requestor_0_s2_xcpt_gf_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_gf_st = dcacheArb_io_requestor_0_s2_xcpt_gf_st;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ae_ld = dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    assign _dcacheArb_io_requestor_0_s2_xcpt_ae_st = dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    assign _dcacheArb_io_requestor_0_s2_gpa = dcacheArb_io_requestor_0_s2_gpa;
    assign _dcacheArb_io_requestor_0_s2_gpa_is_pte = dcacheArb_io_requestor_0_s2_gpa_is_pte;
    assign _dcacheArb_io_requestor_0_ordered = dcacheArb_io_requestor_0_ordered;
    assign _dcacheArb_io_requestor_0_perf_acquire = dcacheArb_io_requestor_0_perf_acquire;
    assign _dcacheArb_io_requestor_0_perf_release = dcacheArb_io_requestor_0_perf_release;
    assign _dcacheArb_io_requestor_0_perf_grant = dcacheArb_io_requestor_0_perf_grant;
    assign _dcacheArb_io_requestor_0_perf_tlbMiss = dcacheArb_io_requestor_0_perf_tlbMiss;
    assign _dcacheArb_io_requestor_0_perf_blocked = dcacheArb_io_requestor_0_perf_blocked;
    assign _dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad = dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad;
    assign _dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW = dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW;
    assign _dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad = dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad;
    assign _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad = dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad;
    assign _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore = dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore;
    assign dcacheArb_io_requestor_0_keep_clock_enabled = _core_io_dmem_keep_clock_enabled;
    assign _dcacheArb_io_requestor_0_clock_enabled = dcacheArb_io_requestor_0_clock_enabled;
    assign dcacheArb_io_mem_req_ready = _dcache_io_cpu_req_ready;
    assign _dcacheArb_io_mem_req_valid = dcacheArb_io_mem_req_valid;
    assign _dcacheArb_io_mem_req_bits_addr = dcacheArb_io_mem_req_bits_addr;
    assign _dcacheArb_io_mem_req_bits_tag = dcacheArb_io_mem_req_bits_tag;
    assign _dcacheArb_io_mem_req_bits_cmd = dcacheArb_io_mem_req_bits_cmd;
    assign _dcacheArb_io_mem_req_bits_size = dcacheArb_io_mem_req_bits_size;
    assign _dcacheArb_io_mem_req_bits_signed = dcacheArb_io_mem_req_bits_signed;
    assign _dcacheArb_io_mem_req_bits_dprv = dcacheArb_io_mem_req_bits_dprv;
    assign _dcacheArb_io_mem_req_bits_dv = dcacheArb_io_mem_req_bits_dv;
    assign _dcacheArb_io_mem_req_bits_phys = dcacheArb_io_mem_req_bits_phys;
    assign _dcacheArb_io_mem_req_bits_no_alloc = dcacheArb_io_mem_req_bits_no_alloc;
    assign _dcacheArb_io_mem_req_bits_no_xcpt = dcacheArb_io_mem_req_bits_no_xcpt;
    assign _dcacheArb_io_mem_req_bits_data = dcacheArb_io_mem_req_bits_data;
    assign _dcacheArb_io_mem_req_bits_mask = dcacheArb_io_mem_req_bits_mask;
    assign _dcacheArb_io_mem_s1_kill = dcacheArb_io_mem_s1_kill;
    assign _dcacheArb_io_mem_s1_data_data = dcacheArb_io_mem_s1_data_data;
    assign _dcacheArb_io_mem_s1_data_mask = dcacheArb_io_mem_s1_data_mask;
    assign dcacheArb_io_mem_s2_nack = _dcache_io_cpu_s2_nack;
    assign dcacheArb_io_mem_s2_nack_cause_raw = _dcache_io_cpu_s2_nack_cause_raw;
    assign _dcacheArb_io_mem_s2_kill = dcacheArb_io_mem_s2_kill;
    assign dcacheArb_io_mem_s2_uncached = _dcache_io_cpu_s2_uncached;
    assign dcacheArb_io_mem_s2_paddr = _dcache_io_cpu_s2_paddr;
    assign dcacheArb_io_mem_resp_valid = _dcache_io_cpu_resp_valid;
    assign dcacheArb_io_mem_resp_bits_addr = _dcache_io_cpu_resp_bits_addr;
    assign dcacheArb_io_mem_resp_bits_tag = _dcache_io_cpu_resp_bits_tag;
    assign dcacheArb_io_mem_resp_bits_cmd = _dcache_io_cpu_resp_bits_cmd;
    assign dcacheArb_io_mem_resp_bits_size = _dcache_io_cpu_resp_bits_size;
    assign dcacheArb_io_mem_resp_bits_signed = _dcache_io_cpu_resp_bits_signed;
    assign dcacheArb_io_mem_resp_bits_dprv = _dcache_io_cpu_resp_bits_dprv;
    assign dcacheArb_io_mem_resp_bits_dv = _dcache_io_cpu_resp_bits_dv;
    assign dcacheArb_io_mem_resp_bits_data = _dcache_io_cpu_resp_bits_data;
    assign dcacheArb_io_mem_resp_bits_mask = _dcache_io_cpu_resp_bits_mask;
    assign dcacheArb_io_mem_resp_bits_replay = _dcache_io_cpu_resp_bits_replay;
    assign dcacheArb_io_mem_resp_bits_has_data = _dcache_io_cpu_resp_bits_has_data;
    assign dcacheArb_io_mem_resp_bits_data_word_bypass = _dcache_io_cpu_resp_bits_data_word_bypass;
    assign dcacheArb_io_mem_resp_bits_data_raw = _dcache_io_cpu_resp_bits_data_raw;
    assign dcacheArb_io_mem_resp_bits_store_data = _dcache_io_cpu_resp_bits_store_data;
    assign dcacheArb_io_mem_replay_next = _dcache_io_cpu_replay_next;
    assign dcacheArb_io_mem_s2_xcpt_ma_ld = _dcache_io_cpu_s2_xcpt_ma_ld;
    assign dcacheArb_io_mem_s2_xcpt_ma_st = _dcache_io_cpu_s2_xcpt_ma_st;
    assign dcacheArb_io_mem_s2_xcpt_pf_ld = _dcache_io_cpu_s2_xcpt_pf_ld;
    assign dcacheArb_io_mem_s2_xcpt_pf_st = _dcache_io_cpu_s2_xcpt_pf_st;
    assign dcacheArb_io_mem_s2_xcpt_gf_ld = _dcache_io_cpu_s2_xcpt_gf_ld;
    assign dcacheArb_io_mem_s2_xcpt_gf_st = _dcache_io_cpu_s2_xcpt_gf_st;
    assign dcacheArb_io_mem_s2_xcpt_ae_ld = _dcache_io_cpu_s2_xcpt_ae_ld;
    assign dcacheArb_io_mem_s2_xcpt_ae_st = _dcache_io_cpu_s2_xcpt_ae_st;
    assign dcacheArb_io_mem_s2_gpa = _dcache_io_cpu_s2_gpa;
    assign dcacheArb_io_mem_s2_gpa_is_pte = _dcache_io_cpu_s2_gpa_is_pte;
    assign dcacheArb_io_mem_ordered = _dcache_io_cpu_ordered;
    assign dcacheArb_io_mem_perf_acquire = _dcache_io_cpu_perf_acquire;
    assign dcacheArb_io_mem_perf_release = _dcache_io_cpu_perf_release;
    assign dcacheArb_io_mem_perf_grant = _dcache_io_cpu_perf_grant;
    assign dcacheArb_io_mem_perf_tlbMiss = _dcache_io_cpu_perf_tlbMiss;
    assign dcacheArb_io_mem_perf_blocked = _dcache_io_cpu_perf_blocked;
    assign dcacheArb_io_mem_perf_canAcceptStoreThenLoad = _dcache_io_cpu_perf_canAcceptStoreThenLoad;
    assign dcacheArb_io_mem_perf_canAcceptStoreThenRMW = _dcache_io_cpu_perf_canAcceptStoreThenRMW;
    assign dcacheArb_io_mem_perf_canAcceptLoadThenLoad = _dcache_io_cpu_perf_canAcceptLoadThenLoad;
    assign dcacheArb_io_mem_perf_storeBufferEmptyAfterLoad = _dcache_io_cpu_perf_storeBufferEmptyAfterLoad;
    assign dcacheArb_io_mem_perf_storeBufferEmptyAfterStore = _dcache_io_cpu_perf_storeBufferEmptyAfterStore;
    assign _dcacheArb_io_mem_keep_clock_enabled = dcacheArb_io_mem_keep_clock_enabled;
    assign dcacheArb_io_mem_clock_enabled = _dcache_io_cpu_clock_enabled;
    
  wire ptw_clock;
    wire ptw_reset;
    wire ptw_io_requestor_0_req_ready;
    wire ptw_io_requestor_0_req_valid;
    wire ptw_io_requestor_0_req_bits_valid;
    wire[20:0] ptw_io_requestor_0_req_bits_bits_addr;
    wire ptw_io_requestor_0_req_bits_bits_need_gpa;
    wire ptw_io_requestor_0_req_bits_bits_vstage1;
    wire ptw_io_requestor_0_req_bits_bits_stage2;
    wire ptw_io_requestor_0_resp_valid;
    wire ptw_io_requestor_0_resp_bits_ae_ptw;
    wire ptw_io_requestor_0_resp_bits_ae_final;
    wire ptw_io_requestor_0_resp_bits_pf;
    wire ptw_io_requestor_0_resp_bits_gf;
    wire ptw_io_requestor_0_resp_bits_hr;
    wire ptw_io_requestor_0_resp_bits_hw;
    wire ptw_io_requestor_0_resp_bits_hx;
    wire[9:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_future;
    wire[43:0] ptw_io_requestor_0_resp_bits_pte_ppn;
    wire[1:0] ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
    wire ptw_io_requestor_0_resp_bits_pte_d;
    wire ptw_io_requestor_0_resp_bits_pte_a;
    wire ptw_io_requestor_0_resp_bits_pte_g;
    wire ptw_io_requestor_0_resp_bits_pte_u;
    wire ptw_io_requestor_0_resp_bits_pte_x;
    wire ptw_io_requestor_0_resp_bits_pte_w;
    wire ptw_io_requestor_0_resp_bits_pte_r;
    wire ptw_io_requestor_0_resp_bits_pte_v;
    wire[1:0] ptw_io_requestor_0_resp_bits_level;
    wire ptw_io_requestor_0_resp_bits_fragmented_superpage;
    wire ptw_io_requestor_0_resp_bits_homogeneous;
    wire ptw_io_requestor_0_resp_bits_gpa_valid;
    wire[32:0] ptw_io_requestor_0_resp_bits_gpa_bits;
    wire ptw_io_requestor_0_resp_bits_gpa_is_pte;
    wire[3:0] ptw_io_requestor_0_ptbr_mode;
    wire[15:0] ptw_io_requestor_0_ptbr_asid;
    wire[43:0] ptw_io_requestor_0_ptbr_ppn;
    wire[3:0] ptw_io_requestor_0_hgatp_mode;
    wire[15:0] ptw_io_requestor_0_hgatp_asid;
    wire[43:0] ptw_io_requestor_0_hgatp_ppn;
    wire[3:0] ptw_io_requestor_0_vsatp_mode;
    wire[15:0] ptw_io_requestor_0_vsatp_asid;
    wire[43:0] ptw_io_requestor_0_vsatp_ppn;
    wire ptw_io_requestor_0_status_debug;
    wire ptw_io_requestor_0_status_cease;
    wire ptw_io_requestor_0_status_wfi;
    wire[31:0] ptw_io_requestor_0_status_isa;
    wire[1:0] ptw_io_requestor_0_status_dprv;
    wire ptw_io_requestor_0_status_dv;
    wire[1:0] ptw_io_requestor_0_status_prv;
    wire ptw_io_requestor_0_status_v;
    wire ptw_io_requestor_0_status_sd;
    wire[22:0] ptw_io_requestor_0_status_zero2;
    wire ptw_io_requestor_0_status_mpv;
    wire ptw_io_requestor_0_status_gva;
    wire ptw_io_requestor_0_status_mbe;
    wire ptw_io_requestor_0_status_sbe;
    wire[1:0] ptw_io_requestor_0_status_sxl;
    wire[1:0] ptw_io_requestor_0_status_uxl;
    wire ptw_io_requestor_0_status_sd_rv32;
    wire[7:0] ptw_io_requestor_0_status_zero1;
    wire ptw_io_requestor_0_status_tsr;
    wire ptw_io_requestor_0_status_tw;
    wire ptw_io_requestor_0_status_tvm;
    wire ptw_io_requestor_0_status_mxr;
    wire ptw_io_requestor_0_status_sum;
    wire ptw_io_requestor_0_status_mprv;
    wire[1:0] ptw_io_requestor_0_status_xs;
    wire[1:0] ptw_io_requestor_0_status_fs;
    wire[1:0] ptw_io_requestor_0_status_mpp;
    wire[1:0] ptw_io_requestor_0_status_vs;
    wire ptw_io_requestor_0_status_spp;
    wire ptw_io_requestor_0_status_mpie;
    wire ptw_io_requestor_0_status_ube;
    wire ptw_io_requestor_0_status_spie;
    wire ptw_io_requestor_0_status_upie;
    wire ptw_io_requestor_0_status_mie;
    wire ptw_io_requestor_0_status_hie;
    wire ptw_io_requestor_0_status_sie;
    wire ptw_io_requestor_0_status_uie;
    wire[29:0] ptw_io_requestor_0_hstatus_zero6;
    wire[1:0] ptw_io_requestor_0_hstatus_vsxl;
    wire[8:0] ptw_io_requestor_0_hstatus_zero5;
    wire ptw_io_requestor_0_hstatus_vtsr;
    wire ptw_io_requestor_0_hstatus_vtw;
    wire ptw_io_requestor_0_hstatus_vtvm;
    wire[1:0] ptw_io_requestor_0_hstatus_zero3;
    wire[5:0] ptw_io_requestor_0_hstatus_vgein;
    wire[1:0] ptw_io_requestor_0_hstatus_zero2;
    wire ptw_io_requestor_0_hstatus_hu;
    wire ptw_io_requestor_0_hstatus_spvp;
    wire ptw_io_requestor_0_hstatus_spv;
    wire ptw_io_requestor_0_hstatus_gva;
    wire ptw_io_requestor_0_hstatus_vsbe;
    wire[4:0] ptw_io_requestor_0_hstatus_zero1;
    wire ptw_io_requestor_0_gstatus_debug;
    wire ptw_io_requestor_0_gstatus_cease;
    wire ptw_io_requestor_0_gstatus_wfi;
    wire[31:0] ptw_io_requestor_0_gstatus_isa;
    wire[1:0] ptw_io_requestor_0_gstatus_dprv;
    wire ptw_io_requestor_0_gstatus_dv;
    wire[1:0] ptw_io_requestor_0_gstatus_prv;
    wire ptw_io_requestor_0_gstatus_v;
    wire ptw_io_requestor_0_gstatus_sd;
    wire[22:0] ptw_io_requestor_0_gstatus_zero2;
    wire ptw_io_requestor_0_gstatus_mpv;
    wire ptw_io_requestor_0_gstatus_gva;
    wire ptw_io_requestor_0_gstatus_mbe;
    wire ptw_io_requestor_0_gstatus_sbe;
    wire[1:0] ptw_io_requestor_0_gstatus_sxl;
    wire[1:0] ptw_io_requestor_0_gstatus_uxl;
    wire ptw_io_requestor_0_gstatus_sd_rv32;
    wire[7:0] ptw_io_requestor_0_gstatus_zero1;
    wire ptw_io_requestor_0_gstatus_tsr;
    wire ptw_io_requestor_0_gstatus_tw;
    wire ptw_io_requestor_0_gstatus_tvm;
    wire ptw_io_requestor_0_gstatus_mxr;
    wire ptw_io_requestor_0_gstatus_sum;
    wire ptw_io_requestor_0_gstatus_mprv;
    wire[1:0] ptw_io_requestor_0_gstatus_xs;
    wire[1:0] ptw_io_requestor_0_gstatus_fs;
    wire[1:0] ptw_io_requestor_0_gstatus_mpp;
    wire[1:0] ptw_io_requestor_0_gstatus_vs;
    wire ptw_io_requestor_0_gstatus_spp;
    wire ptw_io_requestor_0_gstatus_mpie;
    wire ptw_io_requestor_0_gstatus_ube;
    wire ptw_io_requestor_0_gstatus_spie;
    wire ptw_io_requestor_0_gstatus_upie;
    wire ptw_io_requestor_0_gstatus_mie;
    wire ptw_io_requestor_0_gstatus_hie;
    wire ptw_io_requestor_0_gstatus_sie;
    wire ptw_io_requestor_0_gstatus_uie;
    wire ptw_io_requestor_0_pmp_0_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_0_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_0_cfg_a;
    wire ptw_io_requestor_0_pmp_0_cfg_x;
    wire ptw_io_requestor_0_pmp_0_cfg_w;
    wire ptw_io_requestor_0_pmp_0_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_0_addr;
    wire[31:0] ptw_io_requestor_0_pmp_0_mask;
    wire ptw_io_requestor_0_pmp_1_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_1_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_1_cfg_a;
    wire ptw_io_requestor_0_pmp_1_cfg_x;
    wire ptw_io_requestor_0_pmp_1_cfg_w;
    wire ptw_io_requestor_0_pmp_1_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_1_addr;
    wire[31:0] ptw_io_requestor_0_pmp_1_mask;
    wire ptw_io_requestor_0_pmp_2_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_2_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_2_cfg_a;
    wire ptw_io_requestor_0_pmp_2_cfg_x;
    wire ptw_io_requestor_0_pmp_2_cfg_w;
    wire ptw_io_requestor_0_pmp_2_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_2_addr;
    wire[31:0] ptw_io_requestor_0_pmp_2_mask;
    wire ptw_io_requestor_0_pmp_3_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_3_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_3_cfg_a;
    wire ptw_io_requestor_0_pmp_3_cfg_x;
    wire ptw_io_requestor_0_pmp_3_cfg_w;
    wire ptw_io_requestor_0_pmp_3_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_3_addr;
    wire[31:0] ptw_io_requestor_0_pmp_3_mask;
    wire ptw_io_requestor_0_pmp_4_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_4_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_4_cfg_a;
    wire ptw_io_requestor_0_pmp_4_cfg_x;
    wire ptw_io_requestor_0_pmp_4_cfg_w;
    wire ptw_io_requestor_0_pmp_4_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_4_addr;
    wire[31:0] ptw_io_requestor_0_pmp_4_mask;
    wire ptw_io_requestor_0_pmp_5_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_5_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_5_cfg_a;
    wire ptw_io_requestor_0_pmp_5_cfg_x;
    wire ptw_io_requestor_0_pmp_5_cfg_w;
    wire ptw_io_requestor_0_pmp_5_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_5_addr;
    wire[31:0] ptw_io_requestor_0_pmp_5_mask;
    wire ptw_io_requestor_0_pmp_6_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_6_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_6_cfg_a;
    wire ptw_io_requestor_0_pmp_6_cfg_x;
    wire ptw_io_requestor_0_pmp_6_cfg_w;
    wire ptw_io_requestor_0_pmp_6_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_6_addr;
    wire[31:0] ptw_io_requestor_0_pmp_6_mask;
    wire ptw_io_requestor_0_pmp_7_cfg_l;
    wire[1:0] ptw_io_requestor_0_pmp_7_cfg_res;
    wire[1:0] ptw_io_requestor_0_pmp_7_cfg_a;
    wire ptw_io_requestor_0_pmp_7_cfg_x;
    wire ptw_io_requestor_0_pmp_7_cfg_w;
    wire ptw_io_requestor_0_pmp_7_cfg_r;
    wire[29:0] ptw_io_requestor_0_pmp_7_addr;
    wire[31:0] ptw_io_requestor_0_pmp_7_mask;
    wire ptw_io_requestor_0_customCSRs_csrs_0_ren;
    wire ptw_io_requestor_0_customCSRs_csrs_0_wen;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_0_wdata;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_0_value;
    wire ptw_io_requestor_0_customCSRs_csrs_0_stall;
    wire ptw_io_requestor_0_customCSRs_csrs_0_set;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_0_sdata;
    wire ptw_io_requestor_0_customCSRs_csrs_1_ren;
    wire ptw_io_requestor_0_customCSRs_csrs_1_wen;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_1_wdata;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_1_value;
    wire ptw_io_requestor_0_customCSRs_csrs_1_stall;
    wire ptw_io_requestor_0_customCSRs_csrs_1_set;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_1_sdata;
    wire ptw_io_requestor_0_customCSRs_csrs_2_ren;
    wire ptw_io_requestor_0_customCSRs_csrs_2_wen;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_2_wdata;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_2_value;
    wire ptw_io_requestor_0_customCSRs_csrs_2_stall;
    wire ptw_io_requestor_0_customCSRs_csrs_2_set;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_2_sdata;
    wire ptw_io_requestor_0_customCSRs_csrs_3_ren;
    wire ptw_io_requestor_0_customCSRs_csrs_3_wen;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_3_wdata;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_3_value;
    wire ptw_io_requestor_0_customCSRs_csrs_3_stall;
    wire ptw_io_requestor_0_customCSRs_csrs_3_set;
    wire[63:0] ptw_io_requestor_0_customCSRs_csrs_3_sdata;
    wire ptw_io_requestor_1_req_ready;
    wire ptw_io_requestor_1_req_valid;
    wire ptw_io_requestor_1_req_bits_valid;
    wire[20:0] ptw_io_requestor_1_req_bits_bits_addr;
    wire ptw_io_requestor_1_req_bits_bits_need_gpa;
    wire ptw_io_requestor_1_req_bits_bits_vstage1;
    wire ptw_io_requestor_1_req_bits_bits_stage2;
    wire ptw_io_requestor_1_resp_valid;
    wire ptw_io_requestor_1_resp_bits_ae_ptw;
    wire ptw_io_requestor_1_resp_bits_ae_final;
    wire ptw_io_requestor_1_resp_bits_pf;
    wire ptw_io_requestor_1_resp_bits_gf;
    wire ptw_io_requestor_1_resp_bits_hr;
    wire ptw_io_requestor_1_resp_bits_hw;
    wire ptw_io_requestor_1_resp_bits_hx;
    wire[9:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_future;
    wire[43:0] ptw_io_requestor_1_resp_bits_pte_ppn;
    wire[1:0] ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
    wire ptw_io_requestor_1_resp_bits_pte_d;
    wire ptw_io_requestor_1_resp_bits_pte_a;
    wire ptw_io_requestor_1_resp_bits_pte_g;
    wire ptw_io_requestor_1_resp_bits_pte_u;
    wire ptw_io_requestor_1_resp_bits_pte_x;
    wire ptw_io_requestor_1_resp_bits_pte_w;
    wire ptw_io_requestor_1_resp_bits_pte_r;
    wire ptw_io_requestor_1_resp_bits_pte_v;
    wire[1:0] ptw_io_requestor_1_resp_bits_level;
    wire ptw_io_requestor_1_resp_bits_fragmented_superpage;
    wire ptw_io_requestor_1_resp_bits_homogeneous;
    wire ptw_io_requestor_1_resp_bits_gpa_valid;
    wire[32:0] ptw_io_requestor_1_resp_bits_gpa_bits;
    wire ptw_io_requestor_1_resp_bits_gpa_is_pte;
    wire[3:0] ptw_io_requestor_1_ptbr_mode;
    wire[15:0] ptw_io_requestor_1_ptbr_asid;
    wire[43:0] ptw_io_requestor_1_ptbr_ppn;
    wire[3:0] ptw_io_requestor_1_hgatp_mode;
    wire[15:0] ptw_io_requestor_1_hgatp_asid;
    wire[43:0] ptw_io_requestor_1_hgatp_ppn;
    wire[3:0] ptw_io_requestor_1_vsatp_mode;
    wire[15:0] ptw_io_requestor_1_vsatp_asid;
    wire[43:0] ptw_io_requestor_1_vsatp_ppn;
    wire ptw_io_requestor_1_status_debug;
    wire ptw_io_requestor_1_status_cease;
    wire ptw_io_requestor_1_status_wfi;
    wire[31:0] ptw_io_requestor_1_status_isa;
    wire[1:0] ptw_io_requestor_1_status_dprv;
    wire ptw_io_requestor_1_status_dv;
    wire[1:0] ptw_io_requestor_1_status_prv;
    wire ptw_io_requestor_1_status_v;
    wire ptw_io_requestor_1_status_sd;
    wire[22:0] ptw_io_requestor_1_status_zero2;
    wire ptw_io_requestor_1_status_mpv;
    wire ptw_io_requestor_1_status_gva;
    wire ptw_io_requestor_1_status_mbe;
    wire ptw_io_requestor_1_status_sbe;
    wire[1:0] ptw_io_requestor_1_status_sxl;
    wire[1:0] ptw_io_requestor_1_status_uxl;
    wire ptw_io_requestor_1_status_sd_rv32;
    wire[7:0] ptw_io_requestor_1_status_zero1;
    wire ptw_io_requestor_1_status_tsr;
    wire ptw_io_requestor_1_status_tw;
    wire ptw_io_requestor_1_status_tvm;
    wire ptw_io_requestor_1_status_mxr;
    wire ptw_io_requestor_1_status_sum;
    wire ptw_io_requestor_1_status_mprv;
    wire[1:0] ptw_io_requestor_1_status_xs;
    wire[1:0] ptw_io_requestor_1_status_fs;
    wire[1:0] ptw_io_requestor_1_status_mpp;
    wire[1:0] ptw_io_requestor_1_status_vs;
    wire ptw_io_requestor_1_status_spp;
    wire ptw_io_requestor_1_status_mpie;
    wire ptw_io_requestor_1_status_ube;
    wire ptw_io_requestor_1_status_spie;
    wire ptw_io_requestor_1_status_upie;
    wire ptw_io_requestor_1_status_mie;
    wire ptw_io_requestor_1_status_hie;
    wire ptw_io_requestor_1_status_sie;
    wire ptw_io_requestor_1_status_uie;
    wire[29:0] ptw_io_requestor_1_hstatus_zero6;
    wire[1:0] ptw_io_requestor_1_hstatus_vsxl;
    wire[8:0] ptw_io_requestor_1_hstatus_zero5;
    wire ptw_io_requestor_1_hstatus_vtsr;
    wire ptw_io_requestor_1_hstatus_vtw;
    wire ptw_io_requestor_1_hstatus_vtvm;
    wire[1:0] ptw_io_requestor_1_hstatus_zero3;
    wire[5:0] ptw_io_requestor_1_hstatus_vgein;
    wire[1:0] ptw_io_requestor_1_hstatus_zero2;
    wire ptw_io_requestor_1_hstatus_hu;
    wire ptw_io_requestor_1_hstatus_spvp;
    wire ptw_io_requestor_1_hstatus_spv;
    wire ptw_io_requestor_1_hstatus_gva;
    wire ptw_io_requestor_1_hstatus_vsbe;
    wire[4:0] ptw_io_requestor_1_hstatus_zero1;
    wire ptw_io_requestor_1_gstatus_debug;
    wire ptw_io_requestor_1_gstatus_cease;
    wire ptw_io_requestor_1_gstatus_wfi;
    wire[31:0] ptw_io_requestor_1_gstatus_isa;
    wire[1:0] ptw_io_requestor_1_gstatus_dprv;
    wire ptw_io_requestor_1_gstatus_dv;
    wire[1:0] ptw_io_requestor_1_gstatus_prv;
    wire ptw_io_requestor_1_gstatus_v;
    wire ptw_io_requestor_1_gstatus_sd;
    wire[22:0] ptw_io_requestor_1_gstatus_zero2;
    wire ptw_io_requestor_1_gstatus_mpv;
    wire ptw_io_requestor_1_gstatus_gva;
    wire ptw_io_requestor_1_gstatus_mbe;
    wire ptw_io_requestor_1_gstatus_sbe;
    wire[1:0] ptw_io_requestor_1_gstatus_sxl;
    wire[1:0] ptw_io_requestor_1_gstatus_uxl;
    wire ptw_io_requestor_1_gstatus_sd_rv32;
    wire[7:0] ptw_io_requestor_1_gstatus_zero1;
    wire ptw_io_requestor_1_gstatus_tsr;
    wire ptw_io_requestor_1_gstatus_tw;
    wire ptw_io_requestor_1_gstatus_tvm;
    wire ptw_io_requestor_1_gstatus_mxr;
    wire ptw_io_requestor_1_gstatus_sum;
    wire ptw_io_requestor_1_gstatus_mprv;
    wire[1:0] ptw_io_requestor_1_gstatus_xs;
    wire[1:0] ptw_io_requestor_1_gstatus_fs;
    wire[1:0] ptw_io_requestor_1_gstatus_mpp;
    wire[1:0] ptw_io_requestor_1_gstatus_vs;
    wire ptw_io_requestor_1_gstatus_spp;
    wire ptw_io_requestor_1_gstatus_mpie;
    wire ptw_io_requestor_1_gstatus_ube;
    wire ptw_io_requestor_1_gstatus_spie;
    wire ptw_io_requestor_1_gstatus_upie;
    wire ptw_io_requestor_1_gstatus_mie;
    wire ptw_io_requestor_1_gstatus_hie;
    wire ptw_io_requestor_1_gstatus_sie;
    wire ptw_io_requestor_1_gstatus_uie;
    wire ptw_io_requestor_1_pmp_0_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_0_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_0_cfg_a;
    wire ptw_io_requestor_1_pmp_0_cfg_x;
    wire ptw_io_requestor_1_pmp_0_cfg_w;
    wire ptw_io_requestor_1_pmp_0_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_0_addr;
    wire[31:0] ptw_io_requestor_1_pmp_0_mask;
    wire ptw_io_requestor_1_pmp_1_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_1_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_1_cfg_a;
    wire ptw_io_requestor_1_pmp_1_cfg_x;
    wire ptw_io_requestor_1_pmp_1_cfg_w;
    wire ptw_io_requestor_1_pmp_1_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_1_addr;
    wire[31:0] ptw_io_requestor_1_pmp_1_mask;
    wire ptw_io_requestor_1_pmp_2_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_2_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_2_cfg_a;
    wire ptw_io_requestor_1_pmp_2_cfg_x;
    wire ptw_io_requestor_1_pmp_2_cfg_w;
    wire ptw_io_requestor_1_pmp_2_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_2_addr;
    wire[31:0] ptw_io_requestor_1_pmp_2_mask;
    wire ptw_io_requestor_1_pmp_3_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_3_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_3_cfg_a;
    wire ptw_io_requestor_1_pmp_3_cfg_x;
    wire ptw_io_requestor_1_pmp_3_cfg_w;
    wire ptw_io_requestor_1_pmp_3_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_3_addr;
    wire[31:0] ptw_io_requestor_1_pmp_3_mask;
    wire ptw_io_requestor_1_pmp_4_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_4_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_4_cfg_a;
    wire ptw_io_requestor_1_pmp_4_cfg_x;
    wire ptw_io_requestor_1_pmp_4_cfg_w;
    wire ptw_io_requestor_1_pmp_4_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_4_addr;
    wire[31:0] ptw_io_requestor_1_pmp_4_mask;
    wire ptw_io_requestor_1_pmp_5_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_5_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_5_cfg_a;
    wire ptw_io_requestor_1_pmp_5_cfg_x;
    wire ptw_io_requestor_1_pmp_5_cfg_w;
    wire ptw_io_requestor_1_pmp_5_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_5_addr;
    wire[31:0] ptw_io_requestor_1_pmp_5_mask;
    wire ptw_io_requestor_1_pmp_6_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_6_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_6_cfg_a;
    wire ptw_io_requestor_1_pmp_6_cfg_x;
    wire ptw_io_requestor_1_pmp_6_cfg_w;
    wire ptw_io_requestor_1_pmp_6_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_6_addr;
    wire[31:0] ptw_io_requestor_1_pmp_6_mask;
    wire ptw_io_requestor_1_pmp_7_cfg_l;
    wire[1:0] ptw_io_requestor_1_pmp_7_cfg_res;
    wire[1:0] ptw_io_requestor_1_pmp_7_cfg_a;
    wire ptw_io_requestor_1_pmp_7_cfg_x;
    wire ptw_io_requestor_1_pmp_7_cfg_w;
    wire ptw_io_requestor_1_pmp_7_cfg_r;
    wire[29:0] ptw_io_requestor_1_pmp_7_addr;
    wire[31:0] ptw_io_requestor_1_pmp_7_mask;
    wire ptw_io_requestor_1_customCSRs_csrs_0_ren;
    wire ptw_io_requestor_1_customCSRs_csrs_0_wen;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_0_wdata;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_0_value;
    wire ptw_io_requestor_1_customCSRs_csrs_0_stall;
    wire ptw_io_requestor_1_customCSRs_csrs_0_set;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_0_sdata;
    wire ptw_io_requestor_1_customCSRs_csrs_1_ren;
    wire ptw_io_requestor_1_customCSRs_csrs_1_wen;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_1_wdata;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_1_value;
    wire ptw_io_requestor_1_customCSRs_csrs_1_stall;
    wire ptw_io_requestor_1_customCSRs_csrs_1_set;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_1_sdata;
    wire ptw_io_requestor_1_customCSRs_csrs_2_ren;
    wire ptw_io_requestor_1_customCSRs_csrs_2_wen;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_2_wdata;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_2_value;
    wire ptw_io_requestor_1_customCSRs_csrs_2_stall;
    wire ptw_io_requestor_1_customCSRs_csrs_2_set;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_2_sdata;
    wire ptw_io_requestor_1_customCSRs_csrs_3_ren;
    wire ptw_io_requestor_1_customCSRs_csrs_3_wen;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_3_wdata;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_3_value;
    wire ptw_io_requestor_1_customCSRs_csrs_3_stall;
    wire ptw_io_requestor_1_customCSRs_csrs_3_set;
    wire[63:0] ptw_io_requestor_1_customCSRs_csrs_3_sdata;
    wire ptw_io_mem_req_ready;
    wire ptw_io_mem_req_valid;
    wire[33:0] ptw_io_mem_req_bits_addr;
    wire[5:0] ptw_io_mem_req_bits_tag;
    wire[4:0] ptw_io_mem_req_bits_cmd;
    wire[1:0] ptw_io_mem_req_bits_size;
    wire ptw_io_mem_req_bits_signed;
    wire[1:0] ptw_io_mem_req_bits_dprv;
    wire ptw_io_mem_req_bits_dv;
    wire ptw_io_mem_req_bits_phys;
    wire ptw_io_mem_req_bits_no_alloc;
    wire ptw_io_mem_req_bits_no_xcpt;
    wire[63:0] ptw_io_mem_req_bits_data;
    wire[7:0] ptw_io_mem_req_bits_mask;
    wire ptw_io_mem_s1_kill;
    wire[63:0] ptw_io_mem_s1_data_data;
    wire[7:0] ptw_io_mem_s1_data_mask;
    wire ptw_io_mem_s2_nack;
    wire ptw_io_mem_s2_nack_cause_raw;
    wire ptw_io_mem_s2_kill;
    wire ptw_io_mem_s2_uncached;
    wire[31:0] ptw_io_mem_s2_paddr;
    wire ptw_io_mem_resp_valid;
    wire[33:0] ptw_io_mem_resp_bits_addr;
    wire[5:0] ptw_io_mem_resp_bits_tag;
    wire[4:0] ptw_io_mem_resp_bits_cmd;
    wire[1:0] ptw_io_mem_resp_bits_size;
    wire ptw_io_mem_resp_bits_signed;
    wire[1:0] ptw_io_mem_resp_bits_dprv;
    wire ptw_io_mem_resp_bits_dv;
    wire[63:0] ptw_io_mem_resp_bits_data;
    wire[7:0] ptw_io_mem_resp_bits_mask;
    wire ptw_io_mem_resp_bits_replay;
    wire ptw_io_mem_resp_bits_has_data;
    wire[63:0] ptw_io_mem_resp_bits_data_word_bypass;
    wire[63:0] ptw_io_mem_resp_bits_data_raw;
    wire[63:0] ptw_io_mem_resp_bits_store_data;
    wire ptw_io_mem_replay_next;
    wire ptw_io_mem_s2_xcpt_ma_ld;
    wire ptw_io_mem_s2_xcpt_ma_st;
    wire ptw_io_mem_s2_xcpt_pf_ld;
    wire ptw_io_mem_s2_xcpt_pf_st;
    wire ptw_io_mem_s2_xcpt_gf_ld;
    wire ptw_io_mem_s2_xcpt_gf_st;
    wire ptw_io_mem_s2_xcpt_ae_ld;
    wire ptw_io_mem_s2_xcpt_ae_st;
    wire[33:0] ptw_io_mem_s2_gpa;
    wire ptw_io_mem_s2_gpa_is_pte;
    wire ptw_io_mem_ordered;
    wire ptw_io_mem_perf_acquire;
    wire ptw_io_mem_perf_release;
    wire ptw_io_mem_perf_grant;
    wire ptw_io_mem_perf_tlbMiss;
    wire ptw_io_mem_perf_blocked;
    wire ptw_io_mem_perf_canAcceptStoreThenLoad;
    wire ptw_io_mem_perf_canAcceptStoreThenRMW;
    wire ptw_io_mem_perf_canAcceptLoadThenLoad;
    wire ptw_io_mem_perf_storeBufferEmptyAfterLoad;
    wire ptw_io_mem_perf_storeBufferEmptyAfterStore;
    wire ptw_io_mem_keep_clock_enabled;
    wire ptw_io_mem_clock_enabled;
    wire[3:0] ptw_io_dpath_ptbr_mode;
    wire[15:0] ptw_io_dpath_ptbr_asid;
    wire[43:0] ptw_io_dpath_ptbr_ppn;
    wire[3:0] ptw_io_dpath_hgatp_mode;
    wire[15:0] ptw_io_dpath_hgatp_asid;
    wire[43:0] ptw_io_dpath_hgatp_ppn;
    wire[3:0] ptw_io_dpath_vsatp_mode;
    wire[15:0] ptw_io_dpath_vsatp_asid;
    wire[43:0] ptw_io_dpath_vsatp_ppn;
    wire ptw_io_dpath_sfence_valid;
    wire ptw_io_dpath_sfence_bits_rs1;
    wire ptw_io_dpath_sfence_bits_rs2;
    wire[32:0] ptw_io_dpath_sfence_bits_addr;
    wire ptw_io_dpath_sfence_bits_asid;
    wire ptw_io_dpath_sfence_bits_hv;
    wire ptw_io_dpath_sfence_bits_hg;
    wire ptw_io_dpath_status_debug;
    wire ptw_io_dpath_status_cease;
    wire ptw_io_dpath_status_wfi;
    wire[31:0] ptw_io_dpath_status_isa;
    wire[1:0] ptw_io_dpath_status_dprv;
    wire ptw_io_dpath_status_dv;
    wire[1:0] ptw_io_dpath_status_prv;
    wire ptw_io_dpath_status_v;
    wire ptw_io_dpath_status_sd;
    wire[22:0] ptw_io_dpath_status_zero2;
    wire ptw_io_dpath_status_mpv;
    wire ptw_io_dpath_status_gva;
    wire ptw_io_dpath_status_mbe;
    wire ptw_io_dpath_status_sbe;
    wire[1:0] ptw_io_dpath_status_sxl;
    wire[1:0] ptw_io_dpath_status_uxl;
    wire ptw_io_dpath_status_sd_rv32;
    wire[7:0] ptw_io_dpath_status_zero1;
    wire ptw_io_dpath_status_tsr;
    wire ptw_io_dpath_status_tw;
    wire ptw_io_dpath_status_tvm;
    wire ptw_io_dpath_status_mxr;
    wire ptw_io_dpath_status_sum;
    wire ptw_io_dpath_status_mprv;
    wire[1:0] ptw_io_dpath_status_xs;
    wire[1:0] ptw_io_dpath_status_fs;
    wire[1:0] ptw_io_dpath_status_mpp;
    wire[1:0] ptw_io_dpath_status_vs;
    wire ptw_io_dpath_status_spp;
    wire ptw_io_dpath_status_mpie;
    wire ptw_io_dpath_status_ube;
    wire ptw_io_dpath_status_spie;
    wire ptw_io_dpath_status_upie;
    wire ptw_io_dpath_status_mie;
    wire ptw_io_dpath_status_hie;
    wire ptw_io_dpath_status_sie;
    wire ptw_io_dpath_status_uie;
    wire[29:0] ptw_io_dpath_hstatus_zero6;
    wire[1:0] ptw_io_dpath_hstatus_vsxl;
    wire[8:0] ptw_io_dpath_hstatus_zero5;
    wire ptw_io_dpath_hstatus_vtsr;
    wire ptw_io_dpath_hstatus_vtw;
    wire ptw_io_dpath_hstatus_vtvm;
    wire[1:0] ptw_io_dpath_hstatus_zero3;
    wire[5:0] ptw_io_dpath_hstatus_vgein;
    wire[1:0] ptw_io_dpath_hstatus_zero2;
    wire ptw_io_dpath_hstatus_hu;
    wire ptw_io_dpath_hstatus_spvp;
    wire ptw_io_dpath_hstatus_spv;
    wire ptw_io_dpath_hstatus_gva;
    wire ptw_io_dpath_hstatus_vsbe;
    wire[4:0] ptw_io_dpath_hstatus_zero1;
    wire ptw_io_dpath_gstatus_debug;
    wire ptw_io_dpath_gstatus_cease;
    wire ptw_io_dpath_gstatus_wfi;
    wire[31:0] ptw_io_dpath_gstatus_isa;
    wire[1:0] ptw_io_dpath_gstatus_dprv;
    wire ptw_io_dpath_gstatus_dv;
    wire[1:0] ptw_io_dpath_gstatus_prv;
    wire ptw_io_dpath_gstatus_v;
    wire ptw_io_dpath_gstatus_sd;
    wire[22:0] ptw_io_dpath_gstatus_zero2;
    wire ptw_io_dpath_gstatus_mpv;
    wire ptw_io_dpath_gstatus_gva;
    wire ptw_io_dpath_gstatus_mbe;
    wire ptw_io_dpath_gstatus_sbe;
    wire[1:0] ptw_io_dpath_gstatus_sxl;
    wire[1:0] ptw_io_dpath_gstatus_uxl;
    wire ptw_io_dpath_gstatus_sd_rv32;
    wire[7:0] ptw_io_dpath_gstatus_zero1;
    wire ptw_io_dpath_gstatus_tsr;
    wire ptw_io_dpath_gstatus_tw;
    wire ptw_io_dpath_gstatus_tvm;
    wire ptw_io_dpath_gstatus_mxr;
    wire ptw_io_dpath_gstatus_sum;
    wire ptw_io_dpath_gstatus_mprv;
    wire[1:0] ptw_io_dpath_gstatus_xs;
    wire[1:0] ptw_io_dpath_gstatus_fs;
    wire[1:0] ptw_io_dpath_gstatus_mpp;
    wire[1:0] ptw_io_dpath_gstatus_vs;
    wire ptw_io_dpath_gstatus_spp;
    wire ptw_io_dpath_gstatus_mpie;
    wire ptw_io_dpath_gstatus_ube;
    wire ptw_io_dpath_gstatus_spie;
    wire ptw_io_dpath_gstatus_upie;
    wire ptw_io_dpath_gstatus_mie;
    wire ptw_io_dpath_gstatus_hie;
    wire ptw_io_dpath_gstatus_sie;
    wire ptw_io_dpath_gstatus_uie;
    wire ptw_io_dpath_pmp_0_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_0_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_0_cfg_a;
    wire ptw_io_dpath_pmp_0_cfg_x;
    wire ptw_io_dpath_pmp_0_cfg_w;
    wire ptw_io_dpath_pmp_0_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_0_addr;
    wire[31:0] ptw_io_dpath_pmp_0_mask;
    wire ptw_io_dpath_pmp_1_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_1_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_1_cfg_a;
    wire ptw_io_dpath_pmp_1_cfg_x;
    wire ptw_io_dpath_pmp_1_cfg_w;
    wire ptw_io_dpath_pmp_1_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_1_addr;
    wire[31:0] ptw_io_dpath_pmp_1_mask;
    wire ptw_io_dpath_pmp_2_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_2_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_2_cfg_a;
    wire ptw_io_dpath_pmp_2_cfg_x;
    wire ptw_io_dpath_pmp_2_cfg_w;
    wire ptw_io_dpath_pmp_2_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_2_addr;
    wire[31:0] ptw_io_dpath_pmp_2_mask;
    wire ptw_io_dpath_pmp_3_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_3_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_3_cfg_a;
    wire ptw_io_dpath_pmp_3_cfg_x;
    wire ptw_io_dpath_pmp_3_cfg_w;
    wire ptw_io_dpath_pmp_3_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_3_addr;
    wire[31:0] ptw_io_dpath_pmp_3_mask;
    wire ptw_io_dpath_pmp_4_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_4_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_4_cfg_a;
    wire ptw_io_dpath_pmp_4_cfg_x;
    wire ptw_io_dpath_pmp_4_cfg_w;
    wire ptw_io_dpath_pmp_4_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_4_addr;
    wire[31:0] ptw_io_dpath_pmp_4_mask;
    wire ptw_io_dpath_pmp_5_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_5_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_5_cfg_a;
    wire ptw_io_dpath_pmp_5_cfg_x;
    wire ptw_io_dpath_pmp_5_cfg_w;
    wire ptw_io_dpath_pmp_5_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_5_addr;
    wire[31:0] ptw_io_dpath_pmp_5_mask;
    wire ptw_io_dpath_pmp_6_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_6_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_6_cfg_a;
    wire ptw_io_dpath_pmp_6_cfg_x;
    wire ptw_io_dpath_pmp_6_cfg_w;
    wire ptw_io_dpath_pmp_6_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_6_addr;
    wire[31:0] ptw_io_dpath_pmp_6_mask;
    wire ptw_io_dpath_pmp_7_cfg_l;
    wire[1:0] ptw_io_dpath_pmp_7_cfg_res;
    wire[1:0] ptw_io_dpath_pmp_7_cfg_a;
    wire ptw_io_dpath_pmp_7_cfg_x;
    wire ptw_io_dpath_pmp_7_cfg_w;
    wire ptw_io_dpath_pmp_7_cfg_r;
    wire[29:0] ptw_io_dpath_pmp_7_addr;
    wire[31:0] ptw_io_dpath_pmp_7_mask;
    wire ptw_io_dpath_perf_l2miss;
    wire ptw_io_dpath_perf_l2hit;
    wire ptw_io_dpath_perf_pte_miss;
    wire ptw_io_dpath_perf_pte_hit;
    wire ptw_io_dpath_customCSRs_csrs_0_ren;
    wire ptw_io_dpath_customCSRs_csrs_0_wen;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_0_wdata;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_0_value;
    wire ptw_io_dpath_customCSRs_csrs_0_stall;
    wire ptw_io_dpath_customCSRs_csrs_0_set;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_0_sdata;
    wire ptw_io_dpath_customCSRs_csrs_1_ren;
    wire ptw_io_dpath_customCSRs_csrs_1_wen;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_1_wdata;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_1_value;
    wire ptw_io_dpath_customCSRs_csrs_1_stall;
    wire ptw_io_dpath_customCSRs_csrs_1_set;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_1_sdata;
    wire ptw_io_dpath_customCSRs_csrs_2_ren;
    wire ptw_io_dpath_customCSRs_csrs_2_wen;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_2_wdata;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_2_value;
    wire ptw_io_dpath_customCSRs_csrs_2_stall;
    wire ptw_io_dpath_customCSRs_csrs_2_set;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_2_sdata;
    wire ptw_io_dpath_customCSRs_csrs_3_ren;
    wire ptw_io_dpath_customCSRs_csrs_3_wen;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_3_wdata;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_3_value;
    wire ptw_io_dpath_customCSRs_csrs_3_stall;
    wire ptw_io_dpath_customCSRs_csrs_3_set;
    wire[63:0] ptw_io_dpath_customCSRs_csrs_3_sdata;
    wire ptw_io_dpath_clock_enabled;

    wire ptw_pte_v ; 
    wire[9:0] ptw_tmp_reserved_for_future ; 
    wire[1:0] ptw_tmp_reserved_for_software ; 
    wire ptw_tmp_d ; 
    wire ptw_tmp_a ; 
    wire ptw_tmp_g ; 
    wire ptw_tmp_u ; 
    wire ptw_tmp_x ; 
    wire ptw_tmp_w ; 
    wire ptw_tmp_r ; 
    wire ptw__GEN ; 
    wire[9:0] ptw__r_pte_barrier_io_y_reserved_for_future ; 
    wire[43:0] ptw__r_pte_barrier_io_y_ppn ; 
    wire[1:0] ptw__r_pte_barrier_io_y_reserved_for_software ; 
    wire ptw__r_pte_barrier_io_y_d ; 
    wire ptw__r_pte_barrier_io_y_a ; 
    wire ptw__r_pte_barrier_io_y_g ; 
    wire ptw__r_pte_barrier_io_y_u ; 
    wire ptw__r_pte_barrier_io_y_x ; 
    wire ptw__r_pte_barrier_io_y_w ; 
    wire ptw__r_pte_barrier_io_y_r ; 
    wire ptw__r_pte_barrier_io_y_v ; 
    wire[2:0] ptw__state_barrier_io_y ; 
    wire ptw__arb_io_out_valid ; 
    wire ptw__arb_io_out_bits_valid ; 
    wire[20:0] ptw__arb_io_out_bits_bits_addr ; 
    wire ptw__arb_io_out_bits_bits_need_gpa ; 
    wire ptw__arb_io_out_bits_bits_vstage1 ; 
    wire ptw__arb_io_out_bits_bits_stage2 ; 
    wire ptw__arb_io_chosen ; 
    wire[29:0] ptw__pmpHomogeneous_WIRE_addr =30'h0; 
    wire[9:0] ptw__GEN_0 =10'h0; 
    wire[43:0] ptw__GEN_1 =44'h0; 
    wire[33:0] ptw_tag_1 =34'h200000000; 
    wire[31:0] ptw__pmpHomogeneous_WIRE_mask =32'h0; 
    wire[1:0] ptw_r_hgatp_initial_count =2'h0; 
    wire[1:0] ptw_count_1 =2'h0; 
    wire[1:0] ptw__GEN_2 =2'h0; 
    wire[1:0] ptw__pmpHomogeneous_WIRE_cfg_res =2'h0; 
    wire[1:0] ptw__pmpHomogeneous_WIRE_cfg_a =2'h0; 
    wire[1:0] ptw_satp_initial_count =2'h0; 
    wire[1:0] ptw_vsatp_initial_count =2'h0; 
    wire[1:0] ptw_hgatp_initial_count =2'h0; 
    wire[1:0] ptw_resp_gf_count =2'h0; 
    wire[1:0] ptw_r_pte_count =2'h0; 
    wire[1:0] ptw_r_pte_count_1 =2'h0; 
    wire[1:0] ptw_r_pte_count_2 =2'h0; 
    wire ptw__io_dpath_perf_l2hit_output =1'h0; 
    wire ptw__resp_valid_WIRE_0 =1'h0; 
    wire ptw__resp_valid_WIRE_1 =1'h0; 
    wire ptw__GEN_3 =1'h0; 
    wire ptw__GEN_4 =1'h0; 
    wire ptw__GEN_5 =1'h0; 
    wire ptw__GEN_6 =1'h0; 
    wire ptw__GEN_7 =1'h0; 
    wire ptw__GEN_8 =1'h0; 
    wire ptw__GEN_9 =1'h0; 
    wire ptw__GEN_10 =1'h0; 
    wire ptw__pmpHomogeneous_WIRE_cfg_l =1'h0; 
    wire ptw__pmpHomogeneous_WIRE_cfg_x =1'h0; 
    wire ptw__pmpHomogeneous_WIRE_cfg_w =1'h0; 
    wire ptw__pmpHomogeneous_WIRE_cfg_r =1'h0; 
    wire ptw_r_pte_idxs_0 =1'h0; reg[2:0] ptw_state ;  
    wire ptw_arb_clock;
    wire ptw_arb_reset;
    wire ptw_arb_io_in_0_ready;
    wire ptw_arb_io_in_0_valid;
    wire ptw_arb_io_in_0_bits_valid;
    wire[20:0] ptw_arb_io_in_0_bits_bits_addr;
    wire ptw_arb_io_in_0_bits_bits_need_gpa;
    wire ptw_arb_io_in_0_bits_bits_vstage1;
    wire ptw_arb_io_in_0_bits_bits_stage2;
    wire ptw_arb_io_in_1_ready;
    wire ptw_arb_io_in_1_valid;
    wire ptw_arb_io_in_1_bits_valid;
    wire[20:0] ptw_arb_io_in_1_bits_bits_addr;
    wire ptw_arb_io_in_1_bits_bits_need_gpa;
    wire ptw_arb_io_in_1_bits_bits_vstage1;
    wire ptw_arb_io_in_1_bits_bits_stage2;
    wire ptw_arb_io_out_ready;
    wire ptw_arb_io_out_valid;
    wire ptw_arb_io_out_bits_valid;
    wire[20:0] ptw_arb_io_out_bits_bits_addr;
    wire ptw_arb_io_out_bits_bits_need_gpa;
    wire ptw_arb_io_out_bits_bits_vstage1;
    wire ptw_arb_io_out_bits_bits_stage2;
    wire ptw_arb_io_chosen;

    wire ptw_arb_grant_1 = ptw_arb_io_in_0_valid ==1'h0; 
  assign  ptw_arb_io_in_0_ready = ptw_arb_io_out_ready &1'h1; 
  assign  ptw_arb_io_in_1_ready = ptw_arb_grant_1 & ptw_arb_io_out_ready ; 
  assign  ptw_arb_io_out_valid = ptw_arb_grant_1 ==1'h0| ptw_arb_io_in_1_valid ; 
  assign  ptw_arb_io_out_bits_valid = ptw_arb_io_in_0_valid  ?  ptw_arb_io_in_0_bits_valid : ptw_arb_io_in_1_bits_valid ; 
  assign  ptw_arb_io_out_bits_bits_addr = ptw_arb_io_in_0_valid  ?  ptw_arb_io_in_0_bits_bits_addr : ptw_arb_io_in_1_bits_bits_addr ; 
  assign  ptw_arb_io_out_bits_bits_need_gpa = ptw_arb_io_in_0_valid  ?  ptw_arb_io_in_0_bits_bits_need_gpa : ptw_arb_io_in_1_bits_bits_need_gpa ; 
  assign  ptw_arb_io_out_bits_bits_vstage1 = ptw_arb_io_in_0_valid  ?  ptw_arb_io_in_0_bits_bits_vstage1 : ptw_arb_io_in_1_bits_bits_vstage1 ; 
  assign  ptw_arb_io_out_bits_bits_stage2 = ptw_arb_io_in_0_valid  ?  ptw_arb_io_in_0_bits_bits_stage2 : ptw_arb_io_in_1_bits_bits_stage2 ; 
  assign  ptw_arb_io_chosen = ptw_arb_io_in_0_valid  ? 1'h0:1'h1;
    assign ptw_arb_clock = ptw_clock;
    assign ptw_arb_reset = ptw_reset;
    assign ptw_io_requestor_0_req_ready = ptw_arb_io_in_0_ready;
    assign ptw_arb_io_in_0_valid = ptw_io_requestor_0_req_valid;
    assign ptw_arb_io_in_0_bits_valid = ptw_io_requestor_0_req_bits_valid;
    assign ptw_arb_io_in_0_bits_bits_addr = ptw_io_requestor_0_req_bits_bits_addr;
    assign ptw_arb_io_in_0_bits_bits_need_gpa = ptw_io_requestor_0_req_bits_bits_need_gpa;
    assign ptw_arb_io_in_0_bits_bits_vstage1 = ptw_io_requestor_0_req_bits_bits_vstage1;
    assign ptw_arb_io_in_0_bits_bits_stage2 = ptw_io_requestor_0_req_bits_bits_stage2;
    assign ptw_io_requestor_1_req_ready = ptw_arb_io_in_1_ready;
    assign ptw_arb_io_in_1_valid = ptw_io_requestor_1_req_valid;
    assign ptw_arb_io_in_1_bits_valid = ptw_io_requestor_1_req_bits_valid;
    assign ptw_arb_io_in_1_bits_bits_addr = ptw_io_requestor_1_req_bits_bits_addr;
    assign ptw_arb_io_in_1_bits_bits_need_gpa = ptw_io_requestor_1_req_bits_bits_need_gpa;
    assign ptw_arb_io_in_1_bits_bits_vstage1 = ptw_io_requestor_1_req_bits_bits_vstage1;
    assign ptw_arb_io_in_1_bits_bits_stage2 = ptw_io_requestor_1_req_bits_bits_stage2;
    assign ptw_arb_io_out_ready = ptw__GEN;
    assign ptw__arb_io_out_valid = ptw_arb_io_out_valid;
    assign ptw__arb_io_out_bits_valid = ptw_arb_io_out_bits_valid;
    assign ptw__arb_io_out_bits_bits_addr = ptw_arb_io_out_bits_bits_addr;
    assign ptw__arb_io_out_bits_bits_need_gpa = ptw_arb_io_out_bits_bits_need_gpa;
    assign ptw__arb_io_out_bits_bits_vstage1 = ptw_arb_io_out_bits_bits_vstage1;
    assign ptw__arb_io_out_bits_bits_stage2 = ptw_arb_io_out_bits_bits_stage2;
    assign ptw__arb_io_chosen = ptw_arb_io_chosen;
     
    wire ptw_l2_refill_wire ; 
  assign  ptw__GEN = ptw_state ==3'h0& ptw_l2_refill_wire ==1'h0; 
    reg ptw_resp_valid_0 ; 
    reg ptw_resp_valid_1 ; 
    wire ptw_clock_en =(| ptw_state )| ptw_l2_refill_wire | ptw__arb_io_out_valid | ptw_io_dpath_sfence_valid | ptw_io_dpath_customCSRs_csrs_0_value [0]; 
    reg ptw_invalidated ; reg[1:0] ptw_count ; 
    reg ptw_resp_ae_ptw ; 
    reg ptw_resp_ae_final ; 
    reg ptw_resp_pf ; 
    reg ptw_resp_gf ; 
    reg ptw_resp_hr ; 
    reg ptw_resp_hw ; 
    reg ptw_resp_hx ; 
    reg ptw_resp_fragmented_superpage ; reg[20:0] ptw_r_req_addr ; 
    reg ptw_r_req_need_gpa ; 
    reg ptw_r_req_vstage1 ; 
    reg ptw_r_req_stage2 ; 
    reg ptw_r_req_dest ; reg[9:0] ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_2_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_3_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_4_reserved_for_future = ptw_r_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_5_reserved_for_future = ptw_r_pte_reserved_for_future ; reg[43:0] ptw_r_pte_ppn ; reg[1:0] ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_2_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_3_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_4_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_5_reserved_for_software = ptw_r_pte_reserved_for_software ; 
    reg ptw_r_pte_d ; 
    wire ptw_r_pte_pte_2_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_3_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_4_d = ptw_r_pte_d ; 
    wire ptw_r_pte_pte_5_d = ptw_r_pte_d ; 
    reg ptw_r_pte_a ; 
    wire ptw_r_pte_pte_2_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_3_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_4_a = ptw_r_pte_a ; 
    wire ptw_r_pte_pte_5_a = ptw_r_pte_a ; 
    reg ptw_r_pte_g ; 
    wire ptw_r_pte_pte_2_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_3_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_4_g = ptw_r_pte_g ; 
    wire ptw_r_pte_pte_5_g = ptw_r_pte_g ; 
    reg ptw_r_pte_u ; 
    wire ptw_r_pte_pte_2_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_3_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_4_u = ptw_r_pte_u ; 
    wire ptw_r_pte_pte_5_u = ptw_r_pte_u ; 
    reg ptw_r_pte_x ; 
    wire ptw_r_pte_pte_2_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_3_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_4_x = ptw_r_pte_x ; 
    wire ptw_r_pte_pte_5_x = ptw_r_pte_x ; 
    reg ptw_r_pte_w ; 
    wire ptw_r_pte_pte_2_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_3_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_4_w = ptw_r_pte_w ; 
    wire ptw_r_pte_pte_5_w = ptw_r_pte_w ; 
    reg ptw_r_pte_r ; 
    wire ptw_r_pte_pte_2_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_3_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_4_r = ptw_r_pte_r ; 
    wire ptw_r_pte_pte_5_r = ptw_r_pte_r ; 
    reg ptw_r_pte_v ; 
    wire ptw_r_pte_pte_2_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_3_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_4_v = ptw_r_pte_v ; 
    wire ptw_r_pte_pte_5_v = ptw_r_pte_v ; reg[3:0] ptw_r_hgatp_mode ; reg[15:0] ptw_r_hgatp_asid ; reg[43:0] ptw_r_hgatp_ppn ; reg[1:0] ptw_aux_count ; reg[9:0] ptw_aux_pte_reserved_for_future ; 
    wire[9:0] ptw_merged_pte_reserved_for_future = ptw_aux_pte_reserved_for_future ; reg[43:0] ptw_aux_pte_ppn ; reg[1:0] ptw_aux_pte_reserved_for_software ; 
    wire[1:0] ptw_merged_pte_reserved_for_software = ptw_aux_pte_reserved_for_software ; 
    reg ptw_aux_pte_d ; 
    wire ptw_merged_pte_d = ptw_aux_pte_d ; 
    reg ptw_aux_pte_a ; 
    wire ptw_merged_pte_a = ptw_aux_pte_a ; 
    reg ptw_aux_pte_g ; 
    wire ptw_merged_pte_g = ptw_aux_pte_g ; 
    reg ptw_aux_pte_u ; 
    wire ptw_merged_pte_u = ptw_aux_pte_u ; 
    reg ptw_aux_pte_x ; 
    wire ptw_merged_pte_x = ptw_aux_pte_x ; 
    reg ptw_aux_pte_w ; 
    wire ptw_merged_pte_w = ptw_aux_pte_w ; 
    reg ptw_aux_pte_r ; 
    wire ptw_merged_pte_r = ptw_aux_pte_r ; 
    reg ptw_aux_pte_v ; 
    wire ptw_merged_pte_v = ptw_aux_pte_v ; reg[11:0] ptw_gpa_pgoff ; 
    reg ptw_stage2 ; 
    reg ptw_stage2_final ; 
    wire[3:0] ptw_satp_mode = ptw__arb_io_out_bits_bits_vstage1  ?  ptw_io_dpath_vsatp_mode : ptw_io_dpath_ptbr_mode ; 
    wire[15:0] ptw_satp_asid = ptw__arb_io_out_bits_bits_vstage1  ?  ptw_io_dpath_vsatp_asid : ptw_io_dpath_ptbr_asid ; 
    wire[43:0] ptw_satp_ppn = ptw__arb_io_out_bits_bits_vstage1  ?  ptw_io_dpath_vsatp_ppn : ptw_io_dpath_ptbr_ppn ; 
    wire[43:0] ptw_r_pte_pte_5_ppn = ptw_satp_ppn ; 
    wire ptw_do_both_stages = ptw_r_req_vstage1 & ptw_r_req_stage2 ; 
    wire[1:0] ptw_max_count = ptw_count < ptw_aux_count  ?  ptw_aux_count : ptw_count ; 
    wire[43:0] ptw_vpn = ptw_r_req_vstage1 & ptw_stage2  ?  ptw_aux_pte_ppn :{23'h0, ptw_r_req_addr }; 
    reg ptw_mem_resp_valid ; reg[63:0] ptw_mem_resp_data ; 
    wire[63:0] ptw__tmp_WIRE = ptw_mem_resp_data ; 
    wire[9:0] ptw_pte_reserved_for_future = ptw_tmp_reserved_for_future ; 
    wire[1:0] ptw_pte_reserved_for_software = ptw_tmp_reserved_for_software ; 
    wire ptw_pte_d = ptw_tmp_d ; 
    wire ptw_pte_a = ptw_tmp_a ; 
    wire ptw_pte_g = ptw_tmp_g ; 
    wire ptw_pte_u = ptw_tmp_u ; 
    wire ptw_pte_x = ptw_tmp_x ; 
    wire ptw_pte_w = ptw_tmp_w ; 
    wire ptw_pte_r = ptw_tmp_r ; 
    wire ptw_tmp_v = ptw__tmp_WIRE [0]; 
  assign  ptw_tmp_r = ptw__tmp_WIRE [1]; 
  assign  ptw_tmp_w = ptw__tmp_WIRE [2]; 
  assign  ptw_tmp_x = ptw__tmp_WIRE [3]; 
  assign  ptw_tmp_u = ptw__tmp_WIRE [4]; 
  assign  ptw_tmp_g = ptw__tmp_WIRE [5]; 
  assign  ptw_tmp_a = ptw__tmp_WIRE [6]; 
  assign  ptw_tmp_d = ptw__tmp_WIRE [7]; 
  assign  ptw_tmp_reserved_for_software = ptw__tmp_WIRE [9:8]; 
    wire[43:0] ptw_tmp_ppn = ptw__tmp_WIRE [53:10]; 
  assign  ptw_tmp_reserved_for_future = ptw__tmp_WIRE [63:54]; 
    wire[9:0] ptw_aux_pte_pte_reserved_for_future = ptw_pte_reserved_for_future ; 
    wire[1:0] ptw_aux_pte_pte_reserved_for_software = ptw_pte_reserved_for_software ; 
    wire ptw_aux_pte_pte_d = ptw_pte_d ; 
    wire ptw_aux_pte_pte_a = ptw_pte_a ; 
    wire ptw_aux_pte_pte_g = ptw_pte_g ; 
    wire ptw_aux_pte_pte_u = ptw_pte_u ; 
    wire ptw_aux_pte_pte_x = ptw_pte_x ; 
    wire ptw_aux_pte_pte_w = ptw_pte_w ; 
    wire ptw_aux_pte_pte_r = ptw_pte_r ; 
    wire ptw_aux_pte_pte_v = ptw_pte_v ; 
    wire[43:0] ptw_pte_ppn ={23'h0, ptw_do_both_stages & ptw_stage2 ==1'h0 ?  ptw_tmp_ppn [20:0]:{1'h0, ptw_tmp_ppn [19:0]}}; 
    wire ptw__GEN_11 = ptw_tmp_r | ptw_tmp_w | ptw_tmp_x ; 
    wire ptw__GEN_12 = ptw_count <=2'h0&(|( ptw_tmp_ppn [17:9])); 
    wire ptw__GEN_13 = ptw_count <=2'h1&(|( ptw_tmp_ppn [8:0])); 
  assign  ptw_pte_v = ptw__GEN_11  ? ( ptw__GEN_13  ? 1'h0: ptw__GEN_12  ? 1'h0: ptw_tmp_v ): ptw_tmp_v ; 
    wire ptw_invalid_paddr = ptw_do_both_stages & ptw_stage2 ==1'h0 ? (|( ptw_tmp_ppn [43:21])):(|( ptw_tmp_ppn [43:20])); 
    wire[14:0] ptw_idxs_0 = ptw_tmp_ppn [43:29]; 
    wire[14:0] ptw__GEN_14 = ptw_idxs_0 ; 
    wire ptw_invalid_gpa = ptw_do_both_stages & ptw_stage2 ==1'h0&(| ptw__GEN_14 ); 
    wire ptw_traverse = ptw_pte_v & ptw_pte_r ==1'h0& ptw_pte_w ==1'h0& ptw_pte_x ==1'h0& ptw_pte_d ==1'h0& ptw_pte_a ==1'h0& ptw_pte_u ==1'h0& ptw_pte_reserved_for_future ==10'h0& ptw_invalid_paddr ==1'h0& ptw_invalid_gpa ==1'h0& ptw_count <2'h2; reg[6:0] ptw_state_reg ; reg[7:0] ptw_valid ; reg[31:0] ptw_tags_0 ; reg[31:0] ptw_tags_1 ; reg[31:0] ptw_tags_2 ; reg[31:0] ptw_tags_3 ; reg[31:0] ptw_tags_4 ; reg[31:0] ptw_tags_5 ; reg[31:0] ptw_tags_6 ; reg[31:0] ptw_tags_7 ; reg[19:0] ptw_data_0 ; reg[19:0] ptw_data_1 ; reg[19:0] ptw_data_2 ; reg[19:0] ptw_data_3 ; reg[19:0] ptw_data_4 ; reg[19:0] ptw_data_5 ; reg[19:0] ptw_data_6 ; reg[19:0] ptw_data_7 ; 
    wire ptw_can_hit = ptw_count <2'h2&( ptw_r_req_vstage1  ?  ptw_stage2 : ptw_r_req_stage2 ==1'h0); 
    wire[32:0] ptw_tag ={ ptw_r_req_vstage1 ,32'h0}; 
    wire[1:0] ptw_hits_lo_lo ={{1'h0, ptw_tags_1 }== ptw_tag ,{1'h0, ptw_tags_0 }== ptw_tag }; 
    wire[1:0] ptw_hits_lo_hi ={{1'h0, ptw_tags_3 }== ptw_tag ,{1'h0, ptw_tags_2 }== ptw_tag }; 
    wire[3:0] ptw_hits_lo ={ ptw_hits_lo_hi , ptw_hits_lo_lo }; 
    wire[1:0] ptw_hits_hi_lo ={{1'h0, ptw_tags_5 }== ptw_tag ,{1'h0, ptw_tags_4 }== ptw_tag }; 
    wire[1:0] ptw_hits_hi_hi ={{1'h0, ptw_tags_7 }== ptw_tag ,{1'h0, ptw_tags_6 }== ptw_tag }; 
    wire[3:0] ptw_hits_hi ={ ptw_hits_hi_hi , ptw_hits_hi_lo }; 
    wire[7:0] ptw_hits ={ ptw_hits_hi , ptw_hits_lo }& ptw_valid ; 
    wire ptw_pte_cache_hit =(| ptw_hits )& ptw_can_hit ; 
    wire ptw__GEN_15 = ptw_mem_resp_valid & ptw_traverse & ptw_can_hit &(| ptw_hits )==1'h0& ptw_invalidated ==1'h0; 
    wire ptw_r_left_subtree_older = ptw_state_reg [6]; 
    wire[2:0] ptw_r_left_subtree_state = ptw_state_reg [5:3]; 
    wire[2:0] ptw_r_right_subtree_state = ptw_state_reg [2:0]; 
    wire ptw_r_left_subtree_older_1 = ptw_r_left_subtree_state [2]; 
    wire ptw_r_left_subtree_state_1 = ptw_r_left_subtree_state [1]; 
    wire ptw_r_right_subtree_state_1 = ptw_r_left_subtree_state [0]; 
    wire ptw_r_left_subtree_older_2 = ptw_r_right_subtree_state [2]; 
    wire ptw_r_left_subtree_state_2 = ptw_r_right_subtree_state [1]; 
    wire ptw_r_right_subtree_state_2 = ptw_r_right_subtree_state [0]; 
    wire[7:0] ptw__GEN_16 =~ ptw_valid ; 
    wire[2:0] ptw_r =(& ptw_valid ) ? { ptw_r_left_subtree_older , ptw_r_left_subtree_older  ? { ptw_r_left_subtree_older_1 , ptw_r_left_subtree_older_1  ?  ptw_r_left_subtree_state_1 : ptw_r_right_subtree_state_1 }:{ ptw_r_left_subtree_older_2 , ptw_r_left_subtree_older_2  ?  ptw_r_left_subtree_state_2 : ptw_r_right_subtree_state_2 }}: ptw__GEN_16 [0] ? 3'h0: ptw__GEN_16 [1] ? 3'h1: ptw__GEN_16 [2] ? 3'h2: ptw__GEN_16 [3] ? 3'h3: ptw__GEN_16 [4] ? 3'h4: ptw__GEN_16 [5] ? 3'h5: ptw__GEN_16 [6] ? 3'h6:3'h7; 
    wire[2:0] ptw_state_reg_touch_way_sized = ptw_r ; 
    wire[7:0] ptw__GEN_17 = ptw_valid |8'h1<< ptw_r ; 
    wire ptw__GEN_18 = ptw_r ==3'h0; 
    wire ptw__GEN_19 = ptw_r ==3'h1; 
    wire ptw__GEN_20 = ptw_r ==3'h2; 
    wire ptw__GEN_21 = ptw_r ==3'h3; 
    wire ptw__GEN_22 = ptw_r ==3'h4; 
    wire ptw__GEN_23 = ptw_r ==3'h5; 
    wire ptw__GEN_24 = ptw_r ==3'h6; 
    wire ptw__GEN_25 =& ptw_r ; 
    wire ptw__GEN_26 = ptw_r ==3'h0; 
    wire ptw__GEN_27 = ptw_r ==3'h1; 
    wire ptw__GEN_28 = ptw_r ==3'h2; 
    wire ptw__GEN_29 = ptw_r ==3'h3; 
    wire ptw__GEN_30 = ptw_r ==3'h4; 
    wire ptw__GEN_31 = ptw_r ==3'h5; 
    wire ptw__GEN_32 = ptw_r ==3'h6; 
    wire ptw__GEN_33 =& ptw_r ; 
    wire ptw_state_reg_set_left_older = ptw_state_reg_touch_way_sized [2]==1'h0; 
    wire[2:0] ptw_state_reg_left_subtree_state = ptw_state_reg [5:3]; 
    wire[2:0] ptw_state_reg_right_subtree_state = ptw_state_reg [2:0]; 
    wire[1:0] ptw__state_reg_touch_way_sized_1to0 = ptw_state_reg_touch_way_sized [1:0]; 
    wire ptw_state_reg_set_left_older_1 = ptw__state_reg_touch_way_sized_1to0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_1 = ptw_state_reg_left_subtree_state [1]; 
    wire ptw_state_reg_right_subtree_state_1 = ptw_state_reg_left_subtree_state [0]; 
    wire[1:0] ptw_state_reg_hi ={ ptw_state_reg_set_left_older_1 , ptw_state_reg_set_left_older_1  ?  ptw_state_reg_left_subtree_state_1 : ptw__state_reg_touch_way_sized_1to0 [0]==1'h0}; 
    wire[1:0] ptw__state_reg_touch_way_sized_1to0_0 = ptw_state_reg_touch_way_sized [1:0]; 
    wire ptw_state_reg_set_left_older_2 = ptw__state_reg_touch_way_sized_1to0_0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_2 = ptw_state_reg_right_subtree_state [1]; 
    wire ptw_state_reg_right_subtree_state_2 = ptw_state_reg_right_subtree_state [0]; 
    wire[1:0] ptw_state_reg_hi_1 ={ ptw_state_reg_set_left_older_2 , ptw_state_reg_set_left_older_2  ?  ptw_state_reg_left_subtree_state_2 : ptw__state_reg_touch_way_sized_1to0_0 [0]==1'h0}; 
    wire[3:0] ptw_state_reg_hi_2 ={ ptw_state_reg_set_left_older , ptw_state_reg_set_left_older  ?  ptw_state_reg_left_subtree_state :{ ptw_state_reg_hi , ptw_state_reg_set_left_older_1  ?  ptw__state_reg_touch_way_sized_1to0 [0]==1'h0: ptw_state_reg_right_subtree_state_1 }}; 
    wire[6:0] ptw__GEN_34 ={ ptw_state_reg_hi_2 , ptw_state_reg_set_left_older  ? { ptw_state_reg_hi_1 , ptw_state_reg_set_left_older_2  ?  ptw__state_reg_touch_way_sized_1to0_0 [0]==1'h0: ptw_state_reg_right_subtree_state_2 }: ptw_state_reg_right_subtree_state }; 
    wire ptw__GEN_35 = ptw_pte_cache_hit & ptw_state ==3'h1; 
    wire[3:0] ptw_hi = ptw_hits [7:4]; 
    wire[3:0] ptw_lo = ptw_hits [3:0]; 
    wire[3:0] ptw__GEN_36 = ptw_hi | ptw_lo ; 
    wire[1:0] ptw_hi_1 = ptw__GEN_36 [3:2]; 
    wire[1:0] ptw_lo_1 = ptw__GEN_36 [1:0]; 
    wire[1:0] ptw__GEN_37 = ptw_hi_1 | ptw_lo_1 ; 
    wire[2:0] ptw_state_reg_touch_way_sized_1 ={| ptw_hi ,{| ptw_hi_1 , ptw__GEN_37 [1]}}; 
    wire ptw_state_reg_set_left_older_3 = ptw_state_reg_touch_way_sized_1 [2]==1'h0; 
    wire[2:0] ptw_state_reg_left_subtree_state_3 = ptw_state_reg [5:3]; 
    wire[2:0] ptw_state_reg_right_subtree_state_3 = ptw_state_reg [2:0]; 
    wire[1:0] ptw__state_reg_touch_way_sized_1_1to0 = ptw_state_reg_touch_way_sized_1 [1:0]; 
    wire ptw_state_reg_set_left_older_4 = ptw__state_reg_touch_way_sized_1_1to0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_4 = ptw_state_reg_left_subtree_state_3 [1]; 
    wire ptw_state_reg_right_subtree_state_4 = ptw_state_reg_left_subtree_state_3 [0]; 
    wire[1:0] ptw_state_reg_hi_3 ={ ptw_state_reg_set_left_older_4 , ptw_state_reg_set_left_older_4  ?  ptw_state_reg_left_subtree_state_4 : ptw__state_reg_touch_way_sized_1_1to0 [0]==1'h0}; 
    wire[1:0] ptw__state_reg_touch_way_sized_1_1to0_0 = ptw_state_reg_touch_way_sized_1 [1:0]; 
    wire ptw_state_reg_set_left_older_5 = ptw__state_reg_touch_way_sized_1_1to0_0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_5 = ptw_state_reg_right_subtree_state_3 [1]; 
    wire ptw_state_reg_right_subtree_state_5 = ptw_state_reg_right_subtree_state_3 [0]; 
    wire[1:0] ptw_state_reg_hi_4 ={ ptw_state_reg_set_left_older_5 , ptw_state_reg_set_left_older_5  ?  ptw_state_reg_left_subtree_state_5 : ptw__state_reg_touch_way_sized_1_1to0_0 [0]==1'h0}; 
    wire[3:0] ptw_state_reg_hi_5 ={ ptw_state_reg_set_left_older_3 , ptw_state_reg_set_left_older_3  ?  ptw_state_reg_left_subtree_state_3 :{ ptw_state_reg_hi_3 , ptw_state_reg_set_left_older_4  ?  ptw__state_reg_touch_way_sized_1_1to0 [0]==1'h0: ptw_state_reg_right_subtree_state_4 }}; 
    wire[6:0] ptw__GEN_38 ={ ptw_state_reg_hi_5 , ptw_state_reg_set_left_older_3  ? { ptw_state_reg_hi_4 , ptw_state_reg_set_left_older_5  ?  ptw__state_reg_touch_way_sized_1_1to0_0 [0]==1'h0: ptw_state_reg_right_subtree_state_5 }: ptw_state_reg_right_subtree_state_3 }; 
    wire ptw__GEN_39 = ptw_io_dpath_sfence_valid & ptw_io_dpath_sfence_bits_rs1 ==1'h0; 
    wire[19:0] ptw_pte_cache_data =( ptw_hits [0] ?  ptw_data_0 :20'h0)|( ptw_hits [1] ?  ptw_data_1 :20'h0)|( ptw_hits [2] ?  ptw_data_2 :20'h0)|( ptw_hits [3] ?  ptw_data_3 :20'h0)|( ptw_hits [4] ?  ptw_data_4 :20'h0)|( ptw_hits [5] ?  ptw_data_5 :20'h0)|( ptw_hits [6] ?  ptw_data_6 :20'h0)|( ptw_hits [7] ?  ptw_data_7 :20'h0); reg[6:0] ptw_state_reg_1 ; reg[7:0] ptw_valid_1 ; reg[31:0] ptw_tags_1_0 ; reg[31:0] ptw_tags_1_1 ; reg[31:0] ptw_tags_1_2 ; reg[31:0] ptw_tags_1_3 ; reg[31:0] ptw_tags_1_4 ; reg[31:0] ptw_tags_1_5 ; reg[31:0] ptw_tags_1_6 ; reg[31:0] ptw_tags_1_7 ; reg[19:0] ptw_data_1_0 ; reg[19:0] ptw_data_1_1 ; reg[19:0] ptw_data_1_2 ; reg[19:0] ptw_data_1_3 ; reg[19:0] ptw_data_1_4 ; reg[19:0] ptw_data_1_5 ; reg[19:0] ptw_data_1_6 ; reg[19:0] ptw_data_1_7 ; 
    wire ptw_can_hit_1 = ptw_count == ptw_r_hgatp_initial_count & ptw_aux_count <2'h2& ptw_r_req_vstage1 & ptw_stage2 & ptw_stage2_final ==1'h0; 
    wire ptw_can_refill = ptw_do_both_stages & ptw_stage2 ==1'h0& ptw_stage2_final ==1'h0; 
    wire[1:0] ptw_hits_lo_lo_1 ={{2'h0, ptw_tags_1_1 }== ptw_tag_1 ,{2'h0, ptw_tags_1_0 }== ptw_tag_1 }; 
    wire[1:0] ptw_hits_lo_hi_1 ={{2'h0, ptw_tags_1_3 }== ptw_tag_1 ,{2'h0, ptw_tags_1_2 }== ptw_tag_1 }; 
    wire[3:0] ptw_hits_lo_1 ={ ptw_hits_lo_hi_1 , ptw_hits_lo_lo_1 }; 
    wire[1:0] ptw_hits_hi_lo_1 ={{2'h0, ptw_tags_1_5 }== ptw_tag_1 ,{2'h0, ptw_tags_1_4 }== ptw_tag_1 }; 
    wire[1:0] ptw_hits_hi_hi_1 ={{2'h0, ptw_tags_1_7 }== ptw_tag_1 ,{2'h0, ptw_tags_1_6 }== ptw_tag_1 }; 
    wire[3:0] ptw_hits_hi_1 ={ ptw_hits_hi_hi_1 , ptw_hits_hi_lo_1 }; 
    wire[7:0] ptw_hits_1 ={ ptw_hits_hi_1 , ptw_hits_lo_1 }& ptw_valid_1 ; 
    wire ptw_stage2_pte_cache_hit =(| ptw_hits_1 )& ptw_can_hit_1 ; 
    wire ptw__GEN_40 = ptw_mem_resp_valid & ptw_traverse & ptw_can_refill &(| ptw_hits_1 )==1'h0& ptw_invalidated ==1'h0; 
    wire ptw_r_left_subtree_older_3 = ptw_state_reg_1 [6]; 
    wire[2:0] ptw_r_left_subtree_state_3 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_r_right_subtree_state_3 = ptw_state_reg_1 [2:0]; 
    wire ptw_r_left_subtree_older_4 = ptw_r_left_subtree_state_3 [2]; 
    wire ptw_r_left_subtree_state_4 = ptw_r_left_subtree_state_3 [1]; 
    wire ptw_r_right_subtree_state_4 = ptw_r_left_subtree_state_3 [0]; 
    wire ptw_r_left_subtree_older_5 = ptw_r_right_subtree_state_3 [2]; 
    wire ptw_r_left_subtree_state_5 = ptw_r_right_subtree_state_3 [1]; 
    wire ptw_r_right_subtree_state_5 = ptw_r_right_subtree_state_3 [0]; 
    wire[7:0] ptw__GEN_41 =~ ptw_valid_1 ; 
    wire[2:0] ptw_r_1 =(& ptw_valid_1 ) ? { ptw_r_left_subtree_older_3 , ptw_r_left_subtree_older_3  ? { ptw_r_left_subtree_older_4 , ptw_r_left_subtree_older_4  ?  ptw_r_left_subtree_state_4 : ptw_r_right_subtree_state_4 }:{ ptw_r_left_subtree_older_5 , ptw_r_left_subtree_older_5  ?  ptw_r_left_subtree_state_5 : ptw_r_right_subtree_state_5 }}: ptw__GEN_41 [0] ? 3'h0: ptw__GEN_41 [1] ? 3'h1: ptw__GEN_41 [2] ? 3'h2: ptw__GEN_41 [3] ? 3'h3: ptw__GEN_41 [4] ? 3'h4: ptw__GEN_41 [5] ? 3'h5: ptw__GEN_41 [6] ? 3'h6:3'h7; 
    wire[2:0] ptw_state_reg_touch_way_sized_2 = ptw_r_1 ; 
    wire[7:0] ptw__GEN_42 = ptw_valid_1 |8'h1<< ptw_r_1 ; 
    wire ptw__GEN_43 = ptw_r_1 ==3'h0; 
    wire ptw__GEN_44 = ptw_r_1 ==3'h1; 
    wire ptw__GEN_45 = ptw_r_1 ==3'h2; 
    wire ptw__GEN_46 = ptw_r_1 ==3'h3; 
    wire ptw__GEN_47 = ptw_r_1 ==3'h4; 
    wire ptw__GEN_48 = ptw_r_1 ==3'h5; 
    wire ptw__GEN_49 = ptw_r_1 ==3'h6; 
    wire ptw__GEN_50 =& ptw_r_1 ; 
    wire ptw__GEN_51 = ptw_r_1 ==3'h0; 
    wire ptw__GEN_52 = ptw_r_1 ==3'h1; 
    wire ptw__GEN_53 = ptw_r_1 ==3'h2; 
    wire ptw__GEN_54 = ptw_r_1 ==3'h3; 
    wire ptw__GEN_55 = ptw_r_1 ==3'h4; 
    wire ptw__GEN_56 = ptw_r_1 ==3'h5; 
    wire ptw__GEN_57 = ptw_r_1 ==3'h6; 
    wire ptw__GEN_58 =& ptw_r_1 ; 
    wire ptw_state_reg_set_left_older_6 = ptw_state_reg_touch_way_sized_2 [2]==1'h0; 
    wire[2:0] ptw_state_reg_left_subtree_state_6 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_state_reg_right_subtree_state_6 = ptw_state_reg_1 [2:0]; 
    wire[1:0] ptw__state_reg_touch_way_sized_2_1to0 = ptw_state_reg_touch_way_sized_2 [1:0]; 
    wire ptw_state_reg_set_left_older_7 = ptw__state_reg_touch_way_sized_2_1to0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_7 = ptw_state_reg_left_subtree_state_6 [1]; 
    wire ptw_state_reg_right_subtree_state_7 = ptw_state_reg_left_subtree_state_6 [0]; 
    wire[1:0] ptw_state_reg_hi_6 ={ ptw_state_reg_set_left_older_7 , ptw_state_reg_set_left_older_7  ?  ptw_state_reg_left_subtree_state_7 : ptw__state_reg_touch_way_sized_2_1to0 [0]==1'h0}; 
    wire[1:0] ptw__state_reg_touch_way_sized_2_1to0_0 = ptw_state_reg_touch_way_sized_2 [1:0]; 
    wire ptw_state_reg_set_left_older_8 = ptw__state_reg_touch_way_sized_2_1to0_0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_8 = ptw_state_reg_right_subtree_state_6 [1]; 
    wire ptw_state_reg_right_subtree_state_8 = ptw_state_reg_right_subtree_state_6 [0]; 
    wire[1:0] ptw_state_reg_hi_7 ={ ptw_state_reg_set_left_older_8 , ptw_state_reg_set_left_older_8  ?  ptw_state_reg_left_subtree_state_8 : ptw__state_reg_touch_way_sized_2_1to0_0 [0]==1'h0}; 
    wire[3:0] ptw_state_reg_hi_8 ={ ptw_state_reg_set_left_older_6 , ptw_state_reg_set_left_older_6  ?  ptw_state_reg_left_subtree_state_6 :{ ptw_state_reg_hi_6 , ptw_state_reg_set_left_older_7  ?  ptw__state_reg_touch_way_sized_2_1to0 [0]==1'h0: ptw_state_reg_right_subtree_state_7 }}; 
    wire[6:0] ptw__GEN_59 ={ ptw_state_reg_hi_8 , ptw_state_reg_set_left_older_6  ? { ptw_state_reg_hi_7 , ptw_state_reg_set_left_older_8  ?  ptw__state_reg_touch_way_sized_2_1to0_0 [0]==1'h0: ptw_state_reg_right_subtree_state_8 }: ptw_state_reg_right_subtree_state_6 }; 
    wire ptw__GEN_60 = ptw_stage2_pte_cache_hit & ptw_state ==3'h1; 
    wire[3:0] ptw_hi_2 = ptw_hits_1 [7:4]; 
    wire[3:0] ptw_lo_2 = ptw_hits_1 [3:0]; 
    wire[3:0] ptw__GEN_61 = ptw_hi_2 | ptw_lo_2 ; 
    wire[1:0] ptw_hi_3 = ptw__GEN_61 [3:2]; 
    wire[1:0] ptw_lo_3 = ptw__GEN_61 [1:0]; 
    wire[1:0] ptw__GEN_62 = ptw_hi_3 | ptw_lo_3 ; 
    wire[2:0] ptw_state_reg_touch_way_sized_3 ={| ptw_hi_2 ,{| ptw_hi_3 , ptw__GEN_62 [1]}}; 
    wire ptw_state_reg_set_left_older_9 = ptw_state_reg_touch_way_sized_3 [2]==1'h0; 
    wire[2:0] ptw_state_reg_left_subtree_state_9 = ptw_state_reg_1 [5:3]; 
    wire[2:0] ptw_state_reg_right_subtree_state_9 = ptw_state_reg_1 [2:0]; 
    wire[1:0] ptw__state_reg_touch_way_sized_3_1to0 = ptw_state_reg_touch_way_sized_3 [1:0]; 
    wire ptw_state_reg_set_left_older_10 = ptw__state_reg_touch_way_sized_3_1to0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_10 = ptw_state_reg_left_subtree_state_9 [1]; 
    wire ptw_state_reg_right_subtree_state_10 = ptw_state_reg_left_subtree_state_9 [0]; 
    wire[1:0] ptw_state_reg_hi_9 ={ ptw_state_reg_set_left_older_10 , ptw_state_reg_set_left_older_10  ?  ptw_state_reg_left_subtree_state_10 : ptw__state_reg_touch_way_sized_3_1to0 [0]==1'h0}; 
    wire[1:0] ptw__state_reg_touch_way_sized_3_1to0_0 = ptw_state_reg_touch_way_sized_3 [1:0]; 
    wire ptw_state_reg_set_left_older_11 = ptw__state_reg_touch_way_sized_3_1to0_0 [1]==1'h0; 
    wire ptw_state_reg_left_subtree_state_11 = ptw_state_reg_right_subtree_state_9 [1]; 
    wire ptw_state_reg_right_subtree_state_11 = ptw_state_reg_right_subtree_state_9 [0]; 
    wire[1:0] ptw_state_reg_hi_10 ={ ptw_state_reg_set_left_older_11 , ptw_state_reg_set_left_older_11  ?  ptw_state_reg_left_subtree_state_11 : ptw__state_reg_touch_way_sized_3_1to0_0 [0]==1'h0}; 
    wire[3:0] ptw_state_reg_hi_11 ={ ptw_state_reg_set_left_older_9 , ptw_state_reg_set_left_older_9  ?  ptw_state_reg_left_subtree_state_9 :{ ptw_state_reg_hi_9 , ptw_state_reg_set_left_older_10  ?  ptw__state_reg_touch_way_sized_3_1to0 [0]==1'h0: ptw_state_reg_right_subtree_state_10 }}; 
    wire[6:0] ptw__GEN_63 ={ ptw_state_reg_hi_11 , ptw_state_reg_set_left_older_9  ? { ptw_state_reg_hi_10 , ptw_state_reg_set_left_older_11  ?  ptw__state_reg_touch_way_sized_3_1to0_0 [0]==1'h0: ptw_state_reg_right_subtree_state_11 }: ptw_state_reg_right_subtree_state_9 }; 
    wire ptw__GEN_64 = ptw_io_dpath_sfence_valid & ptw_io_dpath_sfence_bits_rs1 ==1'h0; 
    wire[19:0] ptw_stage2_pte_cache_data =( ptw_hits_1 [0] ?  ptw_data_1_0 :20'h0)|( ptw_hits_1 [1] ?  ptw_data_1_1 :20'h0)|( ptw_hits_1 [2] ?  ptw_data_1_2 :20'h0)|( ptw_hits_1 [3] ?  ptw_data_1_3 :20'h0)|( ptw_hits_1 [4] ?  ptw_data_1_4 :20'h0)|( ptw_hits_1 [5] ?  ptw_data_1_5 :20'h0)|( ptw_hits_1 [6] ?  ptw_data_1_6 :20'h0)|( ptw_hits_1 [7] ?  ptw_data_1_7 :20'h0); 
    reg ptw_pte_hit ; 
    wire ptw__io_dpath_perf_pte_miss_output ; 
    wire ptw__io_dpath_perf_pte_hit_output = ptw_pte_hit & ptw_state ==3'h1& ptw__io_dpath_perf_l2hit_output ==1'h0; 
    wire ptw__GEN_65 =( ptw__io_dpath_perf_l2hit_output &( ptw__io_dpath_perf_pte_miss_output | ptw__io_dpath_perf_pte_hit_output ))==1'h0==1'h0; 
    reg ptw_l2_refill ; 
  assign  ptw_l2_refill_wire = ptw_l2_refill ; 
    wire[9:0] ptw_l2_pte_reserved_for_future = ptw__GEN_0 ; 
    wire[43:0] ptw_l2_pte_ppn = ptw__GEN_1 ; 
    wire[1:0] ptw_l2_pte_reserved_for_software = ptw__GEN_2 ; 
    wire ptw_l2_pte_d = ptw__GEN_3 ; 
    wire ptw_l2_pte_a = ptw__GEN_4 ; 
    wire ptw_l2_pte_g = ptw__GEN_5 ; 
    wire ptw_l2_pte_u = ptw__GEN_6 ; 
    wire ptw_l2_pte_x = ptw__GEN_7 ; 
    wire ptw_l2_pte_w = ptw__GEN_8 ; 
    wire ptw_l2_pte_r = ptw__GEN_9 ; 
    wire ptw_l2_pte_v = ptw__GEN_10 ; 
    wire[9:0] ptw_r_pte_pte_reserved_for_future = ptw_l2_pte_reserved_for_future ; 
    wire[9:0] ptw_r_pte_pte_1_reserved_for_future = ptw_l2_pte_reserved_for_future ; 
    wire[1:0] ptw_r_pte_pte_reserved_for_software = ptw_l2_pte_reserved_for_software ; 
    wire[1:0] ptw_r_pte_pte_1_reserved_for_software = ptw_l2_pte_reserved_for_software ; 
    wire ptw_r_pte_pte_d = ptw_l2_pte_d ; 
    wire ptw_r_pte_pte_1_d = ptw_l2_pte_d ; 
    wire ptw_r_pte_pte_a = ptw_l2_pte_a ; 
    wire ptw_r_pte_pte_1_a = ptw_l2_pte_a ; 
    wire ptw_r_pte_pte_g = ptw_l2_pte_g ; 
    wire ptw_r_pte_pte_1_g = ptw_l2_pte_g ; 
    wire ptw_r_pte_pte_u = ptw_l2_pte_u ; 
    wire ptw_r_pte_pte_1_u = ptw_l2_pte_u ; 
    wire ptw_r_pte_pte_x = ptw_l2_pte_x ; 
    wire ptw_r_pte_pte_1_x = ptw_l2_pte_x ; 
    wire ptw_r_pte_pte_w = ptw_l2_pte_w ; 
    wire ptw_r_pte_pte_1_w = ptw_l2_pte_w ; 
    wire ptw_r_pte_pte_r = ptw_l2_pte_r ; 
    wire ptw_r_pte_pte_1_r = ptw_l2_pte_r ; 
    wire ptw_r_pte_pte_v = ptw_l2_pte_v ; 
    wire ptw_r_pte_pte_1_v = ptw_l2_pte_v ; 
    wire[55:0] ptw__GEN_66 ={ ptw_r_pte_ppn ,12'h0}; 
    wire ptw_pmaPgLevelHomogeneous_1 =({1'h0, ptw__GEN_66 ^56'hC000000}&57'h1FFFFFFFC000000)==57'h0|1'h0|({1'h0, ptw__GEN_66 ^56'h60000000}&57'h1FFFFFFE0000000)==57'h0|({1'h0, ptw__GEN_66 ^56'h80000000}&57'h1FFFFFFF0000000)==57'h0; 
    wire[55:0] ptw__GEN_67 ={ ptw_r_pte_ppn ,12'h0}; 
    wire ptw_pmaPgLevelHomogeneous_2 =({1'h0, ptw__GEN_67 }&57'h1FFFFFFFFFFF000)==57'h0|1'h0|({1'h0, ptw__GEN_67 ^56'h3000}&57'h1FFFFFFFFFFF000)==57'h0|({1'h0, ptw__GEN_67 ^56'h10000}&57'h1FFFFFFFFFF0000)==57'h0|({1'h0, ptw__GEN_67 ^56'h2000000}&57'h1FFFFFFFFFF0000)==57'h0|({1'h0, ptw__GEN_67 ^56'hC000000}&57'h1FFFFFFFC000000)==57'h0|({1'h0, ptw__GEN_67 ^56'h60000000}&57'h1FFFFFFE0000000)==57'h0|({1'h0, ptw__GEN_67 ^56'h80000000}&57'h1FFFFFFF0000000)==57'h0; 
    wire ptw_pmaHomogeneous =(& ptw_count ) ?  ptw_pmaPgLevelHomogeneous_2 : ptw_count ==2'h2 ?  ptw_pmaPgLevelHomogeneous_2 : ptw_count ==2'h1 ?  ptw_pmaPgLevelHomogeneous_1 :1'h0; 
    wire[55:0] ptw__GEN_68 ={ ptw_r_pte_ppn ,12'h0}; 
    wire ptw_pmpHomogeneous_maskHomogeneous =(& ptw_count ) ?  ptw_io_dpath_pmp_0_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_0_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_0_mask [20]: ptw_io_dpath_pmp_0_mask [29]; 
    wire[55:0] ptw__GEN_69 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_70 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_71 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_72 =|( ptw__GEN_71 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower = ptw__GEN_68 <{24'h0,~(~{ ptw__pmpHomogeneous_WIRE_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask })<{24'h0,~(~{ ptw__pmpHomogeneous_WIRE_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask })<{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_1 =(& ptw_count ) ?  ptw_io_dpath_pmp_1_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_1_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_1_mask [20]: ptw_io_dpath_pmp_1_mask [29]; 
    wire[55:0] ptw__GEN_73 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_74 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_75 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_76 =|( ptw__GEN_75 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_1 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_1 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_1 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_1 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_1 })<{24'h0,~(~{ ptw_io_dpath_pmp_0_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_1 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_1 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_1 })<{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_1 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_2 =(& ptw_count ) ?  ptw_io_dpath_pmp_2_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_2_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_2_mask [20]: ptw_io_dpath_pmp_2_mask [29]; 
    wire[55:0] ptw__GEN_77 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_78 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_79 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_80 =|( ptw__GEN_79 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_2 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_2 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_2 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_2 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_2 })<{24'h0,~(~{ ptw_io_dpath_pmp_1_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_2 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_2 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_2 })<{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_2 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_3 =(& ptw_count ) ?  ptw_io_dpath_pmp_3_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_3_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_3_mask [20]: ptw_io_dpath_pmp_3_mask [29]; 
    wire[55:0] ptw__GEN_81 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_82 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_83 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_84 =|( ptw__GEN_83 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_3 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_3 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_3 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_3 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_3 })<{24'h0,~(~{ ptw_io_dpath_pmp_2_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_3 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_3 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_3 })<{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_3 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_4 =(& ptw_count ) ?  ptw_io_dpath_pmp_4_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_4_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_4_mask [20]: ptw_io_dpath_pmp_4_mask [29]; 
    wire[55:0] ptw__GEN_85 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_86 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_87 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_88 =|( ptw__GEN_87 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_4 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_4 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_4 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_4 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_4 })<{24'h0,~(~{ ptw_io_dpath_pmp_3_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_4 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_4 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_4 })<{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_4 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_5 =(& ptw_count ) ?  ptw_io_dpath_pmp_5_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_5_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_5_mask [20]: ptw_io_dpath_pmp_5_mask [29]; 
    wire[55:0] ptw__GEN_89 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_90 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_91 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_92 =|( ptw__GEN_91 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_5 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_5 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_5 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_5 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_5 })<{24'h0,~(~{ ptw_io_dpath_pmp_4_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_5 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_5 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_5 })<{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_5 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_6 =(& ptw_count ) ?  ptw_io_dpath_pmp_6_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_6_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_6_mask [20]: ptw_io_dpath_pmp_6_mask [29]; 
    wire[55:0] ptw__GEN_93 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_94 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_95 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_96 =|( ptw__GEN_95 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_6 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_6 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_6 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_6 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_6 })<{24'h0,~(~{ ptw_io_dpath_pmp_5_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_6 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_6 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_6 })<{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_6 }; 
    wire ptw_pmpHomogeneous_maskHomogeneous_7 =(& ptw_count ) ?  ptw_io_dpath_pmp_7_mask [11]: ptw_count ==2'h2 ?  ptw_io_dpath_pmp_7_mask [11]: ptw_count ==2'h1 ?  ptw_io_dpath_pmp_7_mask [20]: ptw_io_dpath_pmp_7_mask [29]; 
    wire[55:0] ptw__GEN_97 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_7_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_98 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_7_addr ,2'h0}|32'h3)}; 
    wire[55:0] ptw__GEN_99 = ptw__GEN_68 ^{24'h0,~(~{ ptw_io_dpath_pmp_7_addr ,2'h0}|32'h3)}; 
    wire ptw__GEN_100 =|( ptw__GEN_99 [55:12]); 
    wire ptw_pmpHomogeneous_beginsAfterLower_7 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)}==1'h0; 
    wire ptw_pmpHomogeneous_beginsAfterUpper_7 = ptw__GEN_68 <{24'h0,~(~{ ptw_io_dpath_pmp_7_addr ,2'h0}|32'h3)}==1'h0; 
    wire[31:0] ptw_pmpHomogeneous_pgMask_7 =(& ptw_count ) ? 32'hFFFFF000: ptw_count ==2'h2 ? 32'hFFFFF000: ptw_count ==2'h1 ? 32'hFFE00000:32'hC0000000; 
    wire ptw_pmpHomogeneous_endsBeforeLower_7 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_7 })<{24'h0,~(~{ ptw_io_dpath_pmp_6_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_7 }; 
    wire ptw_pmpHomogeneous_endsBeforeUpper_7 =( ptw__GEN_68 &{24'h0, ptw_pmpHomogeneous_pgMask_7 })<{24'h0,~(~{ ptw_io_dpath_pmp_7_addr ,2'h0}|32'h3)& ptw_pmpHomogeneous_pgMask_7 }; 
    wire ptw_pmpHomogeneous =( ptw_io_dpath_pmp_0_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous |((& ptw_count ) ?  ptw__GEN_72 : ptw_count ==2'h2 ?  ptw__GEN_72 : ptw_count ==2'h1 ? (|( ptw__GEN_70 [55:21])):(|( ptw__GEN_69 [55:30]))): ptw_io_dpath_pmp_0_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower | ptw_pmpHomogeneous_beginsAfterUpper | ptw_pmpHomogeneous_beginsAfterLower & ptw_pmpHomogeneous_endsBeforeUpper )&1'h1&( ptw_io_dpath_pmp_1_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_1 |((& ptw_count ) ?  ptw__GEN_76 : ptw_count ==2'h2 ?  ptw__GEN_76 : ptw_count ==2'h1 ? (|( ptw__GEN_74 [55:21])):(|( ptw__GEN_73 [55:30]))): ptw_io_dpath_pmp_1_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_1 | ptw_pmpHomogeneous_beginsAfterUpper_1 | ptw_pmpHomogeneous_beginsAfterLower_1 & ptw_pmpHomogeneous_endsBeforeUpper_1 )&( ptw_io_dpath_pmp_2_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_2 |((& ptw_count ) ?  ptw__GEN_80 : ptw_count ==2'h2 ?  ptw__GEN_80 : ptw_count ==2'h1 ? (|( ptw__GEN_78 [55:21])):(|( ptw__GEN_77 [55:30]))): ptw_io_dpath_pmp_2_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_2 | ptw_pmpHomogeneous_beginsAfterUpper_2 | ptw_pmpHomogeneous_beginsAfterLower_2 & ptw_pmpHomogeneous_endsBeforeUpper_2 )&( ptw_io_dpath_pmp_3_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_3 |((& ptw_count ) ?  ptw__GEN_84 : ptw_count ==2'h2 ?  ptw__GEN_84 : ptw_count ==2'h1 ? (|( ptw__GEN_82 [55:21])):(|( ptw__GEN_81 [55:30]))): ptw_io_dpath_pmp_3_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_3 | ptw_pmpHomogeneous_beginsAfterUpper_3 | ptw_pmpHomogeneous_beginsAfterLower_3 & ptw_pmpHomogeneous_endsBeforeUpper_3 )&( ptw_io_dpath_pmp_4_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_4 |((& ptw_count ) ?  ptw__GEN_88 : ptw_count ==2'h2 ?  ptw__GEN_88 : ptw_count ==2'h1 ? (|( ptw__GEN_86 [55:21])):(|( ptw__GEN_85 [55:30]))): ptw_io_dpath_pmp_4_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_4 | ptw_pmpHomogeneous_beginsAfterUpper_4 | ptw_pmpHomogeneous_beginsAfterLower_4 & ptw_pmpHomogeneous_endsBeforeUpper_4 )&( ptw_io_dpath_pmp_5_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_5 |((& ptw_count ) ?  ptw__GEN_92 : ptw_count ==2'h2 ?  ptw__GEN_92 : ptw_count ==2'h1 ? (|( ptw__GEN_90 [55:21])):(|( ptw__GEN_89 [55:30]))): ptw_io_dpath_pmp_5_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_5 | ptw_pmpHomogeneous_beginsAfterUpper_5 | ptw_pmpHomogeneous_beginsAfterLower_5 & ptw_pmpHomogeneous_endsBeforeUpper_5 )&( ptw_io_dpath_pmp_6_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_6 |((& ptw_count ) ?  ptw__GEN_96 : ptw_count ==2'h2 ?  ptw__GEN_96 : ptw_count ==2'h1 ? (|( ptw__GEN_94 [55:21])):(|( ptw__GEN_93 [55:30]))): ptw_io_dpath_pmp_6_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_6 | ptw_pmpHomogeneous_beginsAfterUpper_6 | ptw_pmpHomogeneous_beginsAfterLower_6 & ptw_pmpHomogeneous_endsBeforeUpper_6 )&( ptw_io_dpath_pmp_7_cfg_a [1] ?  ptw_pmpHomogeneous_maskHomogeneous_7 |((& ptw_count ) ?  ptw__GEN_100 : ptw_count ==2'h2 ?  ptw__GEN_100 : ptw_count ==2'h1 ? (|( ptw__GEN_98 [55:21])):(|( ptw__GEN_97 [55:30]))): ptw_io_dpath_pmp_7_cfg_a [0]==1'h0| ptw_pmpHomogeneous_endsBeforeLower_7 | ptw_pmpHomogeneous_beginsAfterUpper_7 | ptw_pmpHomogeneous_beginsAfterLower_7 & ptw_pmpHomogeneous_endsBeforeUpper_7 ); 
    wire ptw_homogeneous = ptw_pmaHomogeneous & ptw_pmpHomogeneous ; 
    wire ptw_io_requestor_0_resp_bits_gpa_bits_truncIdx = ptw_aux_count [0]; 
    wire[55:0] ptw__GEN_101 ={ ptw_stage2_final ==1'h0| ptw_r_req_vstage1 ==1'h0| ptw_aux_count ==2'h2 ?  ptw_aux_pte_ppn :(& ptw_io_requestor_0_resp_bits_gpa_bits_truncIdx ) ? { ptw_aux_pte_ppn [43:9], ptw_r_req_addr [8:0]}:{ ptw_aux_pte_ppn [43:18], ptw_r_req_addr [17:0]}, ptw_gpa_pgoff }; 
    wire ptw_io_requestor_1_resp_bits_gpa_bits_truncIdx = ptw_aux_count [0]; 
    wire[55:0] ptw__GEN_102 ={ ptw_stage2_final ==1'h0| ptw_r_req_vstage1 ==1'h0| ptw_aux_count ==2'h2 ?  ptw_aux_pte_ppn :(& ptw_io_requestor_1_resp_bits_gpa_bits_truncIdx ) ? { ptw_aux_pte_ppn [43:9], ptw_r_req_addr [8:0]}:{ ptw_aux_pte_ppn [43:18], ptw_r_req_addr [17:0]}, ptw_gpa_pgoff }; 
    wire[2:0] ptw_next_state ;  
    wire ptw_state_barrier_clock;
    wire ptw_state_barrier_reset;
    wire[2:0] ptw_state_barrier_io_x;
    wire[2:0] ptw_state_barrier_io_y;

    assign  ptw_state_barrier_io_y = ptw_state_barrier_io_x ;
    assign ptw_state_barrier_clock = ptw_clock;
    assign ptw_state_barrier_reset = ptw_reset;
    assign ptw_state_barrier_io_x = ptw_next_state;
    assign ptw__state_barrier_io_y = ptw_state_barrier_io_y;
     
    wire ptw__GEN_103 =3'h0== ptw_state ; 
    wire ptw__GEN_104 = ptw__GEN & ptw__arb_io_out_valid ; 
    wire[43:0] ptw_aux_ppn = ptw__arb_io_out_bits_bits_vstage1  ?  ptw_io_dpath_vsatp_ppn :{23'h0, ptw__arb_io_out_bits_bits_addr }; 
    wire ptw__GEN_105 = ptw__GEN_103  ? ( ptw__GEN_104  ?  ptw__arb_io_out_bits_bits_stage2 : ptw_stage2 ): ptw_stage2 ; 
    wire ptw__GEN_106 = ptw__arb_io_out_bits_bits_stage2 & ptw__arb_io_out_bits_bits_vstage1 ==1'h0; 
    wire ptw__GEN_107 = ptw__GEN_103  ? ( ptw__GEN_104  ?  ptw__GEN_106 : ptw_stage2_final ): ptw_stage2_final ; 
    wire[1:0] ptw__GEN_108 = ptw__arb_io_out_bits_bits_stage2  ?  ptw_hgatp_initial_count : ptw_satp_initial_count ; 
    wire[1:0] ptw__GEN_109 = ptw__arb_io_out_bits_bits_vstage1  ?  ptw_vsatp_initial_count :2'h0; 
    wire ptw__GEN_110 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h0: ptw_resp_ae_final ): ptw_resp_ae_final ; 
    wire ptw__GEN_111 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h0: ptw_resp_pf ): ptw_resp_pf ; 
    wire[14:0] ptw_resp_gf_idxs_0 = ptw_aux_ppn [43:29]; 
    wire[14:0] ptw__resp_gf_WIRE_0 = ptw_resp_gf_idxs_0 ; 
    wire ptw__GEN_112 =(| ptw__resp_gf_WIRE_0 )& ptw__arb_io_out_bits_bits_stage2 ; 
    wire ptw__GEN_113 = ptw__GEN_103  ? ( ptw__GEN_104  ?  ptw__GEN_112 : ptw_resp_gf ): ptw_resp_gf ; 
    wire ptw__GEN_114 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h1: ptw_resp_hr ): ptw_resp_hr ; 
    wire ptw__GEN_115 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h1: ptw_resp_hw ): ptw_resp_hw ; 
    wire ptw__GEN_116 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h1: ptw_resp_hx ): ptw_resp_hx ; 
    wire ptw__GEN_117 =( ptw__arb_io_out_bits_bits_need_gpa ==1'h0| ptw__arb_io_out_bits_bits_stage2 )==1'h0; 
    wire ptw__GEN_118 =~ ptw__GEN_103 ; 
    wire ptw__GEN_119 =3'h1== ptw_state ; 
    wire ptw__GEN_120 = ptw__GEN_118 & ptw__GEN_119 ; 
    wire ptw__GEN_121 = ptw_stage2 & ptw_count == ptw_r_hgatp_initial_count ; 
    wire[23:0] ptw__GEN_122 = ptw_aux_count ==2'h2 ? { ptw_r_req_addr ,3'h0}:24'h0; 
    wire[2:0] ptw__GEN_123 ={1'h0, ptw_aux_count }+3'h1; 
    wire[43:0] ptw__GEN_124 ={24'h0, ptw_stage2_pte_cache_data }; 
    wire ptw__GEN_125 = ptw__GEN_120 &~ ptw_stage2_pte_cache_hit ; 
    wire[2:0] ptw__GEN_126 ={1'h0, ptw_count }+3'h1; 
    wire ptw__GEN_127 = ptw__GEN_120 & ptw_resp_gf ; 
    wire ptw__GEN_128 = ptw_r_req_dest ==1'h0; 
    wire ptw__GEN_129 =& ptw_r_req_dest ; 
    wire ptw__GEN_130 = ptw__GEN_118 &~ ptw__GEN_119 ; 
    wire ptw__GEN_131 =3'h2== ptw_state ; 
    wire ptw__GEN_132 = ptw__GEN_130 &~ ptw__GEN_131 ; 
    wire ptw__GEN_133 =3'h4== ptw_state ; 
  assign  ptw__io_dpath_perf_pte_miss_output = ptw__GEN_103  ? 1'h0: ptw__GEN_119  ? 1'h0: ptw__GEN_131  ? 1'h0: ptw__GEN_133  ?  ptw_count <2'h2:1'h0; 
    wire ptw__GEN_134 = ptw__GEN_132 & ptw__GEN_133 & ptw_io_mem_s2_xcpt_ae_ld ; 
    wire ptw__GEN_135 = ptw__GEN_103  ? ( ptw__GEN_104  ? 1'h0: ptw_resp_ae_ptw ): ptw__GEN_119  ?  ptw_resp_ae_ptw : ptw__GEN_131  ?  ptw_resp_ae_ptw : ptw__GEN_133  ? ( ptw_io_mem_s2_xcpt_ae_ld  ? 1'h1: ptw_resp_ae_ptw ): ptw_resp_ae_ptw ; 
    wire ptw__GEN_136 = ptw_r_req_dest ==1'h0; 
    wire ptw__GEN_137 =& ptw_r_req_dest ; 
    wire ptw__GEN_138 =3'h7== ptw_state ; 
    wire ptw__GEN_139 = ptw__GEN_132 &~ ptw__GEN_133 & ptw__GEN_138 ; 
    wire ptw__GEN_140 = ptw_r_req_dest ==1'h0; 
    wire ptw__GEN_141 = ptw__GEN_103  ?  ptw__resp_valid_WIRE_0 : ptw__GEN_119  ? ( ptw_resp_gf  ? ( ptw__GEN_128  ? 1'h1: ptw__resp_valid_WIRE_0 ): ptw__resp_valid_WIRE_0 ): ptw__GEN_131  ?  ptw__resp_valid_WIRE_0 : ptw__GEN_133  ? ( ptw_io_mem_s2_xcpt_ae_ld  ? ( ptw__GEN_136  ? 1'h1: ptw__resp_valid_WIRE_0 ): ptw__resp_valid_WIRE_0 ): ptw__GEN_138  ? ( ptw__GEN_140  ? 1'h1: ptw__resp_valid_WIRE_0 ): ptw__resp_valid_WIRE_0 ; 
    wire ptw__GEN_142 =& ptw_r_req_dest ; 
    wire ptw__GEN_143 = ptw__GEN_103  ?  ptw__resp_valid_WIRE_1 : ptw__GEN_119  ? ( ptw_resp_gf  ? ( ptw__GEN_129  ? 1'h1: ptw__resp_valid_WIRE_1 ): ptw__resp_valid_WIRE_1 ): ptw__GEN_131  ?  ptw__resp_valid_WIRE_1 : ptw__GEN_133  ? ( ptw_io_mem_s2_xcpt_ae_ld  ? ( ptw__GEN_137  ? 1'h1: ptw__resp_valid_WIRE_1 ): ptw__resp_valid_WIRE_1 ): ptw__GEN_138  ? ( ptw__GEN_142  ? 1'h1: ptw__resp_valid_WIRE_1 ): ptw__resp_valid_WIRE_1 ; 
    wire ptw__GEN_144 = ptw_homogeneous ==1'h0; 
    wire[1:0] ptw__GEN_145 = ptw__GEN_103  ? ( ptw__GEN_104  ?  ptw__GEN_108 : ptw_count ): ptw__GEN_119  ? ( ptw_stage2_pte_cache_hit  ?  ptw_count : ptw_pte_cache_hit  ?  ptw__GEN_126 [1:0]: ptw_count ): ptw__GEN_131  ?  ptw_count : ptw__GEN_133  ?  ptw_count : ptw__GEN_138  ? ( ptw__GEN_144  ? 2'h2: ptw_count ): ptw_count ; 
    wire[1:0] ptw__GEN_146 = ptw_stage2_final  ?  ptw_max_count :2'h2; 
    wire[43:0] ptw_merged_pte_superpage_mask =(& ptw__GEN_146 ) ? 44'hFFFFFFFFFFF: ptw__GEN_146 ==2'h2 ? 44'hFFFFFFFFFFF: ptw__GEN_146 ==2'h1 ? 44'hFFFFFFFFE00:44'hFFFFFFC0000; 
    wire[43:0] ptw_merged_pte_stage1_ppns_0 ={ ptw_pte_ppn [43:18], ptw_aux_pte_ppn [17:0]}; 
    wire[43:0] ptw_merged_pte_stage1_ppns_1 ={ ptw_pte_ppn [43:9], ptw_aux_pte_ppn [8:0]}; 
    wire[43:0] ptw_merged_pte_stage1_ppn =(& ptw_count ) ?  ptw_pte_ppn : ptw_count ==2'h2 ?  ptw_pte_ppn : ptw_count ==2'h1 ?  ptw_merged_pte_stage1_ppns_1 : ptw_merged_pte_stage1_ppns_0 ; 
    wire[43:0] ptw_merged_pte_ppn = ptw_merged_pte_stage1_ppn & ptw_merged_pte_superpage_mask ; 
    wire ptw__GEN_147 = ptw_state ==3'h1& ptw_stage2_pte_cache_hit ; 
    wire[1:0] ptw_r_pte_lsbs ={1'h0, ptw_r_pte_idxs_0 }; 
    wire[43:0] ptw_r_pte_pte_ppn ={ ptw_r_hgatp_ppn [43:2], ptw_r_pte_lsbs }; 
    wire ptw__GEN_148 = ptw_state ==3'h1& ptw_pte_cache_hit ; 
    wire[43:0] ptw_r_pte_pte_1_ppn ={24'h0, ptw_pte_cache_data }; 
    wire[16:0] ptw_r_pte_idxs_0_1 = ptw_pte_ppn [43:27]; 
    wire[1:0] ptw_r_pte_lsbs_1 = ptw_r_pte_idxs_0_1 [1:0]; 
    wire[43:0] ptw_r_pte_pte_2_ppn ={ ptw_r_hgatp_ppn [43:2], ptw_r_pte_lsbs_1 }; 
    wire ptw__GEN_149 = ptw_traverse ==1'h0& ptw_r_req_vstage1 & ptw_stage2 ; 
    wire ptw__GEN_150 =(& ptw_state )& ptw_homogeneous ==1'h0& ptw_count !=2'h2; 
    wire ptw_r_pte_truncIdx = ptw_count [0]; 
    wire[43:0] ptw_r_pte_pte_3_ppn =(& ptw_r_pte_truncIdx ) ? { ptw_r_pte_ppn [43:9], ptw_r_req_addr [8:0]}:{ ptw_r_pte_ppn [43:18], ptw_r_req_addr [17:0]}; 
    wire ptw__GEN_151 = ptw__GEN & ptw__arb_io_out_valid ; 
    wire[16:0] ptw_r_pte_idxs_0_2 = ptw_io_dpath_vsatp_ppn [43:27]; 
    wire[1:0] ptw_r_pte_lsbs_2 = ptw_r_pte_idxs_0_2 [1:0]; 
    wire[43:0] ptw_r_pte_pte_4_ppn ={ ptw_io_dpath_hgatp_ppn [43:2], ptw_r_pte_lsbs_2 }; 
    wire ptw_do_switch ;  
    wire ptw_r_pte_barrier_clock;
    wire ptw_r_pte_barrier_reset;
    wire[9:0] ptw_r_pte_barrier_io_x_reserved_for_future;
    wire[43:0] ptw_r_pte_barrier_io_x_ppn;
    wire[1:0] ptw_r_pte_barrier_io_x_reserved_for_software;
    wire ptw_r_pte_barrier_io_x_d;
    wire ptw_r_pte_barrier_io_x_a;
    wire ptw_r_pte_barrier_io_x_g;
    wire ptw_r_pte_barrier_io_x_u;
    wire ptw_r_pte_barrier_io_x_x;
    wire ptw_r_pte_barrier_io_x_w;
    wire ptw_r_pte_barrier_io_x_r;
    wire ptw_r_pte_barrier_io_x_v;
    wire[9:0] ptw_r_pte_barrier_io_y_reserved_for_future;
    wire[43:0] ptw_r_pte_barrier_io_y_ppn;
    wire[1:0] ptw_r_pte_barrier_io_y_reserved_for_software;
    wire ptw_r_pte_barrier_io_y_d;
    wire ptw_r_pte_barrier_io_y_a;
    wire ptw_r_pte_barrier_io_y_g;
    wire ptw_r_pte_barrier_io_y_u;
    wire ptw_r_pte_barrier_io_y_x;
    wire ptw_r_pte_barrier_io_y_w;
    wire ptw_r_pte_barrier_io_y_r;
    wire ptw_r_pte_barrier_io_y_v;

    assign  ptw_r_pte_barrier_io_y_reserved_for_future = ptw_r_pte_barrier_io_x_reserved_for_future ; 
  assign  ptw_r_pte_barrier_io_y_ppn = ptw_r_pte_barrier_io_x_ppn ; 
  assign  ptw_r_pte_barrier_io_y_reserved_for_software = ptw_r_pte_barrier_io_x_reserved_for_software ; 
  assign  ptw_r_pte_barrier_io_y_d = ptw_r_pte_barrier_io_x_d ; 
  assign  ptw_r_pte_barrier_io_y_a = ptw_r_pte_barrier_io_x_a ; 
  assign  ptw_r_pte_barrier_io_y_g = ptw_r_pte_barrier_io_x_g ; 
  assign  ptw_r_pte_barrier_io_y_u = ptw_r_pte_barrier_io_x_u ; 
  assign  ptw_r_pte_barrier_io_y_x = ptw_r_pte_barrier_io_x_x ; 
  assign  ptw_r_pte_barrier_io_y_w = ptw_r_pte_barrier_io_x_w ; 
  assign  ptw_r_pte_barrier_io_y_r = ptw_r_pte_barrier_io_x_r ; 
  assign  ptw_r_pte_barrier_io_y_v = ptw_r_pte_barrier_io_x_v ;
    assign ptw_r_pte_barrier_clock = ptw_clock;
    assign ptw_r_pte_barrier_reset = ptw_reset;
    assign ptw_r_pte_barrier_io_x_reserved_for_future = ptw__GEN_147 ? ptw_r_pte_pte_reserved_for_future:ptw__GEN_148 ? ptw_r_pte_pte_1_reserved_for_future:ptw_do_switch ? ptw_r_pte_pte_2_reserved_for_future:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_reserved_for_future:ptw_pte_reserved_for_future):ptw__GEN_150 ? ptw_r_pte_pte_3_reserved_for_future:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_reserved_for_future:ptw_r_pte_pte_5_reserved_for_future):ptw_r_pte_reserved_for_future;
    assign ptw_r_pte_barrier_io_x_ppn = ptw__GEN_147 ? ptw_r_pte_pte_ppn:ptw__GEN_148 ? ptw_r_pte_pte_1_ppn:ptw_do_switch ? ptw_r_pte_pte_2_ppn:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_ppn:ptw_pte_ppn):ptw__GEN_150 ? ptw_r_pte_pte_3_ppn:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_ppn:ptw_r_pte_pte_5_ppn):ptw_r_pte_ppn;
    assign ptw_r_pte_barrier_io_x_reserved_for_software = ptw__GEN_147 ? ptw_r_pte_pte_reserved_for_software:ptw__GEN_148 ? ptw_r_pte_pte_1_reserved_for_software:ptw_do_switch ? ptw_r_pte_pte_2_reserved_for_software:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_reserved_for_software:ptw_pte_reserved_for_software):ptw__GEN_150 ? ptw_r_pte_pte_3_reserved_for_software:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_reserved_for_software:ptw_r_pte_pte_5_reserved_for_software):ptw_r_pte_reserved_for_software;
    assign ptw_r_pte_barrier_io_x_d = ptw__GEN_147 ? ptw_r_pte_pte_d:ptw__GEN_148 ? ptw_r_pte_pte_1_d:ptw_do_switch ? ptw_r_pte_pte_2_d:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_d:ptw_pte_d):ptw__GEN_150 ? ptw_r_pte_pte_3_d:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_d:ptw_r_pte_pte_5_d):ptw_r_pte_d;
    assign ptw_r_pte_barrier_io_x_a = ptw__GEN_147 ? ptw_r_pte_pte_a:ptw__GEN_148 ? ptw_r_pte_pte_1_a:ptw_do_switch ? ptw_r_pte_pte_2_a:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_a:ptw_pte_a):ptw__GEN_150 ? ptw_r_pte_pte_3_a:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_a:ptw_r_pte_pte_5_a):ptw_r_pte_a;
    assign ptw_r_pte_barrier_io_x_g = ptw__GEN_147 ? ptw_r_pte_pte_g:ptw__GEN_148 ? ptw_r_pte_pte_1_g:ptw_do_switch ? ptw_r_pte_pte_2_g:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_g:ptw_pte_g):ptw__GEN_150 ? ptw_r_pte_pte_3_g:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_g:ptw_r_pte_pte_5_g):ptw_r_pte_g;
    assign ptw_r_pte_barrier_io_x_u = ptw__GEN_147 ? ptw_r_pte_pte_u:ptw__GEN_148 ? ptw_r_pte_pte_1_u:ptw_do_switch ? ptw_r_pte_pte_2_u:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_u:ptw_pte_u):ptw__GEN_150 ? ptw_r_pte_pte_3_u:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_u:ptw_r_pte_pte_5_u):ptw_r_pte_u;
    assign ptw_r_pte_barrier_io_x_x = ptw__GEN_147 ? ptw_r_pte_pte_x:ptw__GEN_148 ? ptw_r_pte_pte_1_x:ptw_do_switch ? ptw_r_pte_pte_2_x:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_x:ptw_pte_x):ptw__GEN_150 ? ptw_r_pte_pte_3_x:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_x:ptw_r_pte_pte_5_x):ptw_r_pte_x;
    assign ptw_r_pte_barrier_io_x_w = ptw__GEN_147 ? ptw_r_pte_pte_w:ptw__GEN_148 ? ptw_r_pte_pte_1_w:ptw_do_switch ? ptw_r_pte_pte_2_w:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_w:ptw_pte_w):ptw__GEN_150 ? ptw_r_pte_pte_3_w:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_w:ptw_r_pte_pte_5_w):ptw_r_pte_w;
    assign ptw_r_pte_barrier_io_x_r = ptw__GEN_147 ? ptw_r_pte_pte_r:ptw__GEN_148 ? ptw_r_pte_pte_1_r:ptw_do_switch ? ptw_r_pte_pte_2_r:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_r:ptw_pte_r):ptw__GEN_150 ? ptw_r_pte_pte_3_r:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_r:ptw_r_pte_pte_5_r):ptw_r_pte_r;
    assign ptw_r_pte_barrier_io_x_v = ptw__GEN_147 ? ptw_r_pte_pte_v:ptw__GEN_148 ? ptw_r_pte_pte_1_v:ptw_do_switch ? ptw_r_pte_pte_2_v:ptw_mem_resp_valid ? (ptw__GEN_149 ? ptw_merged_pte_v:ptw_pte_v):ptw__GEN_150 ? ptw_r_pte_pte_3_v:ptw__GEN_151 ? (ptw__arb_io_out_bits_bits_stage2 ? ptw_r_pte_pte_4_v:ptw_r_pte_pte_5_v):ptw_r_pte_v;
    assign ptw__r_pte_barrier_io_y_reserved_for_future = ptw_r_pte_barrier_io_y_reserved_for_future;
    assign ptw__r_pte_barrier_io_y_ppn = ptw_r_pte_barrier_io_y_ppn;
    assign ptw__r_pte_barrier_io_y_reserved_for_software = ptw_r_pte_barrier_io_y_reserved_for_software;
    assign ptw__r_pte_barrier_io_y_d = ptw_r_pte_barrier_io_y_d;
    assign ptw__r_pte_barrier_io_y_a = ptw_r_pte_barrier_io_y_a;
    assign ptw__r_pte_barrier_io_y_g = ptw_r_pte_barrier_io_y_g;
    assign ptw__r_pte_barrier_io_y_u = ptw_r_pte_barrier_io_y_u;
    assign ptw__r_pte_barrier_io_y_x = ptw_r_pte_barrier_io_y_x;
    assign ptw__r_pte_barrier_io_y_w = ptw_r_pte_barrier_io_y_w;
    assign ptw__r_pte_barrier_io_y_r = ptw_r_pte_barrier_io_y_r;
    assign ptw__r_pte_barrier_io_y_v = ptw_r_pte_barrier_io_y_v;
     
    wire ptw__GEN_152 = ptw_state ==3'h5==1'h0; 
    wire ptw__GEN_153 = ptw_do_both_stages & ptw_stage2 ==1'h0; 
    wire[2:0] ptw__GEN_154 ={1'h0, ptw_count }+3'h1; 
    wire ptw__GEN_155 = ptw_mem_resp_valid &~ ptw_traverse ; 
    wire ptw_gf = ptw_stage2 & ptw_stage2_final ==1'h0&( ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_r & ptw_pte_u )==1'h0; 
    wire ptw_ae = ptw_pte_v & ptw_invalid_paddr ; 
    wire ptw_pf = ptw_pte_v &(| ptw_pte_reserved_for_future ); 
    wire ptw_success = ptw_pte_v & ptw_ae ==1'h0& ptw_pf ==1'h0& ptw_gf ==1'h0; 
    wire ptw__GEN_156 = ptw_do_both_stages & ptw_stage2_final ==1'h0& ptw_success ; 
    wire ptw__GEN_157 = ptw__GEN_155 & ptw__GEN_156 ; 
  assign  ptw_do_switch = ptw_mem_resp_valid  ? ( ptw_traverse  ?  ptw__GEN_153 : ptw__GEN_156  ? ( ptw_stage2  ? 1'h0:1'h1):1'h0):1'h0; 
    wire ptw__GEN_158 = ptw__GEN_155 &~ ptw__GEN_156 ; 
    wire ptw__GEN_159 = ptw_r_req_dest ==1'h0; 
    wire ptw__GEN_160 =& ptw_r_req_dest ; 
    wire ptw__GEN_161 = ptw_ae & ptw_count <2'h2& ptw_pte_v & ptw_pte_r ==1'h0& ptw_pte_w ==1'h0& ptw_pte_x ==1'h0& ptw_pte_d ==1'h0& ptw_pte_a ==1'h0& ptw_pte_u ==1'h0& ptw_pte_reserved_for_future ==10'h0; 
    wire ptw__GEN_162 = ptw_pf & ptw_stage2 ==1'h0; 
    wire ptw__GEN_163 = ptw_gf | ptw_pf & ptw_stage2 ; 
    wire ptw__GEN_164 = ptw_stage2 ==1'h0| ptw_pf ==1'h0& ptw_gf ==1'h0& ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_r & ptw_pte_u ; 
    wire ptw__GEN_165 = ptw_stage2 ==1'h0| ptw_pf ==1'h0& ptw_gf ==1'h0& ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_w & ptw_pte_d & ptw_pte_u ; 
    wire ptw__GEN_166 = ptw_stage2 ==1'h0| ptw_pf ==1'h0& ptw_gf ==1'h0& ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_x & ptw_pte_u ; 
    wire ptw__GEN_167 = ptw_state ==3'h4==1'h0; 
  always @( posedge  ptw_clock )
         begin 
             if ( ptw_reset ==1'h0& ptw__GEN_65 )
                 begin 
                     if (1)$error("Assertion failed: PTE Cache Hit/Miss Performance Monitor Events are lower priority than L2TLB Hit event\n    at PTW.scala:395 assert(!(io.dpath.perf.l2hit && (io.dpath.perf.pte_miss || io.dpath.perf.pte_hit)),\n");
                     if (1)$fatal;
                 end 
             if ( ptw__GEN_103 & ptw__GEN_104 & ptw_reset ==1'h0& ptw__GEN_117 )
                 begin 
                     if (1)$error("Assertion failed\n    at PTW.scala:609 assert(!arb.io.out.bits.bits.need_gpa || arb.io.out.bits.bits.stage2)\n");
                     if (1)$fatal;
                 end 
             if (1'h0)
                 begin 
                     if (1)$error("Assertion failed\n    at PTW.scala:685 assert(state === s_req || state === s_wait1)\n");
                     if (1)$fatal;
                 end 
             if ( ptw_mem_resp_valid & ptw_reset ==1'h0& ptw__GEN_152 )
                 begin 
                     if (1)$error("Assertion failed\n    at PTW.scala:691 assert(state === s_wait3)\n");
                     if (1)$fatal;
                 end 
             if ( ptw_io_mem_s2_nack & ptw_reset ==1'h0& ptw__GEN_167 )
                 begin 
                     if (1)$error("Assertion failed\n    at PTW.scala:735 assert(state === s_wait2)\n");
                     if (1)$fatal;
                 end 
         end
  assign  ptw_next_state = ptw_io_mem_s2_nack  ? 3'h1: ptw_mem_resp_valid  ? ( ptw_traverse  ? 3'h1: ptw__GEN_156  ? 3'h1:3'h0): ptw__GEN_103  ? ( ptw__GEN_104  ? ( ptw__arb_io_out_bits_valid  ? 3'h1:3'h0): ptw_state ): ptw__GEN_119  ? ( ptw_resp_gf  ? 3'h0: ptw_stage2_pte_cache_hit  ?  ptw_state : ptw_pte_cache_hit  ?  ptw_state : ptw_io_mem_req_ready  ? 3'h2:3'h1): ptw__GEN_131  ? 3'h4: ptw__GEN_133  ? ( ptw_io_mem_s2_xcpt_ae_ld  ? 3'h0:3'h5): ptw__GEN_138  ? 3'h0: ptw_state ; 
    wire[2:0] ptw__GEN_168 ={1'h0, ptw_count }+3'h1; 
    wire[1:0] ptw__GEN_169 = ptw_traverse  ?  ptw__GEN_168 [1:0]: ptw_count ; 
    wire[43:0] ptw_aux_pte_s1_ppns_0 ={ ptw_pte_ppn [43:18], ptw_r_req_addr [17:0]}; 
    wire[43:0] ptw_aux_pte_s1_ppns_1 ={ ptw_pte_ppn [43:9], ptw_r_req_addr [8:0]}; 
    wire[43:0] ptw_aux_pte_pte_ppn =(& ptw_count ) ?  ptw_pte_ppn : ptw_count ==2'h2 ?  ptw_pte_ppn : ptw_count ==2'h1 ?  ptw_aux_pte_s1_ppns_1 : ptw_aux_pte_s1_ppns_0 ; 
    wire[9:0] ptw__GEN_170 = ptw_traverse  ?  ptw_pte_reserved_for_future : ptw_aux_pte_pte_reserved_for_future ; 
    wire[43:0] ptw__GEN_171 = ptw_traverse  ?  ptw_pte_ppn : ptw_aux_pte_pte_ppn ; 
    wire[1:0] ptw__GEN_172 = ptw_traverse  ?  ptw_pte_reserved_for_software : ptw_aux_pte_pte_reserved_for_software ; 
    wire ptw__GEN_173 = ptw_traverse  ?  ptw_pte_d : ptw_aux_pte_pte_d ; 
    wire ptw__GEN_174 = ptw_traverse  ?  ptw_pte_a : ptw_aux_pte_pte_a ; 
    wire ptw__GEN_175 = ptw_traverse  ?  ptw_pte_g : ptw_aux_pte_pte_g ; 
    wire ptw__GEN_176 = ptw_traverse  ?  ptw_pte_u : ptw_aux_pte_pte_u ; 
    wire ptw__GEN_177 = ptw_traverse  ?  ptw_pte_x : ptw_aux_pte_pte_x ; 
    wire ptw__GEN_178 = ptw_traverse  ?  ptw_pte_w : ptw_aux_pte_pte_w ; 
    wire ptw__GEN_179 = ptw_traverse  ?  ptw_pte_r : ptw_aux_pte_pte_r ; 
    wire ptw__GEN_180 = ptw_traverse  ?  ptw_pte_v : ptw_aux_pte_pte_v ; 
    wire ptw_leaf = ptw_mem_resp_valid & ptw_traverse ==1'h0& ptw_count ==2'h0; 
    wire ptw_leaf_1 = ptw_mem_resp_valid & ptw_traverse ==1'h0& ptw_count ==2'h1; 
    wire ptw_leaf_2 = ptw_mem_resp_valid & ptw_traverse ==1'h0& ptw_count ==2'h2; 
  always @( posedge  ptw_clock )
         begin 
             if ( ptw_reset )
                 begin  
                     ptw_state  <=3'h0; 
                     ptw_state_reg  <=7'h0; 
                     ptw_valid  <=8'h0; 
                     ptw_state_reg_1  <=7'h0; 
                     ptw_valid_1  <=8'h0;
                 end 
              else 
                 begin  
                     ptw_state  <= ptw__state_barrier_io_y ;
                     if ( ptw__GEN_35 ) 
                         ptw_state_reg  <= ptw__GEN_38 ;
                      else 
                         if ( ptw__GEN_15 ) 
                             ptw_state_reg  <= ptw__GEN_34 ;
                          else 
                             begin 
                             end 
                     if ( ptw__GEN_39 ) 
                         ptw_valid  <=8'h0;
                      else 
                         if ( ptw__GEN_15 ) 
                             ptw_valid  <= ptw__GEN_17 ;
                          else 
                             begin 
                             end 
                     if ( ptw__GEN_60 ) 
                         ptw_state_reg_1  <= ptw__GEN_63 ;
                      else 
                         if ( ptw__GEN_40 ) 
                             ptw_state_reg_1  <= ptw__GEN_59 ;
                          else 
                             begin 
                             end 
                     if ( ptw__GEN_64 ) 
                         ptw_valid_1  <=8'h0;
                      else 
                         if ( ptw__GEN_40 ) 
                             ptw_valid_1  <= ptw__GEN_42 ;
                          else 
                             begin 
                             end 
                 end 
         end
  always @( posedge  ptw_clock )
         begin  
             ptw_resp_valid_0  <= ptw_mem_resp_valid  ? ( ptw_traverse  ?  ptw__GEN_141 : ptw__GEN_156  ?  ptw__GEN_141 : ptw__GEN_159  ? 1'h1: ptw__GEN_141 ): ptw__GEN_141 ; 
             ptw_resp_valid_1  <= ptw_mem_resp_valid  ? ( ptw_traverse  ?  ptw__GEN_143 : ptw__GEN_156  ?  ptw__GEN_143 : ptw__GEN_160  ? 1'h1: ptw__GEN_143 ): ptw__GEN_143 ; 
             ptw_invalidated  <= ptw_io_dpath_sfence_valid | ptw_invalidated &(| ptw_state );
             if ( ptw_do_switch )
                 begin  
                     ptw_count  <= ptw_r_hgatp_initial_count ; 
                     ptw_aux_count  <= ptw__GEN_169 ; 
                     ptw_aux_pte_reserved_for_future  <= ptw__GEN_170 ; 
                     ptw_aux_pte_ppn  <= ptw__GEN_171 ; 
                     ptw_aux_pte_reserved_for_software  <= ptw__GEN_172 ; 
                     ptw_aux_pte_d  <= ptw__GEN_173 ; 
                     ptw_aux_pte_a  <= ptw__GEN_174 ; 
                     ptw_aux_pte_g  <= ptw__GEN_175 ; 
                     ptw_aux_pte_u  <= ptw__GEN_176 ; 
                     ptw_aux_pte_x  <= ptw__GEN_177 ; 
                     ptw_aux_pte_w  <= ptw__GEN_178 ; 
                     ptw_aux_pte_r  <= ptw__GEN_179 ; 
                     ptw_aux_pte_v  <= ptw__GEN_180 ; 
                     ptw_stage2  <=1'h1;
                 end 
              else 
                 begin 
                     if ( ptw_mem_resp_valid )
                         begin 
                             if ( ptw_traverse )
                                 begin  
                                     ptw_count  <= ptw__GEN_154 [1:0];
                                     if ( ptw__GEN_103 )
                                         begin 
                                             if ( ptw__GEN_104 ) 
                                                 ptw_stage2  <= ptw__arb_io_out_bits_bits_stage2 ;
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else 
                                         begin 
                                         end 
                                 end 
                              else 
                                 if ( ptw__GEN_156 )
                                     begin 
                                         if ( ptw_stage2 )
                                             begin  
                                                 ptw_count  <= ptw_aux_count ; 
                                                 ptw_stage2  <=1'h0;
                                             end 
                                          else 
                                             if ( ptw__GEN_103 )
                                                 begin 
                                                     if ( ptw__GEN_104 )
                                                         begin  
                                                             ptw_count  <= ptw__GEN_108 ; 
                                                             ptw_stage2  <= ptw__arb_io_out_bits_bits_stage2 ;
                                                         end 
                                                      else 
                                                         begin 
                                                         end 
                                                 end 
                                              else 
                                                 if ( ptw__GEN_119 )
                                                     begin 
                                                         if ( ptw_stage2_pte_cache_hit )
                                                             begin 
                                                             end 
                                                          else 
                                                             if ( ptw_pte_cache_hit ) 
                                                                 ptw_count  <= ptw__GEN_126 [1:0];
                                                              else 
                                                                 begin 
                                                                 end 
                                                     end 
                                                  else 
                                                     if ( ptw__GEN_131 )
                                                         begin 
                                                         end 
                                                      else 
                                                         if ( ptw__GEN_133 )
                                                             begin 
                                                             end 
                                                          else 
                                                             if ( ptw__GEN_138 )
                                                                 begin 
                                                                     if ( ptw__GEN_144 ) 
                                                                         ptw_count  <=2'h2;
                                                                      else 
                                                                         begin 
                                                                         end 
                                                                 end 
                                                              else 
                                                                 begin 
                                                                 end 
                                     end 
                                  else 
                                     begin  
                                         ptw_count  <= ptw_max_count ;
                                         if ( ptw__GEN_103 )
                                             begin 
                                                 if ( ptw__GEN_104 ) 
                                                     ptw_stage2  <= ptw__arb_io_out_bits_bits_stage2 ;
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin 
                                             end 
                                     end 
                         end 
                      else 
                         if ( ptw__GEN_103 )
                             begin 
                                 if ( ptw__GEN_104 )
                                     begin  
                                         ptw_count  <= ptw__GEN_108 ; 
                                         ptw_stage2  <= ptw__arb_io_out_bits_bits_stage2 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             if ( ptw__GEN_119 )
                                 begin 
                                     if ( ptw_stage2_pte_cache_hit )
                                         begin 
                                         end 
                                      else 
                                         if ( ptw_pte_cache_hit ) 
                                             ptw_count  <= ptw__GEN_126 [1:0];
                                          else 
                                             begin 
                                             end 
                                 end 
                              else 
                                 if ( ptw__GEN_131 )
                                     begin 
                                     end 
                                  else 
                                     if ( ptw__GEN_133 )
                                         begin 
                                         end 
                                      else 
                                         if ( ptw__GEN_138 )
                                             begin 
                                                 if ( ptw__GEN_144 ) 
                                                     ptw_count  <=2'h2;
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin 
                                             end 
                     if ( ptw__GEN_103 )
                         begin 
                             if ( ptw__GEN_104 )
                                 begin  
                                     ptw_aux_count  <= ptw__GEN_109 ; 
                                     ptw_aux_pte_reserved_for_future  <=10'h0; 
                                     ptw_aux_pte_ppn  <= ptw_aux_ppn ;
                                 end 
                              else 
                                 begin 
                                 end 
                         end 
                      else 
                         if ( ptw__GEN_119 )
                             begin 
                                 if ( ptw_stage2_pte_cache_hit )
                                     begin  
                                         ptw_aux_count  <= ptw__GEN_123 [1:0]; 
                                         ptw_aux_pte_reserved_for_future  <=10'h0; 
                                         ptw_aux_pte_ppn  <= ptw__GEN_124 ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                 end 
             if ( ptw_mem_resp_valid )
                 begin 
                     if ( ptw_traverse )
                         begin 
                             if ( ptw__GEN_103 )
                                 begin 
                                     if ( ptw__GEN_104 )
                                         begin  
                                             ptw_resp_ae_ptw  <=1'h0; 
                                             ptw_resp_ae_final  <=1'h0; 
                                             ptw_resp_pf  <=1'h0; 
                                             ptw_resp_gf  <= ptw__GEN_112 ; 
                                             ptw_resp_hr  <=1'h1; 
                                             ptw_resp_hw  <=1'h1; 
                                             ptw_resp_hx  <=1'h1; 
                                             ptw_stage2_final  <= ptw__GEN_106 ;
                                         end 
                                      else 
                                         begin 
                                         end 
                                 end 
                              else 
                                 if ( ptw__GEN_119 )
                                     begin 
                                     end 
                                  else 
                                     if ( ptw__GEN_131 )
                                         begin 
                                         end 
                                      else 
                                         if ( ptw__GEN_133 )
                                             begin 
                                                 if ( ptw_io_mem_s2_xcpt_ae_ld ) 
                                                     ptw_resp_ae_ptw  <=1'h1;
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin 
                                             end 
                         end 
                      else 
                         if ( ptw__GEN_156 )
                             begin 
                                 if ( ptw__GEN_103 )
                                     begin 
                                         if ( ptw__GEN_104 )
                                             begin  
                                                 ptw_resp_ae_ptw  <=1'h0; 
                                                 ptw_resp_ae_final  <=1'h0; 
                                                 ptw_resp_pf  <=1'h0; 
                                                 ptw_resp_gf  <= ptw__GEN_112 ; 
                                                 ptw_resp_hr  <=1'h1; 
                                                 ptw_resp_hw  <=1'h1; 
                                                 ptw_resp_hx  <=1'h1;
                                             end 
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     if ( ptw__GEN_119 )
                                         begin 
                                         end 
                                      else 
                                         if ( ptw__GEN_131 )
                                             begin 
                                             end 
                                          else 
                                             if ( ptw__GEN_133 )
                                                 begin 
                                                     if ( ptw_io_mem_s2_xcpt_ae_ld ) 
                                                         ptw_resp_ae_ptw  <=1'h1;
                                                      else 
                                                         begin 
                                                         end 
                                                 end 
                                              else 
                                                 begin 
                                                 end 
                                 if ( ptw_stage2 )
                                     begin 
                                         if ( ptw__GEN_103 )
                                             begin 
                                                 if ( ptw__GEN_104 ) 
                                                     ptw_stage2_final  <= ptw__GEN_106 ;
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else  
                                     ptw_stage2_final  <=1'h1;
                             end 
                          else 
                             begin  
                                 ptw_resp_ae_ptw  <= ptw__GEN_161 ; 
                                 ptw_resp_ae_final  <= ptw_ae ; 
                                 ptw_resp_pf  <= ptw__GEN_162 ; 
                                 ptw_resp_gf  <= ptw__GEN_163 ; 
                                 ptw_resp_hr  <= ptw__GEN_164 ; 
                                 ptw_resp_hw  <= ptw__GEN_165 ; 
                                 ptw_resp_hx  <= ptw__GEN_166 ;
                                 if ( ptw__GEN_103 )
                                     begin 
                                         if ( ptw__GEN_104 ) 
                                             ptw_stage2_final  <= ptw__GEN_106 ;
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                 end 
              else 
                 if ( ptw__GEN_103 )
                     begin 
                         if ( ptw__GEN_104 )
                             begin  
                                 ptw_resp_ae_ptw  <=1'h0; 
                                 ptw_resp_ae_final  <=1'h0; 
                                 ptw_resp_pf  <=1'h0; 
                                 ptw_resp_gf  <= ptw__GEN_112 ; 
                                 ptw_resp_hr  <=1'h1; 
                                 ptw_resp_hw  <=1'h1; 
                                 ptw_resp_hx  <=1'h1; 
                                 ptw_stage2_final  <= ptw__GEN_106 ;
                             end 
                          else 
                             begin 
                             end 
                     end 
                  else 
                     if ( ptw__GEN_119 )
                         begin 
                         end 
                      else 
                         if ( ptw__GEN_131 )
                             begin 
                             end 
                          else 
                             if ( ptw__GEN_133 )
                                 begin 
                                     if ( ptw_io_mem_s2_xcpt_ae_ld ) 
                                         ptw_resp_ae_ptw  <=1'h1;
                                      else 
                                         begin 
                                         end 
                                 end 
                              else 
                                 begin 
                                 end 
             if ( ptw__GEN_103 )
                 begin 
                     if ( ptw__GEN_104 )
                         begin  
                             ptw_resp_fragmented_superpage  <=1'h0; 
                             ptw_r_req_addr  <= ptw__arb_io_out_bits_bits_addr ; 
                             ptw_r_req_need_gpa  <= ptw__arb_io_out_bits_bits_need_gpa ; 
                             ptw_r_req_vstage1  <= ptw__arb_io_out_bits_bits_vstage1 ; 
                             ptw_r_req_stage2  <= ptw__arb_io_out_bits_bits_stage2 ; 
                             ptw_r_req_dest  <= ptw__arb_io_chosen ; 
                             ptw_r_hgatp_mode  <= ptw_io_dpath_hgatp_mode ; 
                             ptw_r_hgatp_asid  <= ptw_io_dpath_hgatp_asid ; 
                             ptw_r_hgatp_ppn  <= ptw_io_dpath_hgatp_ppn ;
                         end 
                      else 
                         begin 
                         end 
                 end 
              else 
                 if ( ptw__GEN_119 )
                     begin 
                         if ( ptw__GEN_121 ) 
                             ptw_gpa_pgoff  <= ptw__GEN_122 [11:0];
                          else 
                             begin 
                             end 
                     end 
                  else 
                     if ( ptw__GEN_131 )
                         begin 
                         end 
                      else 
                         if ( ptw__GEN_133 )
                             begin 
                             end 
                          else 
                             if ( ptw__GEN_138 )
                                 begin 
                                     if ( ptw_do_both_stages ) 
                                         ptw_resp_fragmented_superpage  <=1'h1;
                                      else 
                                         if ( ptw__GEN_144 ) 
                                             ptw_resp_fragmented_superpage  <=1'h1;
                                          else 
                                             begin 
                                             end 
                                 end 
                              else 
                                 begin 
                                 end  
             ptw_r_pte_reserved_for_future  <= ptw__r_pte_barrier_io_y_reserved_for_future ; 
             ptw_r_pte_ppn  <= ptw__r_pte_barrier_io_y_ppn ; 
             ptw_r_pte_reserved_for_software  <= ptw__r_pte_barrier_io_y_reserved_for_software ; 
             ptw_r_pte_d  <= ptw__r_pte_barrier_io_y_d ; 
             ptw_r_pte_a  <= ptw__r_pte_barrier_io_y_a ; 
             ptw_r_pte_g  <= ptw__r_pte_barrier_io_y_g ; 
             ptw_r_pte_u  <= ptw__r_pte_barrier_io_y_u ; 
             ptw_r_pte_x  <= ptw__r_pte_barrier_io_y_x ; 
             ptw_r_pte_w  <= ptw__r_pte_barrier_io_y_w ; 
             ptw_r_pte_r  <= ptw__r_pte_barrier_io_y_r ; 
             ptw_r_pte_v  <= ptw__r_pte_barrier_io_y_v ; 
             ptw_mem_resp_valid  <= ptw_io_mem_resp_valid ; 
             ptw_mem_resp_data  <= ptw_io_mem_resp_bits_data ;
             if ( ptw__GEN_15 )
                 begin 
                     if ( ptw__GEN_18 ) 
                         ptw_tags_0  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_19 ) 
                         ptw_tags_1  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_20 ) 
                         ptw_tags_2  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_21 ) 
                         ptw_tags_3  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_22 ) 
                         ptw_tags_4  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_23 ) 
                         ptw_tags_5  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_24 ) 
                         ptw_tags_6  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_25 ) 
                         ptw_tags_7  <= ptw_tag [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_26 ) 
                         ptw_data_0  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_27 ) 
                         ptw_data_1  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_28 ) 
                         ptw_data_2  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_29 ) 
                         ptw_data_3  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_30 ) 
                         ptw_data_4  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_31 ) 
                         ptw_data_5  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_32 ) 
                         ptw_data_6  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_33 ) 
                         ptw_data_7  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end 
             if ( ptw__GEN_40 )
                 begin 
                     if ( ptw__GEN_43 ) 
                         ptw_tags_1_0  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_44 ) 
                         ptw_tags_1_1  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_45 ) 
                         ptw_tags_1_2  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_46 ) 
                         ptw_tags_1_3  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_47 ) 
                         ptw_tags_1_4  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_48 ) 
                         ptw_tags_1_5  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_49 ) 
                         ptw_tags_1_6  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_50 ) 
                         ptw_tags_1_7  <= ptw_tag_1 [31:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_51 ) 
                         ptw_data_1_0  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_52 ) 
                         ptw_data_1_1  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_53 ) 
                         ptw_data_1_2  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_54 ) 
                         ptw_data_1_3  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_55 ) 
                         ptw_data_1_4  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_56 ) 
                         ptw_data_1_5  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_57 ) 
                         ptw_data_1_6  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                     if ( ptw__GEN_58 ) 
                         ptw_data_1_7  <= ptw_pte_ppn [19:0];
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end  
             ptw_pte_hit  <= ptw__GEN_103  ? 1'h0: ptw__GEN_119  ? ( ptw_stage2_pte_cache_hit  ? 1'h1: ptw_pte_cache_hit ):1'h0; 
             ptw_l2_refill  <= ptw_mem_resp_valid  ? ( ptw_traverse  ? 1'h0: ptw__GEN_156  ? 1'h0: ptw_success & ptw_count ==2'h2& ptw_r_req_need_gpa ==1'h0&( ptw_r_req_vstage1 ==1'h0& ptw_r_req_stage2 ==1'h0| ptw_do_both_stages & ptw_aux_count ==2'h2& ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_w & ptw_pte_d & ptw_pte_u & ptw_pte_v &( ptw_pte_r | ptw_pte_x & ptw_pte_w ==1'h0)& ptw_pte_a & ptw_pte_x & ptw_pte_u )):1'h0;
         end
  assign  ptw_io_requestor_0_resp_valid = ptw_resp_valid_0 ; 
  assign  ptw_io_requestor_0_resp_bits_ae_ptw = ptw_resp_ae_ptw ; 
  assign  ptw_io_requestor_0_resp_bits_ae_final = ptw_resp_ae_final ; 
  assign  ptw_io_requestor_0_resp_bits_pf = ptw_resp_pf ; 
  assign  ptw_io_requestor_0_resp_bits_gf = ptw_resp_gf ; 
  assign  ptw_io_requestor_0_resp_bits_hr = ptw_resp_hr ; 
  assign  ptw_io_requestor_0_resp_bits_hw = ptw_resp_hw ; 
  assign  ptw_io_requestor_0_resp_bits_hx = ptw_resp_hx ; 
  assign  ptw_io_requestor_0_resp_bits_pte_reserved_for_future = ptw_r_pte_reserved_for_future ; 
  assign  ptw_io_requestor_0_resp_bits_pte_ppn = ptw_r_pte_ppn ; 
  assign  ptw_io_requestor_0_resp_bits_pte_reserved_for_software = ptw_r_pte_reserved_for_software ; 
  assign  ptw_io_requestor_0_resp_bits_pte_d = ptw_r_pte_d ; 
  assign  ptw_io_requestor_0_resp_bits_pte_a = ptw_r_pte_a ; 
  assign  ptw_io_requestor_0_resp_bits_pte_g = ptw_r_pte_g ; 
  assign  ptw_io_requestor_0_resp_bits_pte_u = ptw_r_pte_u ; 
  assign  ptw_io_requestor_0_resp_bits_pte_x = ptw_r_pte_x ; 
  assign  ptw_io_requestor_0_resp_bits_pte_w = ptw_r_pte_w ; 
  assign  ptw_io_requestor_0_resp_bits_pte_r = ptw_r_pte_r ; 
  assign  ptw_io_requestor_0_resp_bits_pte_v = ptw_r_pte_v ; 
  assign  ptw_io_requestor_0_resp_bits_level = ptw_max_count ; 
  assign  ptw_io_requestor_0_resp_bits_fragmented_superpage =1'h0; 
  assign  ptw_io_requestor_0_resp_bits_homogeneous = ptw_homogeneous ; 
  assign  ptw_io_requestor_0_resp_bits_gpa_valid = ptw_r_req_need_gpa ; 
  assign  ptw_io_requestor_0_resp_bits_gpa_bits = ptw__GEN_101 [32:0]; 
  assign  ptw_io_requestor_0_resp_bits_gpa_is_pte = ptw_stage2_final ==1'h0; 
  assign  ptw_io_requestor_0_ptbr_mode = ptw_io_dpath_ptbr_mode ; 
  assign  ptw_io_requestor_0_ptbr_asid = ptw_io_dpath_ptbr_asid ; 
  assign  ptw_io_requestor_0_ptbr_ppn = ptw_io_dpath_ptbr_ppn ; 
  assign  ptw_io_requestor_0_hgatp_mode = ptw_io_dpath_hgatp_mode ; 
  assign  ptw_io_requestor_0_hgatp_asid = ptw_io_dpath_hgatp_asid ; 
  assign  ptw_io_requestor_0_hgatp_ppn = ptw_io_dpath_hgatp_ppn ; 
  assign  ptw_io_requestor_0_vsatp_mode = ptw_io_dpath_vsatp_mode ; 
  assign  ptw_io_requestor_0_vsatp_asid = ptw_io_dpath_vsatp_asid ; 
  assign  ptw_io_requestor_0_vsatp_ppn = ptw_io_dpath_vsatp_ppn ; 
  assign  ptw_io_requestor_0_status_debug = ptw_io_dpath_status_debug ; 
  assign  ptw_io_requestor_0_status_cease = ptw_io_dpath_status_cease ; 
  assign  ptw_io_requestor_0_status_wfi = ptw_io_dpath_status_wfi ; 
  assign  ptw_io_requestor_0_status_isa = ptw_io_dpath_status_isa ; 
  assign  ptw_io_requestor_0_status_dprv = ptw_io_dpath_status_dprv ; 
  assign  ptw_io_requestor_0_status_dv = ptw_io_dpath_status_dv ; 
  assign  ptw_io_requestor_0_status_prv = ptw_io_dpath_status_prv ; 
  assign  ptw_io_requestor_0_status_v = ptw_io_dpath_status_v ; 
  assign  ptw_io_requestor_0_status_sd = ptw_io_dpath_status_sd ; 
  assign  ptw_io_requestor_0_status_zero2 = ptw_io_dpath_status_zero2 ; 
  assign  ptw_io_requestor_0_status_mpv = ptw_io_dpath_status_mpv ; 
  assign  ptw_io_requestor_0_status_gva = ptw_io_dpath_status_gva ; 
  assign  ptw_io_requestor_0_status_mbe = ptw_io_dpath_status_mbe ; 
  assign  ptw_io_requestor_0_status_sbe = ptw_io_dpath_status_sbe ; 
  assign  ptw_io_requestor_0_status_sxl = ptw_io_dpath_status_sxl ; 
  assign  ptw_io_requestor_0_status_uxl = ptw_io_dpath_status_uxl ; 
  assign  ptw_io_requestor_0_status_sd_rv32 = ptw_io_dpath_status_sd_rv32 ; 
  assign  ptw_io_requestor_0_status_zero1 = ptw_io_dpath_status_zero1 ; 
  assign  ptw_io_requestor_0_status_tsr = ptw_io_dpath_status_tsr ; 
  assign  ptw_io_requestor_0_status_tw = ptw_io_dpath_status_tw ; 
  assign  ptw_io_requestor_0_status_tvm = ptw_io_dpath_status_tvm ; 
  assign  ptw_io_requestor_0_status_mxr = ptw_io_dpath_status_mxr ; 
  assign  ptw_io_requestor_0_status_sum = ptw_io_dpath_status_sum ; 
  assign  ptw_io_requestor_0_status_mprv = ptw_io_dpath_status_mprv ; 
  assign  ptw_io_requestor_0_status_xs = ptw_io_dpath_status_xs ; 
  assign  ptw_io_requestor_0_status_fs = ptw_io_dpath_status_fs ; 
  assign  ptw_io_requestor_0_status_mpp = ptw_io_dpath_status_mpp ; 
  assign  ptw_io_requestor_0_status_vs = ptw_io_dpath_status_vs ; 
  assign  ptw_io_requestor_0_status_spp = ptw_io_dpath_status_spp ; 
  assign  ptw_io_requestor_0_status_mpie = ptw_io_dpath_status_mpie ; 
  assign  ptw_io_requestor_0_status_ube = ptw_io_dpath_status_ube ; 
  assign  ptw_io_requestor_0_status_spie = ptw_io_dpath_status_spie ; 
  assign  ptw_io_requestor_0_status_upie = ptw_io_dpath_status_upie ; 
  assign  ptw_io_requestor_0_status_mie = ptw_io_dpath_status_mie ; 
  assign  ptw_io_requestor_0_status_hie = ptw_io_dpath_status_hie ; 
  assign  ptw_io_requestor_0_status_sie = ptw_io_dpath_status_sie ; 
  assign  ptw_io_requestor_0_status_uie = ptw_io_dpath_status_uie ; 
  assign  ptw_io_requestor_0_hstatus_zero6 = ptw_io_dpath_hstatus_zero6 ; 
  assign  ptw_io_requestor_0_hstatus_vsxl = ptw_io_dpath_hstatus_vsxl ; 
  assign  ptw_io_requestor_0_hstatus_zero5 = ptw_io_dpath_hstatus_zero5 ; 
  assign  ptw_io_requestor_0_hstatus_vtsr = ptw_io_dpath_hstatus_vtsr ; 
  assign  ptw_io_requestor_0_hstatus_vtw = ptw_io_dpath_hstatus_vtw ; 
  assign  ptw_io_requestor_0_hstatus_vtvm = ptw_io_dpath_hstatus_vtvm ; 
  assign  ptw_io_requestor_0_hstatus_zero3 = ptw_io_dpath_hstatus_zero3 ; 
  assign  ptw_io_requestor_0_hstatus_vgein = ptw_io_dpath_hstatus_vgein ; 
  assign  ptw_io_requestor_0_hstatus_zero2 = ptw_io_dpath_hstatus_zero2 ; 
  assign  ptw_io_requestor_0_hstatus_hu = ptw_io_dpath_hstatus_hu ; 
  assign  ptw_io_requestor_0_hstatus_spvp = ptw_io_dpath_hstatus_spvp ; 
  assign  ptw_io_requestor_0_hstatus_spv = ptw_io_dpath_hstatus_spv ; 
  assign  ptw_io_requestor_0_hstatus_gva = ptw_io_dpath_hstatus_gva ; 
  assign  ptw_io_requestor_0_hstatus_vsbe = ptw_io_dpath_hstatus_vsbe ; 
  assign  ptw_io_requestor_0_hstatus_zero1 = ptw_io_dpath_hstatus_zero1 ; 
  assign  ptw_io_requestor_0_gstatus_debug = ptw_io_dpath_gstatus_debug ; 
  assign  ptw_io_requestor_0_gstatus_cease = ptw_io_dpath_gstatus_cease ; 
  assign  ptw_io_requestor_0_gstatus_wfi = ptw_io_dpath_gstatus_wfi ; 
  assign  ptw_io_requestor_0_gstatus_isa = ptw_io_dpath_gstatus_isa ; 
  assign  ptw_io_requestor_0_gstatus_dprv = ptw_io_dpath_gstatus_dprv ; 
  assign  ptw_io_requestor_0_gstatus_dv = ptw_io_dpath_gstatus_dv ; 
  assign  ptw_io_requestor_0_gstatus_prv = ptw_io_dpath_gstatus_prv ; 
  assign  ptw_io_requestor_0_gstatus_v = ptw_io_dpath_gstatus_v ; 
  assign  ptw_io_requestor_0_gstatus_sd = ptw_io_dpath_gstatus_sd ; 
  assign  ptw_io_requestor_0_gstatus_zero2 = ptw_io_dpath_gstatus_zero2 ; 
  assign  ptw_io_requestor_0_gstatus_mpv = ptw_io_dpath_gstatus_mpv ; 
  assign  ptw_io_requestor_0_gstatus_gva = ptw_io_dpath_gstatus_gva ; 
  assign  ptw_io_requestor_0_gstatus_mbe = ptw_io_dpath_gstatus_mbe ; 
  assign  ptw_io_requestor_0_gstatus_sbe = ptw_io_dpath_gstatus_sbe ; 
  assign  ptw_io_requestor_0_gstatus_sxl = ptw_io_dpath_gstatus_sxl ; 
  assign  ptw_io_requestor_0_gstatus_uxl = ptw_io_dpath_gstatus_uxl ; 
  assign  ptw_io_requestor_0_gstatus_sd_rv32 = ptw_io_dpath_gstatus_sd_rv32 ; 
  assign  ptw_io_requestor_0_gstatus_zero1 = ptw_io_dpath_gstatus_zero1 ; 
  assign  ptw_io_requestor_0_gstatus_tsr = ptw_io_dpath_gstatus_tsr ; 
  assign  ptw_io_requestor_0_gstatus_tw = ptw_io_dpath_gstatus_tw ; 
  assign  ptw_io_requestor_0_gstatus_tvm = ptw_io_dpath_gstatus_tvm ; 
  assign  ptw_io_requestor_0_gstatus_mxr = ptw_io_dpath_gstatus_mxr ; 
  assign  ptw_io_requestor_0_gstatus_sum = ptw_io_dpath_gstatus_sum ; 
  assign  ptw_io_requestor_0_gstatus_mprv = ptw_io_dpath_gstatus_mprv ; 
  assign  ptw_io_requestor_0_gstatus_xs = ptw_io_dpath_gstatus_xs ; 
  assign  ptw_io_requestor_0_gstatus_fs = ptw_io_dpath_gstatus_fs ; 
  assign  ptw_io_requestor_0_gstatus_mpp = ptw_io_dpath_gstatus_mpp ; 
  assign  ptw_io_requestor_0_gstatus_vs = ptw_io_dpath_gstatus_vs ; 
  assign  ptw_io_requestor_0_gstatus_spp = ptw_io_dpath_gstatus_spp ; 
  assign  ptw_io_requestor_0_gstatus_mpie = ptw_io_dpath_gstatus_mpie ; 
  assign  ptw_io_requestor_0_gstatus_ube = ptw_io_dpath_gstatus_ube ; 
  assign  ptw_io_requestor_0_gstatus_spie = ptw_io_dpath_gstatus_spie ; 
  assign  ptw_io_requestor_0_gstatus_upie = ptw_io_dpath_gstatus_upie ; 
  assign  ptw_io_requestor_0_gstatus_mie = ptw_io_dpath_gstatus_mie ; 
  assign  ptw_io_requestor_0_gstatus_hie = ptw_io_dpath_gstatus_hie ; 
  assign  ptw_io_requestor_0_gstatus_sie = ptw_io_dpath_gstatus_sie ; 
  assign  ptw_io_requestor_0_gstatus_uie = ptw_io_dpath_gstatus_uie ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_l = ptw_io_dpath_pmp_0_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_res = ptw_io_dpath_pmp_0_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_a = ptw_io_dpath_pmp_0_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_x = ptw_io_dpath_pmp_0_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_w = ptw_io_dpath_pmp_0_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_0_cfg_r = ptw_io_dpath_pmp_0_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_0_addr = ptw_io_dpath_pmp_0_addr ; 
  assign  ptw_io_requestor_0_pmp_0_mask = ptw_io_dpath_pmp_0_mask ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_l = ptw_io_dpath_pmp_1_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_res = ptw_io_dpath_pmp_1_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_a = ptw_io_dpath_pmp_1_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_x = ptw_io_dpath_pmp_1_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_w = ptw_io_dpath_pmp_1_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_1_cfg_r = ptw_io_dpath_pmp_1_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_1_addr = ptw_io_dpath_pmp_1_addr ; 
  assign  ptw_io_requestor_0_pmp_1_mask = ptw_io_dpath_pmp_1_mask ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_l = ptw_io_dpath_pmp_2_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_res = ptw_io_dpath_pmp_2_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_a = ptw_io_dpath_pmp_2_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_x = ptw_io_dpath_pmp_2_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_w = ptw_io_dpath_pmp_2_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_2_cfg_r = ptw_io_dpath_pmp_2_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_2_addr = ptw_io_dpath_pmp_2_addr ; 
  assign  ptw_io_requestor_0_pmp_2_mask = ptw_io_dpath_pmp_2_mask ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_l = ptw_io_dpath_pmp_3_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_res = ptw_io_dpath_pmp_3_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_a = ptw_io_dpath_pmp_3_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_x = ptw_io_dpath_pmp_3_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_w = ptw_io_dpath_pmp_3_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_3_cfg_r = ptw_io_dpath_pmp_3_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_3_addr = ptw_io_dpath_pmp_3_addr ; 
  assign  ptw_io_requestor_0_pmp_3_mask = ptw_io_dpath_pmp_3_mask ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_l = ptw_io_dpath_pmp_4_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_res = ptw_io_dpath_pmp_4_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_a = ptw_io_dpath_pmp_4_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_x = ptw_io_dpath_pmp_4_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_w = ptw_io_dpath_pmp_4_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_4_cfg_r = ptw_io_dpath_pmp_4_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_4_addr = ptw_io_dpath_pmp_4_addr ; 
  assign  ptw_io_requestor_0_pmp_4_mask = ptw_io_dpath_pmp_4_mask ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_l = ptw_io_dpath_pmp_5_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_res = ptw_io_dpath_pmp_5_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_a = ptw_io_dpath_pmp_5_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_x = ptw_io_dpath_pmp_5_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_w = ptw_io_dpath_pmp_5_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_5_cfg_r = ptw_io_dpath_pmp_5_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_5_addr = ptw_io_dpath_pmp_5_addr ; 
  assign  ptw_io_requestor_0_pmp_5_mask = ptw_io_dpath_pmp_5_mask ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_l = ptw_io_dpath_pmp_6_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_res = ptw_io_dpath_pmp_6_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_a = ptw_io_dpath_pmp_6_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_x = ptw_io_dpath_pmp_6_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_w = ptw_io_dpath_pmp_6_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_6_cfg_r = ptw_io_dpath_pmp_6_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_6_addr = ptw_io_dpath_pmp_6_addr ; 
  assign  ptw_io_requestor_0_pmp_6_mask = ptw_io_dpath_pmp_6_mask ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_l = ptw_io_dpath_pmp_7_cfg_l ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_res = ptw_io_dpath_pmp_7_cfg_res ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_a = ptw_io_dpath_pmp_7_cfg_a ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_x = ptw_io_dpath_pmp_7_cfg_x ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_w = ptw_io_dpath_pmp_7_cfg_w ; 
  assign  ptw_io_requestor_0_pmp_7_cfg_r = ptw_io_dpath_pmp_7_cfg_r ; 
  assign  ptw_io_requestor_0_pmp_7_addr = ptw_io_dpath_pmp_7_addr ; 
  assign  ptw_io_requestor_0_pmp_7_mask = ptw_io_dpath_pmp_7_mask ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_0_ren = ptw_io_dpath_customCSRs_csrs_0_ren ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_0_wen = ptw_io_dpath_customCSRs_csrs_0_wen ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_0_wdata = ptw_io_dpath_customCSRs_csrs_0_wdata ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_0_value = ptw_io_dpath_customCSRs_csrs_0_value ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_1_ren = ptw_io_dpath_customCSRs_csrs_1_ren ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_1_wen = ptw_io_dpath_customCSRs_csrs_1_wen ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_1_wdata = ptw_io_dpath_customCSRs_csrs_1_wdata ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_1_value = ptw_io_dpath_customCSRs_csrs_1_value ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_2_ren = ptw_io_dpath_customCSRs_csrs_2_ren ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_2_wen = ptw_io_dpath_customCSRs_csrs_2_wen ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_2_wdata = ptw_io_dpath_customCSRs_csrs_2_wdata ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_2_value = ptw_io_dpath_customCSRs_csrs_2_value ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_3_ren = ptw_io_dpath_customCSRs_csrs_3_ren ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_3_wen = ptw_io_dpath_customCSRs_csrs_3_wen ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_3_wdata = ptw_io_dpath_customCSRs_csrs_3_wdata ; 
  assign  ptw_io_requestor_0_customCSRs_csrs_3_value = ptw_io_dpath_customCSRs_csrs_3_value ; 
  assign  ptw_io_requestor_1_resp_valid = ptw_resp_valid_1 ; 
  assign  ptw_io_requestor_1_resp_bits_ae_ptw = ptw_resp_ae_ptw ; 
  assign  ptw_io_requestor_1_resp_bits_ae_final = ptw_resp_ae_final ; 
  assign  ptw_io_requestor_1_resp_bits_pf = ptw_resp_pf ; 
  assign  ptw_io_requestor_1_resp_bits_gf = ptw_resp_gf ; 
  assign  ptw_io_requestor_1_resp_bits_hr = ptw_resp_hr ; 
  assign  ptw_io_requestor_1_resp_bits_hw = ptw_resp_hw ; 
  assign  ptw_io_requestor_1_resp_bits_hx = ptw_resp_hx ; 
  assign  ptw_io_requestor_1_resp_bits_pte_reserved_for_future = ptw_r_pte_reserved_for_future ; 
  assign  ptw_io_requestor_1_resp_bits_pte_ppn = ptw_r_pte_ppn ; 
  assign  ptw_io_requestor_1_resp_bits_pte_reserved_for_software = ptw_r_pte_reserved_for_software ; 
  assign  ptw_io_requestor_1_resp_bits_pte_d = ptw_r_pte_d ; 
  assign  ptw_io_requestor_1_resp_bits_pte_a = ptw_r_pte_a ; 
  assign  ptw_io_requestor_1_resp_bits_pte_g = ptw_r_pte_g ; 
  assign  ptw_io_requestor_1_resp_bits_pte_u = ptw_r_pte_u ; 
  assign  ptw_io_requestor_1_resp_bits_pte_x = ptw_r_pte_x ; 
  assign  ptw_io_requestor_1_resp_bits_pte_w = ptw_r_pte_w ; 
  assign  ptw_io_requestor_1_resp_bits_pte_r = ptw_r_pte_r ; 
  assign  ptw_io_requestor_1_resp_bits_pte_v = ptw_r_pte_v ; 
  assign  ptw_io_requestor_1_resp_bits_level = ptw_max_count ; 
  assign  ptw_io_requestor_1_resp_bits_fragmented_superpage =1'h0; 
  assign  ptw_io_requestor_1_resp_bits_homogeneous = ptw_homogeneous ; 
  assign  ptw_io_requestor_1_resp_bits_gpa_valid = ptw_r_req_need_gpa ; 
  assign  ptw_io_requestor_1_resp_bits_gpa_bits = ptw__GEN_102 [32:0]; 
  assign  ptw_io_requestor_1_resp_bits_gpa_is_pte = ptw_stage2_final ==1'h0; 
  assign  ptw_io_requestor_1_ptbr_mode = ptw_io_dpath_ptbr_mode ; 
  assign  ptw_io_requestor_1_ptbr_asid = ptw_io_dpath_ptbr_asid ; 
  assign  ptw_io_requestor_1_ptbr_ppn = ptw_io_dpath_ptbr_ppn ; 
  assign  ptw_io_requestor_1_hgatp_mode = ptw_io_dpath_hgatp_mode ; 
  assign  ptw_io_requestor_1_hgatp_asid = ptw_io_dpath_hgatp_asid ; 
  assign  ptw_io_requestor_1_hgatp_ppn = ptw_io_dpath_hgatp_ppn ; 
  assign  ptw_io_requestor_1_vsatp_mode = ptw_io_dpath_vsatp_mode ; 
  assign  ptw_io_requestor_1_vsatp_asid = ptw_io_dpath_vsatp_asid ; 
  assign  ptw_io_requestor_1_vsatp_ppn = ptw_io_dpath_vsatp_ppn ; 
  assign  ptw_io_requestor_1_status_debug = ptw_io_dpath_status_debug ; 
  assign  ptw_io_requestor_1_status_cease = ptw_io_dpath_status_cease ; 
  assign  ptw_io_requestor_1_status_wfi = ptw_io_dpath_status_wfi ; 
  assign  ptw_io_requestor_1_status_isa = ptw_io_dpath_status_isa ; 
  assign  ptw_io_requestor_1_status_dprv = ptw_io_dpath_status_dprv ; 
  assign  ptw_io_requestor_1_status_dv = ptw_io_dpath_status_dv ; 
  assign  ptw_io_requestor_1_status_prv = ptw_io_dpath_status_prv ; 
  assign  ptw_io_requestor_1_status_v = ptw_io_dpath_status_v ; 
  assign  ptw_io_requestor_1_status_sd = ptw_io_dpath_status_sd ; 
  assign  ptw_io_requestor_1_status_zero2 = ptw_io_dpath_status_zero2 ; 
  assign  ptw_io_requestor_1_status_mpv = ptw_io_dpath_status_mpv ; 
  assign  ptw_io_requestor_1_status_gva = ptw_io_dpath_status_gva ; 
  assign  ptw_io_requestor_1_status_mbe = ptw_io_dpath_status_mbe ; 
  assign  ptw_io_requestor_1_status_sbe = ptw_io_dpath_status_sbe ; 
  assign  ptw_io_requestor_1_status_sxl = ptw_io_dpath_status_sxl ; 
  assign  ptw_io_requestor_1_status_uxl = ptw_io_dpath_status_uxl ; 
  assign  ptw_io_requestor_1_status_sd_rv32 = ptw_io_dpath_status_sd_rv32 ; 
  assign  ptw_io_requestor_1_status_zero1 = ptw_io_dpath_status_zero1 ; 
  assign  ptw_io_requestor_1_status_tsr = ptw_io_dpath_status_tsr ; 
  assign  ptw_io_requestor_1_status_tw = ptw_io_dpath_status_tw ; 
  assign  ptw_io_requestor_1_status_tvm = ptw_io_dpath_status_tvm ; 
  assign  ptw_io_requestor_1_status_mxr = ptw_io_dpath_status_mxr ; 
  assign  ptw_io_requestor_1_status_sum = ptw_io_dpath_status_sum ; 
  assign  ptw_io_requestor_1_status_mprv = ptw_io_dpath_status_mprv ; 
  assign  ptw_io_requestor_1_status_xs = ptw_io_dpath_status_xs ; 
  assign  ptw_io_requestor_1_status_fs = ptw_io_dpath_status_fs ; 
  assign  ptw_io_requestor_1_status_mpp = ptw_io_dpath_status_mpp ; 
  assign  ptw_io_requestor_1_status_vs = ptw_io_dpath_status_vs ; 
  assign  ptw_io_requestor_1_status_spp = ptw_io_dpath_status_spp ; 
  assign  ptw_io_requestor_1_status_mpie = ptw_io_dpath_status_mpie ; 
  assign  ptw_io_requestor_1_status_ube = ptw_io_dpath_status_ube ; 
  assign  ptw_io_requestor_1_status_spie = ptw_io_dpath_status_spie ; 
  assign  ptw_io_requestor_1_status_upie = ptw_io_dpath_status_upie ; 
  assign  ptw_io_requestor_1_status_mie = ptw_io_dpath_status_mie ; 
  assign  ptw_io_requestor_1_status_hie = ptw_io_dpath_status_hie ; 
  assign  ptw_io_requestor_1_status_sie = ptw_io_dpath_status_sie ; 
  assign  ptw_io_requestor_1_status_uie = ptw_io_dpath_status_uie ; 
  assign  ptw_io_requestor_1_hstatus_zero6 = ptw_io_dpath_hstatus_zero6 ; 
  assign  ptw_io_requestor_1_hstatus_vsxl = ptw_io_dpath_hstatus_vsxl ; 
  assign  ptw_io_requestor_1_hstatus_zero5 = ptw_io_dpath_hstatus_zero5 ; 
  assign  ptw_io_requestor_1_hstatus_vtsr = ptw_io_dpath_hstatus_vtsr ; 
  assign  ptw_io_requestor_1_hstatus_vtw = ptw_io_dpath_hstatus_vtw ; 
  assign  ptw_io_requestor_1_hstatus_vtvm = ptw_io_dpath_hstatus_vtvm ; 
  assign  ptw_io_requestor_1_hstatus_zero3 = ptw_io_dpath_hstatus_zero3 ; 
  assign  ptw_io_requestor_1_hstatus_vgein = ptw_io_dpath_hstatus_vgein ; 
  assign  ptw_io_requestor_1_hstatus_zero2 = ptw_io_dpath_hstatus_zero2 ; 
  assign  ptw_io_requestor_1_hstatus_hu = ptw_io_dpath_hstatus_hu ; 
  assign  ptw_io_requestor_1_hstatus_spvp = ptw_io_dpath_hstatus_spvp ; 
  assign  ptw_io_requestor_1_hstatus_spv = ptw_io_dpath_hstatus_spv ; 
  assign  ptw_io_requestor_1_hstatus_gva = ptw_io_dpath_hstatus_gva ; 
  assign  ptw_io_requestor_1_hstatus_vsbe = ptw_io_dpath_hstatus_vsbe ; 
  assign  ptw_io_requestor_1_hstatus_zero1 = ptw_io_dpath_hstatus_zero1 ; 
  assign  ptw_io_requestor_1_gstatus_debug = ptw_io_dpath_gstatus_debug ; 
  assign  ptw_io_requestor_1_gstatus_cease = ptw_io_dpath_gstatus_cease ; 
  assign  ptw_io_requestor_1_gstatus_wfi = ptw_io_dpath_gstatus_wfi ; 
  assign  ptw_io_requestor_1_gstatus_isa = ptw_io_dpath_gstatus_isa ; 
  assign  ptw_io_requestor_1_gstatus_dprv = ptw_io_dpath_gstatus_dprv ; 
  assign  ptw_io_requestor_1_gstatus_dv = ptw_io_dpath_gstatus_dv ; 
  assign  ptw_io_requestor_1_gstatus_prv = ptw_io_dpath_gstatus_prv ; 
  assign  ptw_io_requestor_1_gstatus_v = ptw_io_dpath_gstatus_v ; 
  assign  ptw_io_requestor_1_gstatus_sd = ptw_io_dpath_gstatus_sd ; 
  assign  ptw_io_requestor_1_gstatus_zero2 = ptw_io_dpath_gstatus_zero2 ; 
  assign  ptw_io_requestor_1_gstatus_mpv = ptw_io_dpath_gstatus_mpv ; 
  assign  ptw_io_requestor_1_gstatus_gva = ptw_io_dpath_gstatus_gva ; 
  assign  ptw_io_requestor_1_gstatus_mbe = ptw_io_dpath_gstatus_mbe ; 
  assign  ptw_io_requestor_1_gstatus_sbe = ptw_io_dpath_gstatus_sbe ; 
  assign  ptw_io_requestor_1_gstatus_sxl = ptw_io_dpath_gstatus_sxl ; 
  assign  ptw_io_requestor_1_gstatus_uxl = ptw_io_dpath_gstatus_uxl ; 
  assign  ptw_io_requestor_1_gstatus_sd_rv32 = ptw_io_dpath_gstatus_sd_rv32 ; 
  assign  ptw_io_requestor_1_gstatus_zero1 = ptw_io_dpath_gstatus_zero1 ; 
  assign  ptw_io_requestor_1_gstatus_tsr = ptw_io_dpath_gstatus_tsr ; 
  assign  ptw_io_requestor_1_gstatus_tw = ptw_io_dpath_gstatus_tw ; 
  assign  ptw_io_requestor_1_gstatus_tvm = ptw_io_dpath_gstatus_tvm ; 
  assign  ptw_io_requestor_1_gstatus_mxr = ptw_io_dpath_gstatus_mxr ; 
  assign  ptw_io_requestor_1_gstatus_sum = ptw_io_dpath_gstatus_sum ; 
  assign  ptw_io_requestor_1_gstatus_mprv = ptw_io_dpath_gstatus_mprv ; 
  assign  ptw_io_requestor_1_gstatus_xs = ptw_io_dpath_gstatus_xs ; 
  assign  ptw_io_requestor_1_gstatus_fs = ptw_io_dpath_gstatus_fs ; 
  assign  ptw_io_requestor_1_gstatus_mpp = ptw_io_dpath_gstatus_mpp ; 
  assign  ptw_io_requestor_1_gstatus_vs = ptw_io_dpath_gstatus_vs ; 
  assign  ptw_io_requestor_1_gstatus_spp = ptw_io_dpath_gstatus_spp ; 
  assign  ptw_io_requestor_1_gstatus_mpie = ptw_io_dpath_gstatus_mpie ; 
  assign  ptw_io_requestor_1_gstatus_ube = ptw_io_dpath_gstatus_ube ; 
  assign  ptw_io_requestor_1_gstatus_spie = ptw_io_dpath_gstatus_spie ; 
  assign  ptw_io_requestor_1_gstatus_upie = ptw_io_dpath_gstatus_upie ; 
  assign  ptw_io_requestor_1_gstatus_mie = ptw_io_dpath_gstatus_mie ; 
  assign  ptw_io_requestor_1_gstatus_hie = ptw_io_dpath_gstatus_hie ; 
  assign  ptw_io_requestor_1_gstatus_sie = ptw_io_dpath_gstatus_sie ; 
  assign  ptw_io_requestor_1_gstatus_uie = ptw_io_dpath_gstatus_uie ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_l = ptw_io_dpath_pmp_0_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_res = ptw_io_dpath_pmp_0_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_a = ptw_io_dpath_pmp_0_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_x = ptw_io_dpath_pmp_0_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_w = ptw_io_dpath_pmp_0_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_0_cfg_r = ptw_io_dpath_pmp_0_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_0_addr = ptw_io_dpath_pmp_0_addr ; 
  assign  ptw_io_requestor_1_pmp_0_mask = ptw_io_dpath_pmp_0_mask ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_l = ptw_io_dpath_pmp_1_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_res = ptw_io_dpath_pmp_1_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_a = ptw_io_dpath_pmp_1_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_x = ptw_io_dpath_pmp_1_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_w = ptw_io_dpath_pmp_1_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_1_cfg_r = ptw_io_dpath_pmp_1_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_1_addr = ptw_io_dpath_pmp_1_addr ; 
  assign  ptw_io_requestor_1_pmp_1_mask = ptw_io_dpath_pmp_1_mask ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_l = ptw_io_dpath_pmp_2_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_res = ptw_io_dpath_pmp_2_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_a = ptw_io_dpath_pmp_2_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_x = ptw_io_dpath_pmp_2_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_w = ptw_io_dpath_pmp_2_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_2_cfg_r = ptw_io_dpath_pmp_2_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_2_addr = ptw_io_dpath_pmp_2_addr ; 
  assign  ptw_io_requestor_1_pmp_2_mask = ptw_io_dpath_pmp_2_mask ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_l = ptw_io_dpath_pmp_3_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_res = ptw_io_dpath_pmp_3_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_a = ptw_io_dpath_pmp_3_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_x = ptw_io_dpath_pmp_3_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_w = ptw_io_dpath_pmp_3_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_3_cfg_r = ptw_io_dpath_pmp_3_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_3_addr = ptw_io_dpath_pmp_3_addr ; 
  assign  ptw_io_requestor_1_pmp_3_mask = ptw_io_dpath_pmp_3_mask ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_l = ptw_io_dpath_pmp_4_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_res = ptw_io_dpath_pmp_4_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_a = ptw_io_dpath_pmp_4_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_x = ptw_io_dpath_pmp_4_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_w = ptw_io_dpath_pmp_4_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_4_cfg_r = ptw_io_dpath_pmp_4_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_4_addr = ptw_io_dpath_pmp_4_addr ; 
  assign  ptw_io_requestor_1_pmp_4_mask = ptw_io_dpath_pmp_4_mask ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_l = ptw_io_dpath_pmp_5_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_res = ptw_io_dpath_pmp_5_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_a = ptw_io_dpath_pmp_5_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_x = ptw_io_dpath_pmp_5_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_w = ptw_io_dpath_pmp_5_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_5_cfg_r = ptw_io_dpath_pmp_5_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_5_addr = ptw_io_dpath_pmp_5_addr ; 
  assign  ptw_io_requestor_1_pmp_5_mask = ptw_io_dpath_pmp_5_mask ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_l = ptw_io_dpath_pmp_6_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_res = ptw_io_dpath_pmp_6_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_a = ptw_io_dpath_pmp_6_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_x = ptw_io_dpath_pmp_6_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_w = ptw_io_dpath_pmp_6_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_6_cfg_r = ptw_io_dpath_pmp_6_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_6_addr = ptw_io_dpath_pmp_6_addr ; 
  assign  ptw_io_requestor_1_pmp_6_mask = ptw_io_dpath_pmp_6_mask ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_l = ptw_io_dpath_pmp_7_cfg_l ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_res = ptw_io_dpath_pmp_7_cfg_res ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_a = ptw_io_dpath_pmp_7_cfg_a ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_x = ptw_io_dpath_pmp_7_cfg_x ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_w = ptw_io_dpath_pmp_7_cfg_w ; 
  assign  ptw_io_requestor_1_pmp_7_cfg_r = ptw_io_dpath_pmp_7_cfg_r ; 
  assign  ptw_io_requestor_1_pmp_7_addr = ptw_io_dpath_pmp_7_addr ; 
  assign  ptw_io_requestor_1_pmp_7_mask = ptw_io_dpath_pmp_7_mask ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_0_ren = ptw_io_dpath_customCSRs_csrs_0_ren ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_0_wen = ptw_io_dpath_customCSRs_csrs_0_wen ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_0_wdata = ptw_io_dpath_customCSRs_csrs_0_wdata ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_0_value = ptw_io_dpath_customCSRs_csrs_0_value ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_1_ren = ptw_io_dpath_customCSRs_csrs_1_ren ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_1_wen = ptw_io_dpath_customCSRs_csrs_1_wen ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_1_wdata = ptw_io_dpath_customCSRs_csrs_1_wdata ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_1_value = ptw_io_dpath_customCSRs_csrs_1_value ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_2_ren = ptw_io_dpath_customCSRs_csrs_2_ren ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_2_wen = ptw_io_dpath_customCSRs_csrs_2_wen ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_2_wdata = ptw_io_dpath_customCSRs_csrs_2_wdata ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_2_value = ptw_io_dpath_customCSRs_csrs_2_value ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_3_ren = ptw_io_dpath_customCSRs_csrs_3_ren ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_3_wen = ptw_io_dpath_customCSRs_csrs_3_wen ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_3_wdata = ptw_io_dpath_customCSRs_csrs_3_wdata ; 
  assign  ptw_io_requestor_1_customCSRs_csrs_3_value = ptw_io_dpath_customCSRs_csrs_3_value ; 
  assign  ptw_io_mem_req_valid = ptw_state ==3'h1| ptw_state ==3'h3; 
  assign  ptw_io_mem_req_bits_addr =34'h0; 
  assign  ptw_io_mem_req_bits_tag =6'h0; 
  assign  ptw_io_mem_req_bits_cmd =5'h0; 
  assign  ptw_io_mem_req_bits_size =2'h3; 
  assign  ptw_io_mem_req_bits_signed =1'h0; 
  assign  ptw_io_mem_req_bits_dprv =2'h1; 
  assign  ptw_io_mem_req_bits_dv = ptw_do_both_stages & ptw_stage2 ==1'h0; 
  assign  ptw_io_mem_req_bits_phys =1'h1; 
  assign  ptw_io_mem_req_bits_no_alloc =1'h0; 
  assign  ptw_io_mem_req_bits_no_xcpt =1'h0; 
  assign  ptw_io_mem_req_bits_data =64'h0; 
  assign  ptw_io_mem_req_bits_mask =8'h0; 
  assign  ptw_io_mem_s1_kill = ptw_state !=3'h2|1'h0| ptw_resp_gf ; 
  assign  ptw_io_mem_s1_data_data =64'h0; 
  assign  ptw_io_mem_s1_data_mask =8'h0; 
  assign  ptw_io_mem_s2_kill =1'h0; 
  assign  ptw_io_mem_keep_clock_enabled =1'h0; 
  assign  ptw_io_dpath_perf_l2miss =1'h0; 
  assign  ptw_io_dpath_perf_l2hit = ptw__io_dpath_perf_l2hit_output ; 
  assign  ptw_io_dpath_perf_pte_miss = ptw__io_dpath_perf_pte_miss_output ; 
  assign  ptw_io_dpath_perf_pte_hit = ptw__io_dpath_perf_pte_hit_output ; 
  assign  ptw_io_dpath_customCSRs_csrs_0_stall = ptw_io_requestor_1_customCSRs_csrs_0_stall ; 
  assign  ptw_io_dpath_customCSRs_csrs_0_set = ptw_io_requestor_1_customCSRs_csrs_0_set ; 
  assign  ptw_io_dpath_customCSRs_csrs_0_sdata = ptw_io_requestor_1_customCSRs_csrs_0_sdata ; 
  assign  ptw_io_dpath_customCSRs_csrs_1_stall = ptw_io_requestor_1_customCSRs_csrs_1_stall ; 
  assign  ptw_io_dpath_customCSRs_csrs_1_set = ptw_io_requestor_1_customCSRs_csrs_1_set ; 
  assign  ptw_io_dpath_customCSRs_csrs_1_sdata = ptw_io_requestor_1_customCSRs_csrs_1_sdata ; 
  assign  ptw_io_dpath_customCSRs_csrs_2_stall = ptw_io_requestor_1_customCSRs_csrs_2_stall ; 
  assign  ptw_io_dpath_customCSRs_csrs_2_set = ptw_io_requestor_1_customCSRs_csrs_2_set ; 
  assign  ptw_io_dpath_customCSRs_csrs_2_sdata = ptw_io_requestor_1_customCSRs_csrs_2_sdata ; 
  assign  ptw_io_dpath_customCSRs_csrs_3_stall = ptw_io_requestor_1_customCSRs_csrs_3_stall ; 
  assign  ptw_io_dpath_customCSRs_csrs_3_set = ptw_io_requestor_1_customCSRs_csrs_3_set ; 
  assign  ptw_io_dpath_customCSRs_csrs_3_sdata = ptw_io_requestor_1_customCSRs_csrs_3_sdata ; 
  assign  ptw_io_dpath_clock_enabled =1'h0;
    assign ptw_clock = clock;
    assign ptw_reset = reset;
    assign _ptw_io_requestor_0_req_ready = ptw_io_requestor_0_req_ready;
    assign ptw_io_requestor_0_req_valid = _dcache_io_ptw_req_valid;
    assign ptw_io_requestor_0_req_bits_valid = _dcache_io_ptw_req_bits_valid;
    assign ptw_io_requestor_0_req_bits_bits_addr = _dcache_io_ptw_req_bits_bits_addr;
    assign ptw_io_requestor_0_req_bits_bits_need_gpa = _dcache_io_ptw_req_bits_bits_need_gpa;
    assign ptw_io_requestor_0_req_bits_bits_vstage1 = _dcache_io_ptw_req_bits_bits_vstage1;
    assign ptw_io_requestor_0_req_bits_bits_stage2 = _dcache_io_ptw_req_bits_bits_stage2;
    assign _ptw_io_requestor_0_resp_valid = ptw_io_requestor_0_resp_valid;
    assign _ptw_io_requestor_0_resp_bits_ae_ptw = ptw_io_requestor_0_resp_bits_ae_ptw;
    assign _ptw_io_requestor_0_resp_bits_ae_final = ptw_io_requestor_0_resp_bits_ae_final;
    assign _ptw_io_requestor_0_resp_bits_pf = ptw_io_requestor_0_resp_bits_pf;
    assign _ptw_io_requestor_0_resp_bits_gf = ptw_io_requestor_0_resp_bits_gf;
    assign _ptw_io_requestor_0_resp_bits_hr = ptw_io_requestor_0_resp_bits_hr;
    assign _ptw_io_requestor_0_resp_bits_hw = ptw_io_requestor_0_resp_bits_hw;
    assign _ptw_io_requestor_0_resp_bits_hx = ptw_io_requestor_0_resp_bits_hx;
    assign _ptw_io_requestor_0_resp_bits_pte_reserved_for_future = ptw_io_requestor_0_resp_bits_pte_reserved_for_future;
    assign _ptw_io_requestor_0_resp_bits_pte_ppn = ptw_io_requestor_0_resp_bits_pte_ppn;
    assign _ptw_io_requestor_0_resp_bits_pte_reserved_for_software = ptw_io_requestor_0_resp_bits_pte_reserved_for_software;
    assign _ptw_io_requestor_0_resp_bits_pte_d = ptw_io_requestor_0_resp_bits_pte_d;
    assign _ptw_io_requestor_0_resp_bits_pte_a = ptw_io_requestor_0_resp_bits_pte_a;
    assign _ptw_io_requestor_0_resp_bits_pte_g = ptw_io_requestor_0_resp_bits_pte_g;
    assign _ptw_io_requestor_0_resp_bits_pte_u = ptw_io_requestor_0_resp_bits_pte_u;
    assign _ptw_io_requestor_0_resp_bits_pte_x = ptw_io_requestor_0_resp_bits_pte_x;
    assign _ptw_io_requestor_0_resp_bits_pte_w = ptw_io_requestor_0_resp_bits_pte_w;
    assign _ptw_io_requestor_0_resp_bits_pte_r = ptw_io_requestor_0_resp_bits_pte_r;
    assign _ptw_io_requestor_0_resp_bits_pte_v = ptw_io_requestor_0_resp_bits_pte_v;
    assign _ptw_io_requestor_0_resp_bits_level = ptw_io_requestor_0_resp_bits_level;
    assign _ptw_io_requestor_0_resp_bits_fragmented_superpage = ptw_io_requestor_0_resp_bits_fragmented_superpage;
    assign _ptw_io_requestor_0_resp_bits_homogeneous = ptw_io_requestor_0_resp_bits_homogeneous;
    assign _ptw_io_requestor_0_resp_bits_gpa_valid = ptw_io_requestor_0_resp_bits_gpa_valid;
    assign _ptw_io_requestor_0_resp_bits_gpa_bits = ptw_io_requestor_0_resp_bits_gpa_bits;
    assign _ptw_io_requestor_0_resp_bits_gpa_is_pte = ptw_io_requestor_0_resp_bits_gpa_is_pte;
    assign _ptw_io_requestor_0_ptbr_mode = ptw_io_requestor_0_ptbr_mode;
    assign _ptw_io_requestor_0_ptbr_asid = ptw_io_requestor_0_ptbr_asid;
    assign _ptw_io_requestor_0_ptbr_ppn = ptw_io_requestor_0_ptbr_ppn;
    assign _ptw_io_requestor_0_hgatp_mode = ptw_io_requestor_0_hgatp_mode;
    assign _ptw_io_requestor_0_hgatp_asid = ptw_io_requestor_0_hgatp_asid;
    assign _ptw_io_requestor_0_hgatp_ppn = ptw_io_requestor_0_hgatp_ppn;
    assign _ptw_io_requestor_0_vsatp_mode = ptw_io_requestor_0_vsatp_mode;
    assign _ptw_io_requestor_0_vsatp_asid = ptw_io_requestor_0_vsatp_asid;
    assign _ptw_io_requestor_0_vsatp_ppn = ptw_io_requestor_0_vsatp_ppn;
    assign _ptw_io_requestor_0_status_debug = ptw_io_requestor_0_status_debug;
    assign _ptw_io_requestor_0_status_cease = ptw_io_requestor_0_status_cease;
    assign _ptw_io_requestor_0_status_wfi = ptw_io_requestor_0_status_wfi;
    assign _ptw_io_requestor_0_status_isa = ptw_io_requestor_0_status_isa;
    assign _ptw_io_requestor_0_status_dprv = ptw_io_requestor_0_status_dprv;
    assign _ptw_io_requestor_0_status_dv = ptw_io_requestor_0_status_dv;
    assign _ptw_io_requestor_0_status_prv = ptw_io_requestor_0_status_prv;
    assign _ptw_io_requestor_0_status_v = ptw_io_requestor_0_status_v;
    assign _ptw_io_requestor_0_status_sd = ptw_io_requestor_0_status_sd;
    assign _ptw_io_requestor_0_status_zero2 = ptw_io_requestor_0_status_zero2;
    assign _ptw_io_requestor_0_status_mpv = ptw_io_requestor_0_status_mpv;
    assign _ptw_io_requestor_0_status_gva = ptw_io_requestor_0_status_gva;
    assign _ptw_io_requestor_0_status_mbe = ptw_io_requestor_0_status_mbe;
    assign _ptw_io_requestor_0_status_sbe = ptw_io_requestor_0_status_sbe;
    assign _ptw_io_requestor_0_status_sxl = ptw_io_requestor_0_status_sxl;
    assign _ptw_io_requestor_0_status_uxl = ptw_io_requestor_0_status_uxl;
    assign _ptw_io_requestor_0_status_sd_rv32 = ptw_io_requestor_0_status_sd_rv32;
    assign _ptw_io_requestor_0_status_zero1 = ptw_io_requestor_0_status_zero1;
    assign _ptw_io_requestor_0_status_tsr = ptw_io_requestor_0_status_tsr;
    assign _ptw_io_requestor_0_status_tw = ptw_io_requestor_0_status_tw;
    assign _ptw_io_requestor_0_status_tvm = ptw_io_requestor_0_status_tvm;
    assign _ptw_io_requestor_0_status_mxr = ptw_io_requestor_0_status_mxr;
    assign _ptw_io_requestor_0_status_sum = ptw_io_requestor_0_status_sum;
    assign _ptw_io_requestor_0_status_mprv = ptw_io_requestor_0_status_mprv;
    assign _ptw_io_requestor_0_status_xs = ptw_io_requestor_0_status_xs;
    assign _ptw_io_requestor_0_status_fs = ptw_io_requestor_0_status_fs;
    assign _ptw_io_requestor_0_status_mpp = ptw_io_requestor_0_status_mpp;
    assign _ptw_io_requestor_0_status_vs = ptw_io_requestor_0_status_vs;
    assign _ptw_io_requestor_0_status_spp = ptw_io_requestor_0_status_spp;
    assign _ptw_io_requestor_0_status_mpie = ptw_io_requestor_0_status_mpie;
    assign _ptw_io_requestor_0_status_ube = ptw_io_requestor_0_status_ube;
    assign _ptw_io_requestor_0_status_spie = ptw_io_requestor_0_status_spie;
    assign _ptw_io_requestor_0_status_upie = ptw_io_requestor_0_status_upie;
    assign _ptw_io_requestor_0_status_mie = ptw_io_requestor_0_status_mie;
    assign _ptw_io_requestor_0_status_hie = ptw_io_requestor_0_status_hie;
    assign _ptw_io_requestor_0_status_sie = ptw_io_requestor_0_status_sie;
    assign _ptw_io_requestor_0_status_uie = ptw_io_requestor_0_status_uie;
    assign _ptw_io_requestor_0_hstatus_zero6 = ptw_io_requestor_0_hstatus_zero6;
    assign _ptw_io_requestor_0_hstatus_vsxl = ptw_io_requestor_0_hstatus_vsxl;
    assign _ptw_io_requestor_0_hstatus_zero5 = ptw_io_requestor_0_hstatus_zero5;
    assign _ptw_io_requestor_0_hstatus_vtsr = ptw_io_requestor_0_hstatus_vtsr;
    assign _ptw_io_requestor_0_hstatus_vtw = ptw_io_requestor_0_hstatus_vtw;
    assign _ptw_io_requestor_0_hstatus_vtvm = ptw_io_requestor_0_hstatus_vtvm;
    assign _ptw_io_requestor_0_hstatus_zero3 = ptw_io_requestor_0_hstatus_zero3;
    assign _ptw_io_requestor_0_hstatus_vgein = ptw_io_requestor_0_hstatus_vgein;
    assign _ptw_io_requestor_0_hstatus_zero2 = ptw_io_requestor_0_hstatus_zero2;
    assign _ptw_io_requestor_0_hstatus_hu = ptw_io_requestor_0_hstatus_hu;
    assign _ptw_io_requestor_0_hstatus_spvp = ptw_io_requestor_0_hstatus_spvp;
    assign _ptw_io_requestor_0_hstatus_spv = ptw_io_requestor_0_hstatus_spv;
    assign _ptw_io_requestor_0_hstatus_gva = ptw_io_requestor_0_hstatus_gva;
    assign _ptw_io_requestor_0_hstatus_vsbe = ptw_io_requestor_0_hstatus_vsbe;
    assign _ptw_io_requestor_0_hstatus_zero1 = ptw_io_requestor_0_hstatus_zero1;
    assign _ptw_io_requestor_0_gstatus_debug = ptw_io_requestor_0_gstatus_debug;
    assign _ptw_io_requestor_0_gstatus_cease = ptw_io_requestor_0_gstatus_cease;
    assign _ptw_io_requestor_0_gstatus_wfi = ptw_io_requestor_0_gstatus_wfi;
    assign _ptw_io_requestor_0_gstatus_isa = ptw_io_requestor_0_gstatus_isa;
    assign _ptw_io_requestor_0_gstatus_dprv = ptw_io_requestor_0_gstatus_dprv;
    assign _ptw_io_requestor_0_gstatus_dv = ptw_io_requestor_0_gstatus_dv;
    assign _ptw_io_requestor_0_gstatus_prv = ptw_io_requestor_0_gstatus_prv;
    assign _ptw_io_requestor_0_gstatus_v = ptw_io_requestor_0_gstatus_v;
    assign _ptw_io_requestor_0_gstatus_sd = ptw_io_requestor_0_gstatus_sd;
    assign _ptw_io_requestor_0_gstatus_zero2 = ptw_io_requestor_0_gstatus_zero2;
    assign _ptw_io_requestor_0_gstatus_mpv = ptw_io_requestor_0_gstatus_mpv;
    assign _ptw_io_requestor_0_gstatus_gva = ptw_io_requestor_0_gstatus_gva;
    assign _ptw_io_requestor_0_gstatus_mbe = ptw_io_requestor_0_gstatus_mbe;
    assign _ptw_io_requestor_0_gstatus_sbe = ptw_io_requestor_0_gstatus_sbe;
    assign _ptw_io_requestor_0_gstatus_sxl = ptw_io_requestor_0_gstatus_sxl;
    assign _ptw_io_requestor_0_gstatus_uxl = ptw_io_requestor_0_gstatus_uxl;
    assign _ptw_io_requestor_0_gstatus_sd_rv32 = ptw_io_requestor_0_gstatus_sd_rv32;
    assign _ptw_io_requestor_0_gstatus_zero1 = ptw_io_requestor_0_gstatus_zero1;
    assign _ptw_io_requestor_0_gstatus_tsr = ptw_io_requestor_0_gstatus_tsr;
    assign _ptw_io_requestor_0_gstatus_tw = ptw_io_requestor_0_gstatus_tw;
    assign _ptw_io_requestor_0_gstatus_tvm = ptw_io_requestor_0_gstatus_tvm;
    assign _ptw_io_requestor_0_gstatus_mxr = ptw_io_requestor_0_gstatus_mxr;
    assign _ptw_io_requestor_0_gstatus_sum = ptw_io_requestor_0_gstatus_sum;
    assign _ptw_io_requestor_0_gstatus_mprv = ptw_io_requestor_0_gstatus_mprv;
    assign _ptw_io_requestor_0_gstatus_xs = ptw_io_requestor_0_gstatus_xs;
    assign _ptw_io_requestor_0_gstatus_fs = ptw_io_requestor_0_gstatus_fs;
    assign _ptw_io_requestor_0_gstatus_mpp = ptw_io_requestor_0_gstatus_mpp;
    assign _ptw_io_requestor_0_gstatus_vs = ptw_io_requestor_0_gstatus_vs;
    assign _ptw_io_requestor_0_gstatus_spp = ptw_io_requestor_0_gstatus_spp;
    assign _ptw_io_requestor_0_gstatus_mpie = ptw_io_requestor_0_gstatus_mpie;
    assign _ptw_io_requestor_0_gstatus_ube = ptw_io_requestor_0_gstatus_ube;
    assign _ptw_io_requestor_0_gstatus_spie = ptw_io_requestor_0_gstatus_spie;
    assign _ptw_io_requestor_0_gstatus_upie = ptw_io_requestor_0_gstatus_upie;
    assign _ptw_io_requestor_0_gstatus_mie = ptw_io_requestor_0_gstatus_mie;
    assign _ptw_io_requestor_0_gstatus_hie = ptw_io_requestor_0_gstatus_hie;
    assign _ptw_io_requestor_0_gstatus_sie = ptw_io_requestor_0_gstatus_sie;
    assign _ptw_io_requestor_0_gstatus_uie = ptw_io_requestor_0_gstatus_uie;
    assign _ptw_io_requestor_0_pmp_0_cfg_l = ptw_io_requestor_0_pmp_0_cfg_l;
    assign _ptw_io_requestor_0_pmp_0_cfg_res = ptw_io_requestor_0_pmp_0_cfg_res;
    assign _ptw_io_requestor_0_pmp_0_cfg_a = ptw_io_requestor_0_pmp_0_cfg_a;
    assign _ptw_io_requestor_0_pmp_0_cfg_x = ptw_io_requestor_0_pmp_0_cfg_x;
    assign _ptw_io_requestor_0_pmp_0_cfg_w = ptw_io_requestor_0_pmp_0_cfg_w;
    assign _ptw_io_requestor_0_pmp_0_cfg_r = ptw_io_requestor_0_pmp_0_cfg_r;
    assign _ptw_io_requestor_0_pmp_0_addr = ptw_io_requestor_0_pmp_0_addr;
    assign _ptw_io_requestor_0_pmp_0_mask = ptw_io_requestor_0_pmp_0_mask;
    assign _ptw_io_requestor_0_pmp_1_cfg_l = ptw_io_requestor_0_pmp_1_cfg_l;
    assign _ptw_io_requestor_0_pmp_1_cfg_res = ptw_io_requestor_0_pmp_1_cfg_res;
    assign _ptw_io_requestor_0_pmp_1_cfg_a = ptw_io_requestor_0_pmp_1_cfg_a;
    assign _ptw_io_requestor_0_pmp_1_cfg_x = ptw_io_requestor_0_pmp_1_cfg_x;
    assign _ptw_io_requestor_0_pmp_1_cfg_w = ptw_io_requestor_0_pmp_1_cfg_w;
    assign _ptw_io_requestor_0_pmp_1_cfg_r = ptw_io_requestor_0_pmp_1_cfg_r;
    assign _ptw_io_requestor_0_pmp_1_addr = ptw_io_requestor_0_pmp_1_addr;
    assign _ptw_io_requestor_0_pmp_1_mask = ptw_io_requestor_0_pmp_1_mask;
    assign _ptw_io_requestor_0_pmp_2_cfg_l = ptw_io_requestor_0_pmp_2_cfg_l;
    assign _ptw_io_requestor_0_pmp_2_cfg_res = ptw_io_requestor_0_pmp_2_cfg_res;
    assign _ptw_io_requestor_0_pmp_2_cfg_a = ptw_io_requestor_0_pmp_2_cfg_a;
    assign _ptw_io_requestor_0_pmp_2_cfg_x = ptw_io_requestor_0_pmp_2_cfg_x;
    assign _ptw_io_requestor_0_pmp_2_cfg_w = ptw_io_requestor_0_pmp_2_cfg_w;
    assign _ptw_io_requestor_0_pmp_2_cfg_r = ptw_io_requestor_0_pmp_2_cfg_r;
    assign _ptw_io_requestor_0_pmp_2_addr = ptw_io_requestor_0_pmp_2_addr;
    assign _ptw_io_requestor_0_pmp_2_mask = ptw_io_requestor_0_pmp_2_mask;
    assign _ptw_io_requestor_0_pmp_3_cfg_l = ptw_io_requestor_0_pmp_3_cfg_l;
    assign _ptw_io_requestor_0_pmp_3_cfg_res = ptw_io_requestor_0_pmp_3_cfg_res;
    assign _ptw_io_requestor_0_pmp_3_cfg_a = ptw_io_requestor_0_pmp_3_cfg_a;
    assign _ptw_io_requestor_0_pmp_3_cfg_x = ptw_io_requestor_0_pmp_3_cfg_x;
    assign _ptw_io_requestor_0_pmp_3_cfg_w = ptw_io_requestor_0_pmp_3_cfg_w;
    assign _ptw_io_requestor_0_pmp_3_cfg_r = ptw_io_requestor_0_pmp_3_cfg_r;
    assign _ptw_io_requestor_0_pmp_3_addr = ptw_io_requestor_0_pmp_3_addr;
    assign _ptw_io_requestor_0_pmp_3_mask = ptw_io_requestor_0_pmp_3_mask;
    assign _ptw_io_requestor_0_pmp_4_cfg_l = ptw_io_requestor_0_pmp_4_cfg_l;
    assign _ptw_io_requestor_0_pmp_4_cfg_res = ptw_io_requestor_0_pmp_4_cfg_res;
    assign _ptw_io_requestor_0_pmp_4_cfg_a = ptw_io_requestor_0_pmp_4_cfg_a;
    assign _ptw_io_requestor_0_pmp_4_cfg_x = ptw_io_requestor_0_pmp_4_cfg_x;
    assign _ptw_io_requestor_0_pmp_4_cfg_w = ptw_io_requestor_0_pmp_4_cfg_w;
    assign _ptw_io_requestor_0_pmp_4_cfg_r = ptw_io_requestor_0_pmp_4_cfg_r;
    assign _ptw_io_requestor_0_pmp_4_addr = ptw_io_requestor_0_pmp_4_addr;
    assign _ptw_io_requestor_0_pmp_4_mask = ptw_io_requestor_0_pmp_4_mask;
    assign _ptw_io_requestor_0_pmp_5_cfg_l = ptw_io_requestor_0_pmp_5_cfg_l;
    assign _ptw_io_requestor_0_pmp_5_cfg_res = ptw_io_requestor_0_pmp_5_cfg_res;
    assign _ptw_io_requestor_0_pmp_5_cfg_a = ptw_io_requestor_0_pmp_5_cfg_a;
    assign _ptw_io_requestor_0_pmp_5_cfg_x = ptw_io_requestor_0_pmp_5_cfg_x;
    assign _ptw_io_requestor_0_pmp_5_cfg_w = ptw_io_requestor_0_pmp_5_cfg_w;
    assign _ptw_io_requestor_0_pmp_5_cfg_r = ptw_io_requestor_0_pmp_5_cfg_r;
    assign _ptw_io_requestor_0_pmp_5_addr = ptw_io_requestor_0_pmp_5_addr;
    assign _ptw_io_requestor_0_pmp_5_mask = ptw_io_requestor_0_pmp_5_mask;
    assign _ptw_io_requestor_0_pmp_6_cfg_l = ptw_io_requestor_0_pmp_6_cfg_l;
    assign _ptw_io_requestor_0_pmp_6_cfg_res = ptw_io_requestor_0_pmp_6_cfg_res;
    assign _ptw_io_requestor_0_pmp_6_cfg_a = ptw_io_requestor_0_pmp_6_cfg_a;
    assign _ptw_io_requestor_0_pmp_6_cfg_x = ptw_io_requestor_0_pmp_6_cfg_x;
    assign _ptw_io_requestor_0_pmp_6_cfg_w = ptw_io_requestor_0_pmp_6_cfg_w;
    assign _ptw_io_requestor_0_pmp_6_cfg_r = ptw_io_requestor_0_pmp_6_cfg_r;
    assign _ptw_io_requestor_0_pmp_6_addr = ptw_io_requestor_0_pmp_6_addr;
    assign _ptw_io_requestor_0_pmp_6_mask = ptw_io_requestor_0_pmp_6_mask;
    assign _ptw_io_requestor_0_pmp_7_cfg_l = ptw_io_requestor_0_pmp_7_cfg_l;
    assign _ptw_io_requestor_0_pmp_7_cfg_res = ptw_io_requestor_0_pmp_7_cfg_res;
    assign _ptw_io_requestor_0_pmp_7_cfg_a = ptw_io_requestor_0_pmp_7_cfg_a;
    assign _ptw_io_requestor_0_pmp_7_cfg_x = ptw_io_requestor_0_pmp_7_cfg_x;
    assign _ptw_io_requestor_0_pmp_7_cfg_w = ptw_io_requestor_0_pmp_7_cfg_w;
    assign _ptw_io_requestor_0_pmp_7_cfg_r = ptw_io_requestor_0_pmp_7_cfg_r;
    assign _ptw_io_requestor_0_pmp_7_addr = ptw_io_requestor_0_pmp_7_addr;
    assign _ptw_io_requestor_0_pmp_7_mask = ptw_io_requestor_0_pmp_7_mask;
    assign _ptw_io_requestor_0_customCSRs_csrs_0_ren = ptw_io_requestor_0_customCSRs_csrs_0_ren;
    assign _ptw_io_requestor_0_customCSRs_csrs_0_wen = ptw_io_requestor_0_customCSRs_csrs_0_wen;
    assign _ptw_io_requestor_0_customCSRs_csrs_0_wdata = ptw_io_requestor_0_customCSRs_csrs_0_wdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_0_value = ptw_io_requestor_0_customCSRs_csrs_0_value;
    assign ptw_io_requestor_0_customCSRs_csrs_0_stall = _dcache_io_ptw_customCSRs_csrs_0_stall;
    assign ptw_io_requestor_0_customCSRs_csrs_0_set = _dcache_io_ptw_customCSRs_csrs_0_set;
    assign ptw_io_requestor_0_customCSRs_csrs_0_sdata = _dcache_io_ptw_customCSRs_csrs_0_sdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_1_ren = ptw_io_requestor_0_customCSRs_csrs_1_ren;
    assign _ptw_io_requestor_0_customCSRs_csrs_1_wen = ptw_io_requestor_0_customCSRs_csrs_1_wen;
    assign _ptw_io_requestor_0_customCSRs_csrs_1_wdata = ptw_io_requestor_0_customCSRs_csrs_1_wdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_1_value = ptw_io_requestor_0_customCSRs_csrs_1_value;
    assign ptw_io_requestor_0_customCSRs_csrs_1_stall = _dcache_io_ptw_customCSRs_csrs_1_stall;
    assign ptw_io_requestor_0_customCSRs_csrs_1_set = _dcache_io_ptw_customCSRs_csrs_1_set;
    assign ptw_io_requestor_0_customCSRs_csrs_1_sdata = _dcache_io_ptw_customCSRs_csrs_1_sdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_2_ren = ptw_io_requestor_0_customCSRs_csrs_2_ren;
    assign _ptw_io_requestor_0_customCSRs_csrs_2_wen = ptw_io_requestor_0_customCSRs_csrs_2_wen;
    assign _ptw_io_requestor_0_customCSRs_csrs_2_wdata = ptw_io_requestor_0_customCSRs_csrs_2_wdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_2_value = ptw_io_requestor_0_customCSRs_csrs_2_value;
    assign ptw_io_requestor_0_customCSRs_csrs_2_stall = _dcache_io_ptw_customCSRs_csrs_2_stall;
    assign ptw_io_requestor_0_customCSRs_csrs_2_set = _dcache_io_ptw_customCSRs_csrs_2_set;
    assign ptw_io_requestor_0_customCSRs_csrs_2_sdata = _dcache_io_ptw_customCSRs_csrs_2_sdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_3_ren = ptw_io_requestor_0_customCSRs_csrs_3_ren;
    assign _ptw_io_requestor_0_customCSRs_csrs_3_wen = ptw_io_requestor_0_customCSRs_csrs_3_wen;
    assign _ptw_io_requestor_0_customCSRs_csrs_3_wdata = ptw_io_requestor_0_customCSRs_csrs_3_wdata;
    assign _ptw_io_requestor_0_customCSRs_csrs_3_value = ptw_io_requestor_0_customCSRs_csrs_3_value;
    assign ptw_io_requestor_0_customCSRs_csrs_3_stall = _dcache_io_ptw_customCSRs_csrs_3_stall;
    assign ptw_io_requestor_0_customCSRs_csrs_3_set = _dcache_io_ptw_customCSRs_csrs_3_set;
    assign ptw_io_requestor_0_customCSRs_csrs_3_sdata = _dcache_io_ptw_customCSRs_csrs_3_sdata;
    assign _ptw_io_requestor_1_req_ready = ptw_io_requestor_1_req_ready;
    assign ptw_io_requestor_1_req_valid = _frontend_io_ptw_req_valid;
    assign ptw_io_requestor_1_req_bits_valid = _frontend_io_ptw_req_bits_valid;
    assign ptw_io_requestor_1_req_bits_bits_addr = _frontend_io_ptw_req_bits_bits_addr;
    assign ptw_io_requestor_1_req_bits_bits_need_gpa = _frontend_io_ptw_req_bits_bits_need_gpa;
    assign ptw_io_requestor_1_req_bits_bits_vstage1 = _frontend_io_ptw_req_bits_bits_vstage1;
    assign ptw_io_requestor_1_req_bits_bits_stage2 = _frontend_io_ptw_req_bits_bits_stage2;
    assign _ptw_io_requestor_1_resp_valid = ptw_io_requestor_1_resp_valid;
    assign _ptw_io_requestor_1_resp_bits_ae_ptw = ptw_io_requestor_1_resp_bits_ae_ptw;
    assign _ptw_io_requestor_1_resp_bits_ae_final = ptw_io_requestor_1_resp_bits_ae_final;
    assign _ptw_io_requestor_1_resp_bits_pf = ptw_io_requestor_1_resp_bits_pf;
    assign _ptw_io_requestor_1_resp_bits_gf = ptw_io_requestor_1_resp_bits_gf;
    assign _ptw_io_requestor_1_resp_bits_hr = ptw_io_requestor_1_resp_bits_hr;
    assign _ptw_io_requestor_1_resp_bits_hw = ptw_io_requestor_1_resp_bits_hw;
    assign _ptw_io_requestor_1_resp_bits_hx = ptw_io_requestor_1_resp_bits_hx;
    assign _ptw_io_requestor_1_resp_bits_pte_reserved_for_future = ptw_io_requestor_1_resp_bits_pte_reserved_for_future;
    assign _ptw_io_requestor_1_resp_bits_pte_ppn = ptw_io_requestor_1_resp_bits_pte_ppn;
    assign _ptw_io_requestor_1_resp_bits_pte_reserved_for_software = ptw_io_requestor_1_resp_bits_pte_reserved_for_software;
    assign _ptw_io_requestor_1_resp_bits_pte_d = ptw_io_requestor_1_resp_bits_pte_d;
    assign _ptw_io_requestor_1_resp_bits_pte_a = ptw_io_requestor_1_resp_bits_pte_a;
    assign _ptw_io_requestor_1_resp_bits_pte_g = ptw_io_requestor_1_resp_bits_pte_g;
    assign _ptw_io_requestor_1_resp_bits_pte_u = ptw_io_requestor_1_resp_bits_pte_u;
    assign _ptw_io_requestor_1_resp_bits_pte_x = ptw_io_requestor_1_resp_bits_pte_x;
    assign _ptw_io_requestor_1_resp_bits_pte_w = ptw_io_requestor_1_resp_bits_pte_w;
    assign _ptw_io_requestor_1_resp_bits_pte_r = ptw_io_requestor_1_resp_bits_pte_r;
    assign _ptw_io_requestor_1_resp_bits_pte_v = ptw_io_requestor_1_resp_bits_pte_v;
    assign _ptw_io_requestor_1_resp_bits_level = ptw_io_requestor_1_resp_bits_level;
    assign _ptw_io_requestor_1_resp_bits_fragmented_superpage = ptw_io_requestor_1_resp_bits_fragmented_superpage;
    assign _ptw_io_requestor_1_resp_bits_homogeneous = ptw_io_requestor_1_resp_bits_homogeneous;
    assign _ptw_io_requestor_1_resp_bits_gpa_valid = ptw_io_requestor_1_resp_bits_gpa_valid;
    assign _ptw_io_requestor_1_resp_bits_gpa_bits = ptw_io_requestor_1_resp_bits_gpa_bits;
    assign _ptw_io_requestor_1_resp_bits_gpa_is_pte = ptw_io_requestor_1_resp_bits_gpa_is_pte;
    assign _ptw_io_requestor_1_ptbr_mode = ptw_io_requestor_1_ptbr_mode;
    assign _ptw_io_requestor_1_ptbr_asid = ptw_io_requestor_1_ptbr_asid;
    assign _ptw_io_requestor_1_ptbr_ppn = ptw_io_requestor_1_ptbr_ppn;
    assign _ptw_io_requestor_1_hgatp_mode = ptw_io_requestor_1_hgatp_mode;
    assign _ptw_io_requestor_1_hgatp_asid = ptw_io_requestor_1_hgatp_asid;
    assign _ptw_io_requestor_1_hgatp_ppn = ptw_io_requestor_1_hgatp_ppn;
    assign _ptw_io_requestor_1_vsatp_mode = ptw_io_requestor_1_vsatp_mode;
    assign _ptw_io_requestor_1_vsatp_asid = ptw_io_requestor_1_vsatp_asid;
    assign _ptw_io_requestor_1_vsatp_ppn = ptw_io_requestor_1_vsatp_ppn;
    assign _ptw_io_requestor_1_status_debug = ptw_io_requestor_1_status_debug;
    assign _ptw_io_requestor_1_status_cease = ptw_io_requestor_1_status_cease;
    assign _ptw_io_requestor_1_status_wfi = ptw_io_requestor_1_status_wfi;
    assign _ptw_io_requestor_1_status_isa = ptw_io_requestor_1_status_isa;
    assign _ptw_io_requestor_1_status_dprv = ptw_io_requestor_1_status_dprv;
    assign _ptw_io_requestor_1_status_dv = ptw_io_requestor_1_status_dv;
    assign _ptw_io_requestor_1_status_prv = ptw_io_requestor_1_status_prv;
    assign _ptw_io_requestor_1_status_v = ptw_io_requestor_1_status_v;
    assign _ptw_io_requestor_1_status_sd = ptw_io_requestor_1_status_sd;
    assign _ptw_io_requestor_1_status_zero2 = ptw_io_requestor_1_status_zero2;
    assign _ptw_io_requestor_1_status_mpv = ptw_io_requestor_1_status_mpv;
    assign _ptw_io_requestor_1_status_gva = ptw_io_requestor_1_status_gva;
    assign _ptw_io_requestor_1_status_mbe = ptw_io_requestor_1_status_mbe;
    assign _ptw_io_requestor_1_status_sbe = ptw_io_requestor_1_status_sbe;
    assign _ptw_io_requestor_1_status_sxl = ptw_io_requestor_1_status_sxl;
    assign _ptw_io_requestor_1_status_uxl = ptw_io_requestor_1_status_uxl;
    assign _ptw_io_requestor_1_status_sd_rv32 = ptw_io_requestor_1_status_sd_rv32;
    assign _ptw_io_requestor_1_status_zero1 = ptw_io_requestor_1_status_zero1;
    assign _ptw_io_requestor_1_status_tsr = ptw_io_requestor_1_status_tsr;
    assign _ptw_io_requestor_1_status_tw = ptw_io_requestor_1_status_tw;
    assign _ptw_io_requestor_1_status_tvm = ptw_io_requestor_1_status_tvm;
    assign _ptw_io_requestor_1_status_mxr = ptw_io_requestor_1_status_mxr;
    assign _ptw_io_requestor_1_status_sum = ptw_io_requestor_1_status_sum;
    assign _ptw_io_requestor_1_status_mprv = ptw_io_requestor_1_status_mprv;
    assign _ptw_io_requestor_1_status_xs = ptw_io_requestor_1_status_xs;
    assign _ptw_io_requestor_1_status_fs = ptw_io_requestor_1_status_fs;
    assign _ptw_io_requestor_1_status_mpp = ptw_io_requestor_1_status_mpp;
    assign _ptw_io_requestor_1_status_vs = ptw_io_requestor_1_status_vs;
    assign _ptw_io_requestor_1_status_spp = ptw_io_requestor_1_status_spp;
    assign _ptw_io_requestor_1_status_mpie = ptw_io_requestor_1_status_mpie;
    assign _ptw_io_requestor_1_status_ube = ptw_io_requestor_1_status_ube;
    assign _ptw_io_requestor_1_status_spie = ptw_io_requestor_1_status_spie;
    assign _ptw_io_requestor_1_status_upie = ptw_io_requestor_1_status_upie;
    assign _ptw_io_requestor_1_status_mie = ptw_io_requestor_1_status_mie;
    assign _ptw_io_requestor_1_status_hie = ptw_io_requestor_1_status_hie;
    assign _ptw_io_requestor_1_status_sie = ptw_io_requestor_1_status_sie;
    assign _ptw_io_requestor_1_status_uie = ptw_io_requestor_1_status_uie;
    assign _ptw_io_requestor_1_hstatus_zero6 = ptw_io_requestor_1_hstatus_zero6;
    assign _ptw_io_requestor_1_hstatus_vsxl = ptw_io_requestor_1_hstatus_vsxl;
    assign _ptw_io_requestor_1_hstatus_zero5 = ptw_io_requestor_1_hstatus_zero5;
    assign _ptw_io_requestor_1_hstatus_vtsr = ptw_io_requestor_1_hstatus_vtsr;
    assign _ptw_io_requestor_1_hstatus_vtw = ptw_io_requestor_1_hstatus_vtw;
    assign _ptw_io_requestor_1_hstatus_vtvm = ptw_io_requestor_1_hstatus_vtvm;
    assign _ptw_io_requestor_1_hstatus_zero3 = ptw_io_requestor_1_hstatus_zero3;
    assign _ptw_io_requestor_1_hstatus_vgein = ptw_io_requestor_1_hstatus_vgein;
    assign _ptw_io_requestor_1_hstatus_zero2 = ptw_io_requestor_1_hstatus_zero2;
    assign _ptw_io_requestor_1_hstatus_hu = ptw_io_requestor_1_hstatus_hu;
    assign _ptw_io_requestor_1_hstatus_spvp = ptw_io_requestor_1_hstatus_spvp;
    assign _ptw_io_requestor_1_hstatus_spv = ptw_io_requestor_1_hstatus_spv;
    assign _ptw_io_requestor_1_hstatus_gva = ptw_io_requestor_1_hstatus_gva;
    assign _ptw_io_requestor_1_hstatus_vsbe = ptw_io_requestor_1_hstatus_vsbe;
    assign _ptw_io_requestor_1_hstatus_zero1 = ptw_io_requestor_1_hstatus_zero1;
    assign _ptw_io_requestor_1_gstatus_debug = ptw_io_requestor_1_gstatus_debug;
    assign _ptw_io_requestor_1_gstatus_cease = ptw_io_requestor_1_gstatus_cease;
    assign _ptw_io_requestor_1_gstatus_wfi = ptw_io_requestor_1_gstatus_wfi;
    assign _ptw_io_requestor_1_gstatus_isa = ptw_io_requestor_1_gstatus_isa;
    assign _ptw_io_requestor_1_gstatus_dprv = ptw_io_requestor_1_gstatus_dprv;
    assign _ptw_io_requestor_1_gstatus_dv = ptw_io_requestor_1_gstatus_dv;
    assign _ptw_io_requestor_1_gstatus_prv = ptw_io_requestor_1_gstatus_prv;
    assign _ptw_io_requestor_1_gstatus_v = ptw_io_requestor_1_gstatus_v;
    assign _ptw_io_requestor_1_gstatus_sd = ptw_io_requestor_1_gstatus_sd;
    assign _ptw_io_requestor_1_gstatus_zero2 = ptw_io_requestor_1_gstatus_zero2;
    assign _ptw_io_requestor_1_gstatus_mpv = ptw_io_requestor_1_gstatus_mpv;
    assign _ptw_io_requestor_1_gstatus_gva = ptw_io_requestor_1_gstatus_gva;
    assign _ptw_io_requestor_1_gstatus_mbe = ptw_io_requestor_1_gstatus_mbe;
    assign _ptw_io_requestor_1_gstatus_sbe = ptw_io_requestor_1_gstatus_sbe;
    assign _ptw_io_requestor_1_gstatus_sxl = ptw_io_requestor_1_gstatus_sxl;
    assign _ptw_io_requestor_1_gstatus_uxl = ptw_io_requestor_1_gstatus_uxl;
    assign _ptw_io_requestor_1_gstatus_sd_rv32 = ptw_io_requestor_1_gstatus_sd_rv32;
    assign _ptw_io_requestor_1_gstatus_zero1 = ptw_io_requestor_1_gstatus_zero1;
    assign _ptw_io_requestor_1_gstatus_tsr = ptw_io_requestor_1_gstatus_tsr;
    assign _ptw_io_requestor_1_gstatus_tw = ptw_io_requestor_1_gstatus_tw;
    assign _ptw_io_requestor_1_gstatus_tvm = ptw_io_requestor_1_gstatus_tvm;
    assign _ptw_io_requestor_1_gstatus_mxr = ptw_io_requestor_1_gstatus_mxr;
    assign _ptw_io_requestor_1_gstatus_sum = ptw_io_requestor_1_gstatus_sum;
    assign _ptw_io_requestor_1_gstatus_mprv = ptw_io_requestor_1_gstatus_mprv;
    assign _ptw_io_requestor_1_gstatus_xs = ptw_io_requestor_1_gstatus_xs;
    assign _ptw_io_requestor_1_gstatus_fs = ptw_io_requestor_1_gstatus_fs;
    assign _ptw_io_requestor_1_gstatus_mpp = ptw_io_requestor_1_gstatus_mpp;
    assign _ptw_io_requestor_1_gstatus_vs = ptw_io_requestor_1_gstatus_vs;
    assign _ptw_io_requestor_1_gstatus_spp = ptw_io_requestor_1_gstatus_spp;
    assign _ptw_io_requestor_1_gstatus_mpie = ptw_io_requestor_1_gstatus_mpie;
    assign _ptw_io_requestor_1_gstatus_ube = ptw_io_requestor_1_gstatus_ube;
    assign _ptw_io_requestor_1_gstatus_spie = ptw_io_requestor_1_gstatus_spie;
    assign _ptw_io_requestor_1_gstatus_upie = ptw_io_requestor_1_gstatus_upie;
    assign _ptw_io_requestor_1_gstatus_mie = ptw_io_requestor_1_gstatus_mie;
    assign _ptw_io_requestor_1_gstatus_hie = ptw_io_requestor_1_gstatus_hie;
    assign _ptw_io_requestor_1_gstatus_sie = ptw_io_requestor_1_gstatus_sie;
    assign _ptw_io_requestor_1_gstatus_uie = ptw_io_requestor_1_gstatus_uie;
    assign _ptw_io_requestor_1_pmp_0_cfg_l = ptw_io_requestor_1_pmp_0_cfg_l;
    assign _ptw_io_requestor_1_pmp_0_cfg_res = ptw_io_requestor_1_pmp_0_cfg_res;
    assign _ptw_io_requestor_1_pmp_0_cfg_a = ptw_io_requestor_1_pmp_0_cfg_a;
    assign _ptw_io_requestor_1_pmp_0_cfg_x = ptw_io_requestor_1_pmp_0_cfg_x;
    assign _ptw_io_requestor_1_pmp_0_cfg_w = ptw_io_requestor_1_pmp_0_cfg_w;
    assign _ptw_io_requestor_1_pmp_0_cfg_r = ptw_io_requestor_1_pmp_0_cfg_r;
    assign _ptw_io_requestor_1_pmp_0_addr = ptw_io_requestor_1_pmp_0_addr;
    assign _ptw_io_requestor_1_pmp_0_mask = ptw_io_requestor_1_pmp_0_mask;
    assign _ptw_io_requestor_1_pmp_1_cfg_l = ptw_io_requestor_1_pmp_1_cfg_l;
    assign _ptw_io_requestor_1_pmp_1_cfg_res = ptw_io_requestor_1_pmp_1_cfg_res;
    assign _ptw_io_requestor_1_pmp_1_cfg_a = ptw_io_requestor_1_pmp_1_cfg_a;
    assign _ptw_io_requestor_1_pmp_1_cfg_x = ptw_io_requestor_1_pmp_1_cfg_x;
    assign _ptw_io_requestor_1_pmp_1_cfg_w = ptw_io_requestor_1_pmp_1_cfg_w;
    assign _ptw_io_requestor_1_pmp_1_cfg_r = ptw_io_requestor_1_pmp_1_cfg_r;
    assign _ptw_io_requestor_1_pmp_1_addr = ptw_io_requestor_1_pmp_1_addr;
    assign _ptw_io_requestor_1_pmp_1_mask = ptw_io_requestor_1_pmp_1_mask;
    assign _ptw_io_requestor_1_pmp_2_cfg_l = ptw_io_requestor_1_pmp_2_cfg_l;
    assign _ptw_io_requestor_1_pmp_2_cfg_res = ptw_io_requestor_1_pmp_2_cfg_res;
    assign _ptw_io_requestor_1_pmp_2_cfg_a = ptw_io_requestor_1_pmp_2_cfg_a;
    assign _ptw_io_requestor_1_pmp_2_cfg_x = ptw_io_requestor_1_pmp_2_cfg_x;
    assign _ptw_io_requestor_1_pmp_2_cfg_w = ptw_io_requestor_1_pmp_2_cfg_w;
    assign _ptw_io_requestor_1_pmp_2_cfg_r = ptw_io_requestor_1_pmp_2_cfg_r;
    assign _ptw_io_requestor_1_pmp_2_addr = ptw_io_requestor_1_pmp_2_addr;
    assign _ptw_io_requestor_1_pmp_2_mask = ptw_io_requestor_1_pmp_2_mask;
    assign _ptw_io_requestor_1_pmp_3_cfg_l = ptw_io_requestor_1_pmp_3_cfg_l;
    assign _ptw_io_requestor_1_pmp_3_cfg_res = ptw_io_requestor_1_pmp_3_cfg_res;
    assign _ptw_io_requestor_1_pmp_3_cfg_a = ptw_io_requestor_1_pmp_3_cfg_a;
    assign _ptw_io_requestor_1_pmp_3_cfg_x = ptw_io_requestor_1_pmp_3_cfg_x;
    assign _ptw_io_requestor_1_pmp_3_cfg_w = ptw_io_requestor_1_pmp_3_cfg_w;
    assign _ptw_io_requestor_1_pmp_3_cfg_r = ptw_io_requestor_1_pmp_3_cfg_r;
    assign _ptw_io_requestor_1_pmp_3_addr = ptw_io_requestor_1_pmp_3_addr;
    assign _ptw_io_requestor_1_pmp_3_mask = ptw_io_requestor_1_pmp_3_mask;
    assign _ptw_io_requestor_1_pmp_4_cfg_l = ptw_io_requestor_1_pmp_4_cfg_l;
    assign _ptw_io_requestor_1_pmp_4_cfg_res = ptw_io_requestor_1_pmp_4_cfg_res;
    assign _ptw_io_requestor_1_pmp_4_cfg_a = ptw_io_requestor_1_pmp_4_cfg_a;
    assign _ptw_io_requestor_1_pmp_4_cfg_x = ptw_io_requestor_1_pmp_4_cfg_x;
    assign _ptw_io_requestor_1_pmp_4_cfg_w = ptw_io_requestor_1_pmp_4_cfg_w;
    assign _ptw_io_requestor_1_pmp_4_cfg_r = ptw_io_requestor_1_pmp_4_cfg_r;
    assign _ptw_io_requestor_1_pmp_4_addr = ptw_io_requestor_1_pmp_4_addr;
    assign _ptw_io_requestor_1_pmp_4_mask = ptw_io_requestor_1_pmp_4_mask;
    assign _ptw_io_requestor_1_pmp_5_cfg_l = ptw_io_requestor_1_pmp_5_cfg_l;
    assign _ptw_io_requestor_1_pmp_5_cfg_res = ptw_io_requestor_1_pmp_5_cfg_res;
    assign _ptw_io_requestor_1_pmp_5_cfg_a = ptw_io_requestor_1_pmp_5_cfg_a;
    assign _ptw_io_requestor_1_pmp_5_cfg_x = ptw_io_requestor_1_pmp_5_cfg_x;
    assign _ptw_io_requestor_1_pmp_5_cfg_w = ptw_io_requestor_1_pmp_5_cfg_w;
    assign _ptw_io_requestor_1_pmp_5_cfg_r = ptw_io_requestor_1_pmp_5_cfg_r;
    assign _ptw_io_requestor_1_pmp_5_addr = ptw_io_requestor_1_pmp_5_addr;
    assign _ptw_io_requestor_1_pmp_5_mask = ptw_io_requestor_1_pmp_5_mask;
    assign _ptw_io_requestor_1_pmp_6_cfg_l = ptw_io_requestor_1_pmp_6_cfg_l;
    assign _ptw_io_requestor_1_pmp_6_cfg_res = ptw_io_requestor_1_pmp_6_cfg_res;
    assign _ptw_io_requestor_1_pmp_6_cfg_a = ptw_io_requestor_1_pmp_6_cfg_a;
    assign _ptw_io_requestor_1_pmp_6_cfg_x = ptw_io_requestor_1_pmp_6_cfg_x;
    assign _ptw_io_requestor_1_pmp_6_cfg_w = ptw_io_requestor_1_pmp_6_cfg_w;
    assign _ptw_io_requestor_1_pmp_6_cfg_r = ptw_io_requestor_1_pmp_6_cfg_r;
    assign _ptw_io_requestor_1_pmp_6_addr = ptw_io_requestor_1_pmp_6_addr;
    assign _ptw_io_requestor_1_pmp_6_mask = ptw_io_requestor_1_pmp_6_mask;
    assign _ptw_io_requestor_1_pmp_7_cfg_l = ptw_io_requestor_1_pmp_7_cfg_l;
    assign _ptw_io_requestor_1_pmp_7_cfg_res = ptw_io_requestor_1_pmp_7_cfg_res;
    assign _ptw_io_requestor_1_pmp_7_cfg_a = ptw_io_requestor_1_pmp_7_cfg_a;
    assign _ptw_io_requestor_1_pmp_7_cfg_x = ptw_io_requestor_1_pmp_7_cfg_x;
    assign _ptw_io_requestor_1_pmp_7_cfg_w = ptw_io_requestor_1_pmp_7_cfg_w;
    assign _ptw_io_requestor_1_pmp_7_cfg_r = ptw_io_requestor_1_pmp_7_cfg_r;
    assign _ptw_io_requestor_1_pmp_7_addr = ptw_io_requestor_1_pmp_7_addr;
    assign _ptw_io_requestor_1_pmp_7_mask = ptw_io_requestor_1_pmp_7_mask;
    assign _ptw_io_requestor_1_customCSRs_csrs_0_ren = ptw_io_requestor_1_customCSRs_csrs_0_ren;
    assign _ptw_io_requestor_1_customCSRs_csrs_0_wen = ptw_io_requestor_1_customCSRs_csrs_0_wen;
    assign _ptw_io_requestor_1_customCSRs_csrs_0_wdata = ptw_io_requestor_1_customCSRs_csrs_0_wdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_0_value = ptw_io_requestor_1_customCSRs_csrs_0_value;
    assign ptw_io_requestor_1_customCSRs_csrs_0_stall = _frontend_io_ptw_customCSRs_csrs_0_stall;
    assign ptw_io_requestor_1_customCSRs_csrs_0_set = _frontend_io_ptw_customCSRs_csrs_0_set;
    assign ptw_io_requestor_1_customCSRs_csrs_0_sdata = _frontend_io_ptw_customCSRs_csrs_0_sdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_1_ren = ptw_io_requestor_1_customCSRs_csrs_1_ren;
    assign _ptw_io_requestor_1_customCSRs_csrs_1_wen = ptw_io_requestor_1_customCSRs_csrs_1_wen;
    assign _ptw_io_requestor_1_customCSRs_csrs_1_wdata = ptw_io_requestor_1_customCSRs_csrs_1_wdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_1_value = ptw_io_requestor_1_customCSRs_csrs_1_value;
    assign ptw_io_requestor_1_customCSRs_csrs_1_stall = _frontend_io_ptw_customCSRs_csrs_1_stall;
    assign ptw_io_requestor_1_customCSRs_csrs_1_set = _frontend_io_ptw_customCSRs_csrs_1_set;
    assign ptw_io_requestor_1_customCSRs_csrs_1_sdata = _frontend_io_ptw_customCSRs_csrs_1_sdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_2_ren = ptw_io_requestor_1_customCSRs_csrs_2_ren;
    assign _ptw_io_requestor_1_customCSRs_csrs_2_wen = ptw_io_requestor_1_customCSRs_csrs_2_wen;
    assign _ptw_io_requestor_1_customCSRs_csrs_2_wdata = ptw_io_requestor_1_customCSRs_csrs_2_wdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_2_value = ptw_io_requestor_1_customCSRs_csrs_2_value;
    assign ptw_io_requestor_1_customCSRs_csrs_2_stall = _frontend_io_ptw_customCSRs_csrs_2_stall;
    assign ptw_io_requestor_1_customCSRs_csrs_2_set = _frontend_io_ptw_customCSRs_csrs_2_set;
    assign ptw_io_requestor_1_customCSRs_csrs_2_sdata = _frontend_io_ptw_customCSRs_csrs_2_sdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_3_ren = ptw_io_requestor_1_customCSRs_csrs_3_ren;
    assign _ptw_io_requestor_1_customCSRs_csrs_3_wen = ptw_io_requestor_1_customCSRs_csrs_3_wen;
    assign _ptw_io_requestor_1_customCSRs_csrs_3_wdata = ptw_io_requestor_1_customCSRs_csrs_3_wdata;
    assign _ptw_io_requestor_1_customCSRs_csrs_3_value = ptw_io_requestor_1_customCSRs_csrs_3_value;
    assign ptw_io_requestor_1_customCSRs_csrs_3_stall = _frontend_io_ptw_customCSRs_csrs_3_stall;
    assign ptw_io_requestor_1_customCSRs_csrs_3_set = _frontend_io_ptw_customCSRs_csrs_3_set;
    assign ptw_io_requestor_1_customCSRs_csrs_3_sdata = _frontend_io_ptw_customCSRs_csrs_3_sdata;
    assign ptw_io_mem_req_ready = 1'h0;
    assign ptw_io_mem_s2_nack = 1'h0;
    assign ptw_io_mem_s2_nack_cause_raw = 1'h0;
    assign ptw_io_mem_s2_uncached = 1'h0;
    assign ptw_io_mem_s2_paddr = 32'h0;
    assign ptw_io_mem_resp_valid = 1'h0;
    assign ptw_io_mem_resp_bits_addr = 34'h0;
    assign ptw_io_mem_resp_bits_tag = 6'h0;
    assign ptw_io_mem_resp_bits_cmd = 5'h0;
    assign ptw_io_mem_resp_bits_size = 2'h0;
    assign ptw_io_mem_resp_bits_signed = 1'h0;
    assign ptw_io_mem_resp_bits_dprv = 2'h0;
    assign ptw_io_mem_resp_bits_dv = 1'h0;
    assign ptw_io_mem_resp_bits_data = 64'h0;
    assign ptw_io_mem_resp_bits_mask = 8'h0;
    assign ptw_io_mem_resp_bits_replay = 1'h0;
    assign ptw_io_mem_resp_bits_has_data = 1'h0;
    assign ptw_io_mem_resp_bits_data_word_bypass = 64'h0;
    assign ptw_io_mem_resp_bits_data_raw = 64'h0;
    assign ptw_io_mem_resp_bits_store_data = 64'h0;
    assign ptw_io_mem_replay_next = 1'h0;
    assign ptw_io_mem_s2_xcpt_ma_ld = 1'h0;
    assign ptw_io_mem_s2_xcpt_ma_st = 1'h0;
    assign ptw_io_mem_s2_xcpt_pf_ld = 1'h0;
    assign ptw_io_mem_s2_xcpt_pf_st = 1'h0;
    assign ptw_io_mem_s2_xcpt_gf_ld = 1'h0;
    assign ptw_io_mem_s2_xcpt_gf_st = 1'h0;
    assign ptw_io_mem_s2_xcpt_ae_ld = 1'h0;
    assign ptw_io_mem_s2_xcpt_ae_st = 1'h0;
    assign ptw_io_mem_s2_gpa = 34'h0;
    assign ptw_io_mem_s2_gpa_is_pte = 1'h0;
    assign ptw_io_mem_ordered = 1'h0;
    assign ptw_io_mem_perf_acquire = 1'h0;
    assign ptw_io_mem_perf_release = 1'h0;
    assign ptw_io_mem_perf_grant = 1'h0;
    assign ptw_io_mem_perf_tlbMiss = 1'h0;
    assign ptw_io_mem_perf_blocked = 1'h0;
    assign ptw_io_mem_perf_canAcceptStoreThenLoad = 1'h0;
    assign ptw_io_mem_perf_canAcceptStoreThenRMW = 1'h0;
    assign ptw_io_mem_perf_canAcceptLoadThenLoad = 1'h0;
    assign ptw_io_mem_perf_storeBufferEmptyAfterLoad = 1'h0;
    assign ptw_io_mem_perf_storeBufferEmptyAfterStore = 1'h0;
    assign ptw_io_mem_clock_enabled = 1'h0;
    assign ptw_io_dpath_ptbr_mode = _core_io_ptw_ptbr_mode;
    assign ptw_io_dpath_ptbr_asid = _core_io_ptw_ptbr_asid;
    assign ptw_io_dpath_ptbr_ppn = _core_io_ptw_ptbr_ppn;
    assign ptw_io_dpath_hgatp_mode = _core_io_ptw_hgatp_mode;
    assign ptw_io_dpath_hgatp_asid = _core_io_ptw_hgatp_asid;
    assign ptw_io_dpath_hgatp_ppn = _core_io_ptw_hgatp_ppn;
    assign ptw_io_dpath_vsatp_mode = _core_io_ptw_vsatp_mode;
    assign ptw_io_dpath_vsatp_asid = _core_io_ptw_vsatp_asid;
    assign ptw_io_dpath_vsatp_ppn = _core_io_ptw_vsatp_ppn;
    assign ptw_io_dpath_sfence_valid = _core_io_ptw_sfence_valid;
    assign ptw_io_dpath_sfence_bits_rs1 = _core_io_ptw_sfence_bits_rs1;
    assign ptw_io_dpath_sfence_bits_rs2 = _core_io_ptw_sfence_bits_rs2;
    assign ptw_io_dpath_sfence_bits_addr = _core_io_ptw_sfence_bits_addr;
    assign ptw_io_dpath_sfence_bits_asid = _core_io_ptw_sfence_bits_asid;
    assign ptw_io_dpath_sfence_bits_hv = _core_io_ptw_sfence_bits_hv;
    assign ptw_io_dpath_sfence_bits_hg = _core_io_ptw_sfence_bits_hg;
    assign ptw_io_dpath_status_debug = _core_io_ptw_status_debug;
    assign ptw_io_dpath_status_cease = _core_io_ptw_status_cease;
    assign ptw_io_dpath_status_wfi = _core_io_ptw_status_wfi;
    assign ptw_io_dpath_status_isa = _core_io_ptw_status_isa;
    assign ptw_io_dpath_status_dprv = _core_io_ptw_status_dprv;
    assign ptw_io_dpath_status_dv = _core_io_ptw_status_dv;
    assign ptw_io_dpath_status_prv = _core_io_ptw_status_prv;
    assign ptw_io_dpath_status_v = _core_io_ptw_status_v;
    assign ptw_io_dpath_status_sd = _core_io_ptw_status_sd;
    assign ptw_io_dpath_status_zero2 = _core_io_ptw_status_zero2;
    assign ptw_io_dpath_status_mpv = _core_io_ptw_status_mpv;
    assign ptw_io_dpath_status_gva = _core_io_ptw_status_gva;
    assign ptw_io_dpath_status_mbe = _core_io_ptw_status_mbe;
    assign ptw_io_dpath_status_sbe = _core_io_ptw_status_sbe;
    assign ptw_io_dpath_status_sxl = _core_io_ptw_status_sxl;
    assign ptw_io_dpath_status_uxl = _core_io_ptw_status_uxl;
    assign ptw_io_dpath_status_sd_rv32 = _core_io_ptw_status_sd_rv32;
    assign ptw_io_dpath_status_zero1 = _core_io_ptw_status_zero1;
    assign ptw_io_dpath_status_tsr = _core_io_ptw_status_tsr;
    assign ptw_io_dpath_status_tw = _core_io_ptw_status_tw;
    assign ptw_io_dpath_status_tvm = _core_io_ptw_status_tvm;
    assign ptw_io_dpath_status_mxr = _core_io_ptw_status_mxr;
    assign ptw_io_dpath_status_sum = _core_io_ptw_status_sum;
    assign ptw_io_dpath_status_mprv = _core_io_ptw_status_mprv;
    assign ptw_io_dpath_status_xs = _core_io_ptw_status_xs;
    assign ptw_io_dpath_status_fs = _core_io_ptw_status_fs;
    assign ptw_io_dpath_status_mpp = _core_io_ptw_status_mpp;
    assign ptw_io_dpath_status_vs = _core_io_ptw_status_vs;
    assign ptw_io_dpath_status_spp = _core_io_ptw_status_spp;
    assign ptw_io_dpath_status_mpie = _core_io_ptw_status_mpie;
    assign ptw_io_dpath_status_ube = _core_io_ptw_status_ube;
    assign ptw_io_dpath_status_spie = _core_io_ptw_status_spie;
    assign ptw_io_dpath_status_upie = _core_io_ptw_status_upie;
    assign ptw_io_dpath_status_mie = _core_io_ptw_status_mie;
    assign ptw_io_dpath_status_hie = _core_io_ptw_status_hie;
    assign ptw_io_dpath_status_sie = _core_io_ptw_status_sie;
    assign ptw_io_dpath_status_uie = _core_io_ptw_status_uie;
    assign ptw_io_dpath_hstatus_zero6 = _core_io_ptw_hstatus_zero6;
    assign ptw_io_dpath_hstatus_vsxl = _core_io_ptw_hstatus_vsxl;
    assign ptw_io_dpath_hstatus_zero5 = _core_io_ptw_hstatus_zero5;
    assign ptw_io_dpath_hstatus_vtsr = _core_io_ptw_hstatus_vtsr;
    assign ptw_io_dpath_hstatus_vtw = _core_io_ptw_hstatus_vtw;
    assign ptw_io_dpath_hstatus_vtvm = _core_io_ptw_hstatus_vtvm;
    assign ptw_io_dpath_hstatus_zero3 = _core_io_ptw_hstatus_zero3;
    assign ptw_io_dpath_hstatus_vgein = _core_io_ptw_hstatus_vgein;
    assign ptw_io_dpath_hstatus_zero2 = _core_io_ptw_hstatus_zero2;
    assign ptw_io_dpath_hstatus_hu = _core_io_ptw_hstatus_hu;
    assign ptw_io_dpath_hstatus_spvp = _core_io_ptw_hstatus_spvp;
    assign ptw_io_dpath_hstatus_spv = _core_io_ptw_hstatus_spv;
    assign ptw_io_dpath_hstatus_gva = _core_io_ptw_hstatus_gva;
    assign ptw_io_dpath_hstatus_vsbe = _core_io_ptw_hstatus_vsbe;
    assign ptw_io_dpath_hstatus_zero1 = _core_io_ptw_hstatus_zero1;
    assign ptw_io_dpath_gstatus_debug = _core_io_ptw_gstatus_debug;
    assign ptw_io_dpath_gstatus_cease = _core_io_ptw_gstatus_cease;
    assign ptw_io_dpath_gstatus_wfi = _core_io_ptw_gstatus_wfi;
    assign ptw_io_dpath_gstatus_isa = _core_io_ptw_gstatus_isa;
    assign ptw_io_dpath_gstatus_dprv = _core_io_ptw_gstatus_dprv;
    assign ptw_io_dpath_gstatus_dv = _core_io_ptw_gstatus_dv;
    assign ptw_io_dpath_gstatus_prv = _core_io_ptw_gstatus_prv;
    assign ptw_io_dpath_gstatus_v = _core_io_ptw_gstatus_v;
    assign ptw_io_dpath_gstatus_sd = _core_io_ptw_gstatus_sd;
    assign ptw_io_dpath_gstatus_zero2 = _core_io_ptw_gstatus_zero2;
    assign ptw_io_dpath_gstatus_mpv = _core_io_ptw_gstatus_mpv;
    assign ptw_io_dpath_gstatus_gva = _core_io_ptw_gstatus_gva;
    assign ptw_io_dpath_gstatus_mbe = _core_io_ptw_gstatus_mbe;
    assign ptw_io_dpath_gstatus_sbe = _core_io_ptw_gstatus_sbe;
    assign ptw_io_dpath_gstatus_sxl = _core_io_ptw_gstatus_sxl;
    assign ptw_io_dpath_gstatus_uxl = _core_io_ptw_gstatus_uxl;
    assign ptw_io_dpath_gstatus_sd_rv32 = _core_io_ptw_gstatus_sd_rv32;
    assign ptw_io_dpath_gstatus_zero1 = _core_io_ptw_gstatus_zero1;
    assign ptw_io_dpath_gstatus_tsr = _core_io_ptw_gstatus_tsr;
    assign ptw_io_dpath_gstatus_tw = _core_io_ptw_gstatus_tw;
    assign ptw_io_dpath_gstatus_tvm = _core_io_ptw_gstatus_tvm;
    assign ptw_io_dpath_gstatus_mxr = _core_io_ptw_gstatus_mxr;
    assign ptw_io_dpath_gstatus_sum = _core_io_ptw_gstatus_sum;
    assign ptw_io_dpath_gstatus_mprv = _core_io_ptw_gstatus_mprv;
    assign ptw_io_dpath_gstatus_xs = _core_io_ptw_gstatus_xs;
    assign ptw_io_dpath_gstatus_fs = _core_io_ptw_gstatus_fs;
    assign ptw_io_dpath_gstatus_mpp = _core_io_ptw_gstatus_mpp;
    assign ptw_io_dpath_gstatus_vs = _core_io_ptw_gstatus_vs;
    assign ptw_io_dpath_gstatus_spp = _core_io_ptw_gstatus_spp;
    assign ptw_io_dpath_gstatus_mpie = _core_io_ptw_gstatus_mpie;
    assign ptw_io_dpath_gstatus_ube = _core_io_ptw_gstatus_ube;
    assign ptw_io_dpath_gstatus_spie = _core_io_ptw_gstatus_spie;
    assign ptw_io_dpath_gstatus_upie = _core_io_ptw_gstatus_upie;
    assign ptw_io_dpath_gstatus_mie = _core_io_ptw_gstatus_mie;
    assign ptw_io_dpath_gstatus_hie = _core_io_ptw_gstatus_hie;
    assign ptw_io_dpath_gstatus_sie = _core_io_ptw_gstatus_sie;
    assign ptw_io_dpath_gstatus_uie = _core_io_ptw_gstatus_uie;
    assign ptw_io_dpath_pmp_0_cfg_l = _core_io_ptw_pmp_0_cfg_l;
    assign ptw_io_dpath_pmp_0_cfg_res = _core_io_ptw_pmp_0_cfg_res;
    assign ptw_io_dpath_pmp_0_cfg_a = _core_io_ptw_pmp_0_cfg_a;
    assign ptw_io_dpath_pmp_0_cfg_x = _core_io_ptw_pmp_0_cfg_x;
    assign ptw_io_dpath_pmp_0_cfg_w = _core_io_ptw_pmp_0_cfg_w;
    assign ptw_io_dpath_pmp_0_cfg_r = _core_io_ptw_pmp_0_cfg_r;
    assign ptw_io_dpath_pmp_0_addr = _core_io_ptw_pmp_0_addr;
    assign ptw_io_dpath_pmp_0_mask = _core_io_ptw_pmp_0_mask;
    assign ptw_io_dpath_pmp_1_cfg_l = _core_io_ptw_pmp_1_cfg_l;
    assign ptw_io_dpath_pmp_1_cfg_res = _core_io_ptw_pmp_1_cfg_res;
    assign ptw_io_dpath_pmp_1_cfg_a = _core_io_ptw_pmp_1_cfg_a;
    assign ptw_io_dpath_pmp_1_cfg_x = _core_io_ptw_pmp_1_cfg_x;
    assign ptw_io_dpath_pmp_1_cfg_w = _core_io_ptw_pmp_1_cfg_w;
    assign ptw_io_dpath_pmp_1_cfg_r = _core_io_ptw_pmp_1_cfg_r;
    assign ptw_io_dpath_pmp_1_addr = _core_io_ptw_pmp_1_addr;
    assign ptw_io_dpath_pmp_1_mask = _core_io_ptw_pmp_1_mask;
    assign ptw_io_dpath_pmp_2_cfg_l = _core_io_ptw_pmp_2_cfg_l;
    assign ptw_io_dpath_pmp_2_cfg_res = _core_io_ptw_pmp_2_cfg_res;
    assign ptw_io_dpath_pmp_2_cfg_a = _core_io_ptw_pmp_2_cfg_a;
    assign ptw_io_dpath_pmp_2_cfg_x = _core_io_ptw_pmp_2_cfg_x;
    assign ptw_io_dpath_pmp_2_cfg_w = _core_io_ptw_pmp_2_cfg_w;
    assign ptw_io_dpath_pmp_2_cfg_r = _core_io_ptw_pmp_2_cfg_r;
    assign ptw_io_dpath_pmp_2_addr = _core_io_ptw_pmp_2_addr;
    assign ptw_io_dpath_pmp_2_mask = _core_io_ptw_pmp_2_mask;
    assign ptw_io_dpath_pmp_3_cfg_l = _core_io_ptw_pmp_3_cfg_l;
    assign ptw_io_dpath_pmp_3_cfg_res = _core_io_ptw_pmp_3_cfg_res;
    assign ptw_io_dpath_pmp_3_cfg_a = _core_io_ptw_pmp_3_cfg_a;
    assign ptw_io_dpath_pmp_3_cfg_x = _core_io_ptw_pmp_3_cfg_x;
    assign ptw_io_dpath_pmp_3_cfg_w = _core_io_ptw_pmp_3_cfg_w;
    assign ptw_io_dpath_pmp_3_cfg_r = _core_io_ptw_pmp_3_cfg_r;
    assign ptw_io_dpath_pmp_3_addr = _core_io_ptw_pmp_3_addr;
    assign ptw_io_dpath_pmp_3_mask = _core_io_ptw_pmp_3_mask;
    assign ptw_io_dpath_pmp_4_cfg_l = _core_io_ptw_pmp_4_cfg_l;
    assign ptw_io_dpath_pmp_4_cfg_res = _core_io_ptw_pmp_4_cfg_res;
    assign ptw_io_dpath_pmp_4_cfg_a = _core_io_ptw_pmp_4_cfg_a;
    assign ptw_io_dpath_pmp_4_cfg_x = _core_io_ptw_pmp_4_cfg_x;
    assign ptw_io_dpath_pmp_4_cfg_w = _core_io_ptw_pmp_4_cfg_w;
    assign ptw_io_dpath_pmp_4_cfg_r = _core_io_ptw_pmp_4_cfg_r;
    assign ptw_io_dpath_pmp_4_addr = _core_io_ptw_pmp_4_addr;
    assign ptw_io_dpath_pmp_4_mask = _core_io_ptw_pmp_4_mask;
    assign ptw_io_dpath_pmp_5_cfg_l = _core_io_ptw_pmp_5_cfg_l;
    assign ptw_io_dpath_pmp_5_cfg_res = _core_io_ptw_pmp_5_cfg_res;
    assign ptw_io_dpath_pmp_5_cfg_a = _core_io_ptw_pmp_5_cfg_a;
    assign ptw_io_dpath_pmp_5_cfg_x = _core_io_ptw_pmp_5_cfg_x;
    assign ptw_io_dpath_pmp_5_cfg_w = _core_io_ptw_pmp_5_cfg_w;
    assign ptw_io_dpath_pmp_5_cfg_r = _core_io_ptw_pmp_5_cfg_r;
    assign ptw_io_dpath_pmp_5_addr = _core_io_ptw_pmp_5_addr;
    assign ptw_io_dpath_pmp_5_mask = _core_io_ptw_pmp_5_mask;
    assign ptw_io_dpath_pmp_6_cfg_l = _core_io_ptw_pmp_6_cfg_l;
    assign ptw_io_dpath_pmp_6_cfg_res = _core_io_ptw_pmp_6_cfg_res;
    assign ptw_io_dpath_pmp_6_cfg_a = _core_io_ptw_pmp_6_cfg_a;
    assign ptw_io_dpath_pmp_6_cfg_x = _core_io_ptw_pmp_6_cfg_x;
    assign ptw_io_dpath_pmp_6_cfg_w = _core_io_ptw_pmp_6_cfg_w;
    assign ptw_io_dpath_pmp_6_cfg_r = _core_io_ptw_pmp_6_cfg_r;
    assign ptw_io_dpath_pmp_6_addr = _core_io_ptw_pmp_6_addr;
    assign ptw_io_dpath_pmp_6_mask = _core_io_ptw_pmp_6_mask;
    assign ptw_io_dpath_pmp_7_cfg_l = _core_io_ptw_pmp_7_cfg_l;
    assign ptw_io_dpath_pmp_7_cfg_res = _core_io_ptw_pmp_7_cfg_res;
    assign ptw_io_dpath_pmp_7_cfg_a = _core_io_ptw_pmp_7_cfg_a;
    assign ptw_io_dpath_pmp_7_cfg_x = _core_io_ptw_pmp_7_cfg_x;
    assign ptw_io_dpath_pmp_7_cfg_w = _core_io_ptw_pmp_7_cfg_w;
    assign ptw_io_dpath_pmp_7_cfg_r = _core_io_ptw_pmp_7_cfg_r;
    assign ptw_io_dpath_pmp_7_addr = _core_io_ptw_pmp_7_addr;
    assign ptw_io_dpath_pmp_7_mask = _core_io_ptw_pmp_7_mask;
    assign _ptw_io_dpath_perf_l2miss = ptw_io_dpath_perf_l2miss;
    assign _ptw_io_dpath_perf_l2hit = ptw_io_dpath_perf_l2hit;
    assign _ptw_io_dpath_perf_pte_miss = ptw_io_dpath_perf_pte_miss;
    assign _ptw_io_dpath_perf_pte_hit = ptw_io_dpath_perf_pte_hit;
    assign ptw_io_dpath_customCSRs_csrs_0_ren = _core_io_ptw_customCSRs_csrs_0_ren;
    assign ptw_io_dpath_customCSRs_csrs_0_wen = _core_io_ptw_customCSRs_csrs_0_wen;
    assign ptw_io_dpath_customCSRs_csrs_0_wdata = _core_io_ptw_customCSRs_csrs_0_wdata;
    assign ptw_io_dpath_customCSRs_csrs_0_value = _core_io_ptw_customCSRs_csrs_0_value;
    assign _ptw_io_dpath_customCSRs_csrs_0_stall = ptw_io_dpath_customCSRs_csrs_0_stall;
    assign _ptw_io_dpath_customCSRs_csrs_0_set = ptw_io_dpath_customCSRs_csrs_0_set;
    assign _ptw_io_dpath_customCSRs_csrs_0_sdata = ptw_io_dpath_customCSRs_csrs_0_sdata;
    assign ptw_io_dpath_customCSRs_csrs_1_ren = _core_io_ptw_customCSRs_csrs_1_ren;
    assign ptw_io_dpath_customCSRs_csrs_1_wen = _core_io_ptw_customCSRs_csrs_1_wen;
    assign ptw_io_dpath_customCSRs_csrs_1_wdata = _core_io_ptw_customCSRs_csrs_1_wdata;
    assign ptw_io_dpath_customCSRs_csrs_1_value = _core_io_ptw_customCSRs_csrs_1_value;
    assign _ptw_io_dpath_customCSRs_csrs_1_stall = ptw_io_dpath_customCSRs_csrs_1_stall;
    assign _ptw_io_dpath_customCSRs_csrs_1_set = ptw_io_dpath_customCSRs_csrs_1_set;
    assign _ptw_io_dpath_customCSRs_csrs_1_sdata = ptw_io_dpath_customCSRs_csrs_1_sdata;
    assign ptw_io_dpath_customCSRs_csrs_2_ren = _core_io_ptw_customCSRs_csrs_2_ren;
    assign ptw_io_dpath_customCSRs_csrs_2_wen = _core_io_ptw_customCSRs_csrs_2_wen;
    assign ptw_io_dpath_customCSRs_csrs_2_wdata = _core_io_ptw_customCSRs_csrs_2_wdata;
    assign ptw_io_dpath_customCSRs_csrs_2_value = _core_io_ptw_customCSRs_csrs_2_value;
    assign _ptw_io_dpath_customCSRs_csrs_2_stall = ptw_io_dpath_customCSRs_csrs_2_stall;
    assign _ptw_io_dpath_customCSRs_csrs_2_set = ptw_io_dpath_customCSRs_csrs_2_set;
    assign _ptw_io_dpath_customCSRs_csrs_2_sdata = ptw_io_dpath_customCSRs_csrs_2_sdata;
    assign ptw_io_dpath_customCSRs_csrs_3_ren = _core_io_ptw_customCSRs_csrs_3_ren;
    assign ptw_io_dpath_customCSRs_csrs_3_wen = _core_io_ptw_customCSRs_csrs_3_wen;
    assign ptw_io_dpath_customCSRs_csrs_3_wdata = _core_io_ptw_customCSRs_csrs_3_wdata;
    assign ptw_io_dpath_customCSRs_csrs_3_value = _core_io_ptw_customCSRs_csrs_3_value;
    assign _ptw_io_dpath_customCSRs_csrs_3_stall = ptw_io_dpath_customCSRs_csrs_3_stall;
    assign _ptw_io_dpath_customCSRs_csrs_3_set = ptw_io_dpath_customCSRs_csrs_3_set;
    assign _ptw_io_dpath_customCSRs_csrs_3_sdata = ptw_io_dpath_customCSRs_csrs_3_sdata;
    assign _ptw_io_dpath_clock_enabled = ptw_io_dpath_clock_enabled;
    
  wire core_clock;
    wire core_reset;
    wire core_io_hartid;
    wire[31:0] core_io_reset_vector;
    wire core_io_interrupts_debug;
    wire core_io_interrupts_mtip;
    wire core_io_interrupts_msip;
    wire core_io_interrupts_meip;
    wire core_io_imem_might_request;
    wire core_io_imem_clock_enabled;
    wire core_io_imem_req_valid;
    wire[33:0] core_io_imem_req_bits_pc;
    wire core_io_imem_req_bits_speculative;
    wire core_io_imem_sfence_valid;
    wire core_io_imem_sfence_bits_rs1;
    wire core_io_imem_sfence_bits_rs2;
    wire[32:0] core_io_imem_sfence_bits_addr;
    wire core_io_imem_sfence_bits_asid;
    wire core_io_imem_sfence_bits_hv;
    wire core_io_imem_sfence_bits_hg;
    wire core_io_imem_resp_ready;
    wire core_io_imem_resp_valid;
    wire[1:0] core_io_imem_resp_bits_btb_cfiType;
    wire core_io_imem_resp_bits_btb_taken;
    wire[1:0] core_io_imem_resp_bits_btb_mask;
    wire core_io_imem_resp_bits_btb_bridx;
    wire[32:0] core_io_imem_resp_bits_btb_target;
    wire core_io_imem_resp_bits_btb_entry;
    wire[7:0] core_io_imem_resp_bits_btb_bht_history;
    wire core_io_imem_resp_bits_btb_bht_value;
    wire[33:0] core_io_imem_resp_bits_pc;
    wire[31:0] core_io_imem_resp_bits_data;
    wire[1:0] core_io_imem_resp_bits_mask;
    wire core_io_imem_resp_bits_xcpt_pf_inst;
    wire core_io_imem_resp_bits_xcpt_gf_inst;
    wire core_io_imem_resp_bits_xcpt_ae_inst;
    wire core_io_imem_resp_bits_replay;
    wire core_io_imem_gpa_valid;
    wire[33:0] core_io_imem_gpa_bits;
    wire core_io_imem_btb_update_valid;
    wire[1:0] core_io_imem_btb_update_bits_prediction_cfiType;
    wire core_io_imem_btb_update_bits_prediction_taken;
    wire[1:0] core_io_imem_btb_update_bits_prediction_mask;
    wire core_io_imem_btb_update_bits_prediction_bridx;
    wire[32:0] core_io_imem_btb_update_bits_prediction_target;
    wire core_io_imem_btb_update_bits_prediction_entry;
    wire[7:0] core_io_imem_btb_update_bits_prediction_bht_history;
    wire core_io_imem_btb_update_bits_prediction_bht_value;
    wire[32:0] core_io_imem_btb_update_bits_pc;
    wire[32:0] core_io_imem_btb_update_bits_target;
    wire core_io_imem_btb_update_bits_taken;
    wire core_io_imem_btb_update_bits_isValid;
    wire[32:0] core_io_imem_btb_update_bits_br_pc;
    wire[1:0] core_io_imem_btb_update_bits_cfiType;
    wire core_io_imem_bht_update_valid;
    wire[7:0] core_io_imem_bht_update_bits_prediction_history;
    wire core_io_imem_bht_update_bits_prediction_value;
    wire[32:0] core_io_imem_bht_update_bits_pc;
    wire core_io_imem_bht_update_bits_branch;
    wire core_io_imem_bht_update_bits_taken;
    wire core_io_imem_bht_update_bits_mispredict;
    wire core_io_imem_ras_update_valid;
    wire[1:0] core_io_imem_ras_update_bits_cfiType;
    wire[32:0] core_io_imem_ras_update_bits_returnAddr;
    wire core_io_imem_flush_icache;
    wire[33:0] core_io_imem_npc;
    wire core_io_imem_perf_acquire;
    wire core_io_imem_perf_tlbMiss;
    wire core_io_imem_progress;
    wire core_io_dmem_req_ready;
    wire core_io_dmem_req_valid;
    wire[33:0] core_io_dmem_req_bits_addr;
    wire[5:0] core_io_dmem_req_bits_tag;
    wire[4:0] core_io_dmem_req_bits_cmd;
    wire[1:0] core_io_dmem_req_bits_size;
    wire core_io_dmem_req_bits_signed;
    wire[1:0] core_io_dmem_req_bits_dprv;
    wire core_io_dmem_req_bits_dv;
    wire core_io_dmem_req_bits_phys;
    wire core_io_dmem_req_bits_no_alloc;
    wire core_io_dmem_req_bits_no_xcpt;
    wire[63:0] core_io_dmem_req_bits_data;
    wire[7:0] core_io_dmem_req_bits_mask;
    wire core_io_dmem_s1_kill;
    wire[63:0] core_io_dmem_s1_data_data;
    wire[7:0] core_io_dmem_s1_data_mask;
    wire core_io_dmem_s2_nack;
    wire core_io_dmem_s2_nack_cause_raw;
    wire core_io_dmem_s2_kill;
    wire core_io_dmem_s2_uncached;
    wire[31:0] core_io_dmem_s2_paddr;
    wire core_io_dmem_resp_valid;
    wire[33:0] core_io_dmem_resp_bits_addr;
    wire[5:0] core_io_dmem_resp_bits_tag;
    wire[4:0] core_io_dmem_resp_bits_cmd;
    wire[1:0] core_io_dmem_resp_bits_size;
    wire core_io_dmem_resp_bits_signed;
    wire[1:0] core_io_dmem_resp_bits_dprv;
    wire core_io_dmem_resp_bits_dv;
    wire[63:0] core_io_dmem_resp_bits_data;
    wire[7:0] core_io_dmem_resp_bits_mask;
    wire core_io_dmem_resp_bits_replay;
    wire core_io_dmem_resp_bits_has_data;
    wire[63:0] core_io_dmem_resp_bits_data_word_bypass;
    wire[63:0] core_io_dmem_resp_bits_data_raw;
    wire[63:0] core_io_dmem_resp_bits_store_data;
    wire core_io_dmem_replay_next;
    wire core_io_dmem_s2_xcpt_ma_ld;
    wire core_io_dmem_s2_xcpt_ma_st;
    wire core_io_dmem_s2_xcpt_pf_ld;
    wire core_io_dmem_s2_xcpt_pf_st;
    wire core_io_dmem_s2_xcpt_gf_ld;
    wire core_io_dmem_s2_xcpt_gf_st;
    wire core_io_dmem_s2_xcpt_ae_ld;
    wire core_io_dmem_s2_xcpt_ae_st;
    wire[33:0] core_io_dmem_s2_gpa;
    wire core_io_dmem_s2_gpa_is_pte;
    wire core_io_dmem_ordered;
    wire core_io_dmem_perf_acquire;
    wire core_io_dmem_perf_release;
    wire core_io_dmem_perf_grant;
    wire core_io_dmem_perf_tlbMiss;
    wire core_io_dmem_perf_blocked;
    wire core_io_dmem_perf_canAcceptStoreThenLoad;
    wire core_io_dmem_perf_canAcceptStoreThenRMW;
    wire core_io_dmem_perf_canAcceptLoadThenLoad;
    wire core_io_dmem_perf_storeBufferEmptyAfterLoad;
    wire core_io_dmem_perf_storeBufferEmptyAfterStore;
    wire core_io_dmem_keep_clock_enabled;
    wire core_io_dmem_clock_enabled;
    wire[3:0] core_io_ptw_ptbr_mode;
    wire[15:0] core_io_ptw_ptbr_asid;
    wire[43:0] core_io_ptw_ptbr_ppn;
    wire[3:0] core_io_ptw_hgatp_mode;
    wire[15:0] core_io_ptw_hgatp_asid;
    wire[43:0] core_io_ptw_hgatp_ppn;
    wire[3:0] core_io_ptw_vsatp_mode;
    wire[15:0] core_io_ptw_vsatp_asid;
    wire[43:0] core_io_ptw_vsatp_ppn;
    wire core_io_ptw_sfence_valid;
    wire core_io_ptw_sfence_bits_rs1;
    wire core_io_ptw_sfence_bits_rs2;
    wire[32:0] core_io_ptw_sfence_bits_addr;
    wire core_io_ptw_sfence_bits_asid;
    wire core_io_ptw_sfence_bits_hv;
    wire core_io_ptw_sfence_bits_hg;
    wire core_io_ptw_status_debug;
    wire core_io_ptw_status_cease;
    wire core_io_ptw_status_wfi;
    wire[31:0] core_io_ptw_status_isa;
    wire[1:0] core_io_ptw_status_dprv;
    wire core_io_ptw_status_dv;
    wire[1:0] core_io_ptw_status_prv;
    wire core_io_ptw_status_v;
    wire core_io_ptw_status_sd;
    wire[22:0] core_io_ptw_status_zero2;
    wire core_io_ptw_status_mpv;
    wire core_io_ptw_status_gva;
    wire core_io_ptw_status_mbe;
    wire core_io_ptw_status_sbe;
    wire[1:0] core_io_ptw_status_sxl;
    wire[1:0] core_io_ptw_status_uxl;
    wire core_io_ptw_status_sd_rv32;
    wire[7:0] core_io_ptw_status_zero1;
    wire core_io_ptw_status_tsr;
    wire core_io_ptw_status_tw;
    wire core_io_ptw_status_tvm;
    wire core_io_ptw_status_mxr;
    wire core_io_ptw_status_sum;
    wire core_io_ptw_status_mprv;
    wire[1:0] core_io_ptw_status_xs;
    wire[1:0] core_io_ptw_status_fs;
    wire[1:0] core_io_ptw_status_mpp;
    wire[1:0] core_io_ptw_status_vs;
    wire core_io_ptw_status_spp;
    wire core_io_ptw_status_mpie;
    wire core_io_ptw_status_ube;
    wire core_io_ptw_status_spie;
    wire core_io_ptw_status_upie;
    wire core_io_ptw_status_mie;
    wire core_io_ptw_status_hie;
    wire core_io_ptw_status_sie;
    wire core_io_ptw_status_uie;
    wire[29:0] core_io_ptw_hstatus_zero6;
    wire[1:0] core_io_ptw_hstatus_vsxl;
    wire[8:0] core_io_ptw_hstatus_zero5;
    wire core_io_ptw_hstatus_vtsr;
    wire core_io_ptw_hstatus_vtw;
    wire core_io_ptw_hstatus_vtvm;
    wire[1:0] core_io_ptw_hstatus_zero3;
    wire[5:0] core_io_ptw_hstatus_vgein;
    wire[1:0] core_io_ptw_hstatus_zero2;
    wire core_io_ptw_hstatus_hu;
    wire core_io_ptw_hstatus_spvp;
    wire core_io_ptw_hstatus_spv;
    wire core_io_ptw_hstatus_gva;
    wire core_io_ptw_hstatus_vsbe;
    wire[4:0] core_io_ptw_hstatus_zero1;
    wire core_io_ptw_gstatus_debug;
    wire core_io_ptw_gstatus_cease;
    wire core_io_ptw_gstatus_wfi;
    wire[31:0] core_io_ptw_gstatus_isa;
    wire[1:0] core_io_ptw_gstatus_dprv;
    wire core_io_ptw_gstatus_dv;
    wire[1:0] core_io_ptw_gstatus_prv;
    wire core_io_ptw_gstatus_v;
    wire core_io_ptw_gstatus_sd;
    wire[22:0] core_io_ptw_gstatus_zero2;
    wire core_io_ptw_gstatus_mpv;
    wire core_io_ptw_gstatus_gva;
    wire core_io_ptw_gstatus_mbe;
    wire core_io_ptw_gstatus_sbe;
    wire[1:0] core_io_ptw_gstatus_sxl;
    wire[1:0] core_io_ptw_gstatus_uxl;
    wire core_io_ptw_gstatus_sd_rv32;
    wire[7:0] core_io_ptw_gstatus_zero1;
    wire core_io_ptw_gstatus_tsr;
    wire core_io_ptw_gstatus_tw;
    wire core_io_ptw_gstatus_tvm;
    wire core_io_ptw_gstatus_mxr;
    wire core_io_ptw_gstatus_sum;
    wire core_io_ptw_gstatus_mprv;
    wire[1:0] core_io_ptw_gstatus_xs;
    wire[1:0] core_io_ptw_gstatus_fs;
    wire[1:0] core_io_ptw_gstatus_mpp;
    wire[1:0] core_io_ptw_gstatus_vs;
    wire core_io_ptw_gstatus_spp;
    wire core_io_ptw_gstatus_mpie;
    wire core_io_ptw_gstatus_ube;
    wire core_io_ptw_gstatus_spie;
    wire core_io_ptw_gstatus_upie;
    wire core_io_ptw_gstatus_mie;
    wire core_io_ptw_gstatus_hie;
    wire core_io_ptw_gstatus_sie;
    wire core_io_ptw_gstatus_uie;
    wire core_io_ptw_pmp_0_cfg_l;
    wire[1:0] core_io_ptw_pmp_0_cfg_res;
    wire[1:0] core_io_ptw_pmp_0_cfg_a;
    wire core_io_ptw_pmp_0_cfg_x;
    wire core_io_ptw_pmp_0_cfg_w;
    wire core_io_ptw_pmp_0_cfg_r;
    wire[29:0] core_io_ptw_pmp_0_addr;
    wire[31:0] core_io_ptw_pmp_0_mask;
    wire core_io_ptw_pmp_1_cfg_l;
    wire[1:0] core_io_ptw_pmp_1_cfg_res;
    wire[1:0] core_io_ptw_pmp_1_cfg_a;
    wire core_io_ptw_pmp_1_cfg_x;
    wire core_io_ptw_pmp_1_cfg_w;
    wire core_io_ptw_pmp_1_cfg_r;
    wire[29:0] core_io_ptw_pmp_1_addr;
    wire[31:0] core_io_ptw_pmp_1_mask;
    wire core_io_ptw_pmp_2_cfg_l;
    wire[1:0] core_io_ptw_pmp_2_cfg_res;
    wire[1:0] core_io_ptw_pmp_2_cfg_a;
    wire core_io_ptw_pmp_2_cfg_x;
    wire core_io_ptw_pmp_2_cfg_w;
    wire core_io_ptw_pmp_2_cfg_r;
    wire[29:0] core_io_ptw_pmp_2_addr;
    wire[31:0] core_io_ptw_pmp_2_mask;
    wire core_io_ptw_pmp_3_cfg_l;
    wire[1:0] core_io_ptw_pmp_3_cfg_res;
    wire[1:0] core_io_ptw_pmp_3_cfg_a;
    wire core_io_ptw_pmp_3_cfg_x;
    wire core_io_ptw_pmp_3_cfg_w;
    wire core_io_ptw_pmp_3_cfg_r;
    wire[29:0] core_io_ptw_pmp_3_addr;
    wire[31:0] core_io_ptw_pmp_3_mask;
    wire core_io_ptw_pmp_4_cfg_l;
    wire[1:0] core_io_ptw_pmp_4_cfg_res;
    wire[1:0] core_io_ptw_pmp_4_cfg_a;
    wire core_io_ptw_pmp_4_cfg_x;
    wire core_io_ptw_pmp_4_cfg_w;
    wire core_io_ptw_pmp_4_cfg_r;
    wire[29:0] core_io_ptw_pmp_4_addr;
    wire[31:0] core_io_ptw_pmp_4_mask;
    wire core_io_ptw_pmp_5_cfg_l;
    wire[1:0] core_io_ptw_pmp_5_cfg_res;
    wire[1:0] core_io_ptw_pmp_5_cfg_a;
    wire core_io_ptw_pmp_5_cfg_x;
    wire core_io_ptw_pmp_5_cfg_w;
    wire core_io_ptw_pmp_5_cfg_r;
    wire[29:0] core_io_ptw_pmp_5_addr;
    wire[31:0] core_io_ptw_pmp_5_mask;
    wire core_io_ptw_pmp_6_cfg_l;
    wire[1:0] core_io_ptw_pmp_6_cfg_res;
    wire[1:0] core_io_ptw_pmp_6_cfg_a;
    wire core_io_ptw_pmp_6_cfg_x;
    wire core_io_ptw_pmp_6_cfg_w;
    wire core_io_ptw_pmp_6_cfg_r;
    wire[29:0] core_io_ptw_pmp_6_addr;
    wire[31:0] core_io_ptw_pmp_6_mask;
    wire core_io_ptw_pmp_7_cfg_l;
    wire[1:0] core_io_ptw_pmp_7_cfg_res;
    wire[1:0] core_io_ptw_pmp_7_cfg_a;
    wire core_io_ptw_pmp_7_cfg_x;
    wire core_io_ptw_pmp_7_cfg_w;
    wire core_io_ptw_pmp_7_cfg_r;
    wire[29:0] core_io_ptw_pmp_7_addr;
    wire[31:0] core_io_ptw_pmp_7_mask;
    wire core_io_ptw_perf_l2miss;
    wire core_io_ptw_perf_l2hit;
    wire core_io_ptw_perf_pte_miss;
    wire core_io_ptw_perf_pte_hit;
    wire core_io_ptw_customCSRs_csrs_0_ren;
    wire core_io_ptw_customCSRs_csrs_0_wen;
    wire[63:0] core_io_ptw_customCSRs_csrs_0_wdata;
    wire[63:0] core_io_ptw_customCSRs_csrs_0_value;
    wire core_io_ptw_customCSRs_csrs_0_stall;
    wire core_io_ptw_customCSRs_csrs_0_set;
    wire[63:0] core_io_ptw_customCSRs_csrs_0_sdata;
    wire core_io_ptw_customCSRs_csrs_1_ren;
    wire core_io_ptw_customCSRs_csrs_1_wen;
    wire[63:0] core_io_ptw_customCSRs_csrs_1_wdata;
    wire[63:0] core_io_ptw_customCSRs_csrs_1_value;
    wire core_io_ptw_customCSRs_csrs_1_stall;
    wire core_io_ptw_customCSRs_csrs_1_set;
    wire[63:0] core_io_ptw_customCSRs_csrs_1_sdata;
    wire core_io_ptw_customCSRs_csrs_2_ren;
    wire core_io_ptw_customCSRs_csrs_2_wen;
    wire[63:0] core_io_ptw_customCSRs_csrs_2_wdata;
    wire[63:0] core_io_ptw_customCSRs_csrs_2_value;
    wire core_io_ptw_customCSRs_csrs_2_stall;
    wire core_io_ptw_customCSRs_csrs_2_set;
    wire[63:0] core_io_ptw_customCSRs_csrs_2_sdata;
    wire core_io_ptw_customCSRs_csrs_3_ren;
    wire core_io_ptw_customCSRs_csrs_3_wen;
    wire[63:0] core_io_ptw_customCSRs_csrs_3_wdata;
    wire[63:0] core_io_ptw_customCSRs_csrs_3_value;
    wire core_io_ptw_customCSRs_csrs_3_stall;
    wire core_io_ptw_customCSRs_csrs_3_set;
    wire[63:0] core_io_ptw_customCSRs_csrs_3_sdata;
    wire core_io_ptw_clock_enabled;
    wire core_io_fpu_hartid;
    wire[63:0] core_io_fpu_time;
    wire[31:0] core_io_fpu_inst;
    wire[63:0] core_io_fpu_fromint_data;
    wire[2:0] core_io_fpu_fcsr_rm;
    wire core_io_fpu_fcsr_flags_valid;
    wire[4:0] core_io_fpu_fcsr_flags_bits;
    wire[63:0] core_io_fpu_toint_data;
    wire core_io_fpu_dmem_resp_val;
    wire[2:0] core_io_fpu_dmem_resp_type;
    wire[4:0] core_io_fpu_dmem_resp_tag;
    wire core_io_fpu_valid;
    wire core_io_fpu_fcsr_rdy;
    wire core_io_fpu_nack_mem;
    wire core_io_fpu_illegal_rm;
    wire core_io_fpu_killx;
    wire core_io_fpu_killm;
    wire core_io_fpu_dec_ldst;
    wire core_io_fpu_dec_wen;
    wire core_io_fpu_dec_ren1;
    wire core_io_fpu_dec_ren2;
    wire core_io_fpu_dec_ren3;
    wire core_io_fpu_dec_swap12;
    wire core_io_fpu_dec_swap23;
    wire[1:0] core_io_fpu_dec_typeTagIn;
    wire[1:0] core_io_fpu_dec_typeTagOut;
    wire core_io_fpu_dec_fromint;
    wire core_io_fpu_dec_toint;
    wire core_io_fpu_dec_fastpipe;
    wire core_io_fpu_dec_fma;
    wire core_io_fpu_dec_div;
    wire core_io_fpu_dec_sqrt;
    wire core_io_fpu_dec_wflags;
    wire core_io_fpu_sboard_set;
    wire core_io_fpu_sboard_clr;
    wire[4:0] core_io_fpu_sboard_clra;
    wire core_io_fpu_keep_clock_enabled;
    wire core_io_rocc_cmd_ready;
    wire core_io_rocc_cmd_valid;
    wire[6:0] core_io_rocc_cmd_bits_inst_funct;
    wire[4:0] core_io_rocc_cmd_bits_inst_rs2;
    wire[4:0] core_io_rocc_cmd_bits_inst_rs1;
    wire core_io_rocc_cmd_bits_inst_xd;
    wire core_io_rocc_cmd_bits_inst_xs1;
    wire core_io_rocc_cmd_bits_inst_xs2;
    wire[4:0] core_io_rocc_cmd_bits_inst_rd;
    wire[6:0] core_io_rocc_cmd_bits_inst_opcode;
    wire[63:0] core_io_rocc_cmd_bits_rs1;
    wire[63:0] core_io_rocc_cmd_bits_rs2;
    wire core_io_rocc_cmd_bits_status_debug;
    wire core_io_rocc_cmd_bits_status_cease;
    wire core_io_rocc_cmd_bits_status_wfi;
    wire[31:0] core_io_rocc_cmd_bits_status_isa;
    wire[1:0] core_io_rocc_cmd_bits_status_dprv;
    wire core_io_rocc_cmd_bits_status_dv;
    wire[1:0] core_io_rocc_cmd_bits_status_prv;
    wire core_io_rocc_cmd_bits_status_v;
    wire core_io_rocc_cmd_bits_status_sd;
    wire[22:0] core_io_rocc_cmd_bits_status_zero2;
    wire core_io_rocc_cmd_bits_status_mpv;
    wire core_io_rocc_cmd_bits_status_gva;
    wire core_io_rocc_cmd_bits_status_mbe;
    wire core_io_rocc_cmd_bits_status_sbe;
    wire[1:0] core_io_rocc_cmd_bits_status_sxl;
    wire[1:0] core_io_rocc_cmd_bits_status_uxl;
    wire core_io_rocc_cmd_bits_status_sd_rv32;
    wire[7:0] core_io_rocc_cmd_bits_status_zero1;
    wire core_io_rocc_cmd_bits_status_tsr;
    wire core_io_rocc_cmd_bits_status_tw;
    wire core_io_rocc_cmd_bits_status_tvm;
    wire core_io_rocc_cmd_bits_status_mxr;
    wire core_io_rocc_cmd_bits_status_sum;
    wire core_io_rocc_cmd_bits_status_mprv;
    wire[1:0] core_io_rocc_cmd_bits_status_xs;
    wire[1:0] core_io_rocc_cmd_bits_status_fs;
    wire[1:0] core_io_rocc_cmd_bits_status_mpp;
    wire[1:0] core_io_rocc_cmd_bits_status_vs;
    wire core_io_rocc_cmd_bits_status_spp;
    wire core_io_rocc_cmd_bits_status_mpie;
    wire core_io_rocc_cmd_bits_status_ube;
    wire core_io_rocc_cmd_bits_status_spie;
    wire core_io_rocc_cmd_bits_status_upie;
    wire core_io_rocc_cmd_bits_status_mie;
    wire core_io_rocc_cmd_bits_status_hie;
    wire core_io_rocc_cmd_bits_status_sie;
    wire core_io_rocc_cmd_bits_status_uie;
    wire core_io_rocc_resp_ready;
    wire core_io_rocc_resp_valid;
    wire[4:0] core_io_rocc_resp_bits_rd;
    wire[63:0] core_io_rocc_resp_bits_data;
    wire core_io_rocc_mem_req_ready;
    wire core_io_rocc_mem_req_valid;
    wire[33:0] core_io_rocc_mem_req_bits_addr;
    wire[5:0] core_io_rocc_mem_req_bits_tag;
    wire[4:0] core_io_rocc_mem_req_bits_cmd;
    wire[1:0] core_io_rocc_mem_req_bits_size;
    wire core_io_rocc_mem_req_bits_signed;
    wire[1:0] core_io_rocc_mem_req_bits_dprv;
    wire core_io_rocc_mem_req_bits_dv;
    wire core_io_rocc_mem_req_bits_phys;
    wire core_io_rocc_mem_req_bits_no_alloc;
    wire core_io_rocc_mem_req_bits_no_xcpt;
    wire[63:0] core_io_rocc_mem_req_bits_data;
    wire[7:0] core_io_rocc_mem_req_bits_mask;
    wire core_io_rocc_mem_s1_kill;
    wire[63:0] core_io_rocc_mem_s1_data_data;
    wire[7:0] core_io_rocc_mem_s1_data_mask;
    wire core_io_rocc_mem_s2_nack;
    wire core_io_rocc_mem_s2_nack_cause_raw;
    wire core_io_rocc_mem_s2_kill;
    wire core_io_rocc_mem_s2_uncached;
    wire[31:0] core_io_rocc_mem_s2_paddr;
    wire core_io_rocc_mem_resp_valid;
    wire[33:0] core_io_rocc_mem_resp_bits_addr;
    wire[5:0] core_io_rocc_mem_resp_bits_tag;
    wire[4:0] core_io_rocc_mem_resp_bits_cmd;
    wire[1:0] core_io_rocc_mem_resp_bits_size;
    wire core_io_rocc_mem_resp_bits_signed;
    wire[1:0] core_io_rocc_mem_resp_bits_dprv;
    wire core_io_rocc_mem_resp_bits_dv;
    wire[63:0] core_io_rocc_mem_resp_bits_data;
    wire[7:0] core_io_rocc_mem_resp_bits_mask;
    wire core_io_rocc_mem_resp_bits_replay;
    wire core_io_rocc_mem_resp_bits_has_data;
    wire[63:0] core_io_rocc_mem_resp_bits_data_word_bypass;
    wire[63:0] core_io_rocc_mem_resp_bits_data_raw;
    wire[63:0] core_io_rocc_mem_resp_bits_store_data;
    wire core_io_rocc_mem_replay_next;
    wire core_io_rocc_mem_s2_xcpt_ma_ld;
    wire core_io_rocc_mem_s2_xcpt_ma_st;
    wire core_io_rocc_mem_s2_xcpt_pf_ld;
    wire core_io_rocc_mem_s2_xcpt_pf_st;
    wire core_io_rocc_mem_s2_xcpt_gf_ld;
    wire core_io_rocc_mem_s2_xcpt_gf_st;
    wire core_io_rocc_mem_s2_xcpt_ae_ld;
    wire core_io_rocc_mem_s2_xcpt_ae_st;
    wire[33:0] core_io_rocc_mem_s2_gpa;
    wire core_io_rocc_mem_s2_gpa_is_pte;
    wire core_io_rocc_mem_ordered;
    wire core_io_rocc_mem_perf_acquire;
    wire core_io_rocc_mem_perf_release;
    wire core_io_rocc_mem_perf_grant;
    wire core_io_rocc_mem_perf_tlbMiss;
    wire core_io_rocc_mem_perf_blocked;
    wire core_io_rocc_mem_perf_canAcceptStoreThenLoad;
    wire core_io_rocc_mem_perf_canAcceptStoreThenRMW;
    wire core_io_rocc_mem_perf_canAcceptLoadThenLoad;
    wire core_io_rocc_mem_perf_storeBufferEmptyAfterLoad;
    wire core_io_rocc_mem_perf_storeBufferEmptyAfterStore;
    wire core_io_rocc_mem_keep_clock_enabled;
    wire core_io_rocc_mem_clock_enabled;
    wire core_io_rocc_busy;
    wire core_io_rocc_interrupt;
    wire core_io_rocc_exception;
    wire core_io_trace_insns_0_valid;
    wire[33:0] core_io_trace_insns_0_iaddr;
    wire[31:0] core_io_trace_insns_0_insn;
    wire[2:0] core_io_trace_insns_0_priv;
    wire core_io_trace_insns_0_exception;
    wire core_io_trace_insns_0_interrupt;
    wire[63:0] core_io_trace_insns_0_cause;
    wire[33:0] core_io_trace_insns_0_tval;
    wire[63:0] core_io_trace_time;
    wire core_io_bpwatch_0_valid_0;
    wire core_io_bpwatch_0_rvalid_0;
    wire core_io_bpwatch_0_wvalid_0;
    wire core_io_bpwatch_0_ivalid_0;
    wire[2:0] core_io_bpwatch_0_action;
    wire core_io_cease;
    wire core_io_wfi;
    wire core_io_traceStall;

    wire[31:0] core__csr_io_time_31to0 ; 
    wire core__GEN ; 
    wire[2:0] core__GEN_0 ; 
    wire[11:0] core__wb_reg_inst_31to20 ; 
    wire[39:0] core__GEN_1 ; 
    wire[33:0] core__GEN_2 ; 
    wire core__GEN_3 ; 
    wire[31:0] core__GEN_4 ; 
    wire core__GEN_5 ; 
    wire[4:0] core__GEN_6 ; 
    wire core__GEN_7 ; 
    wire core__GEN_8 ; 
    wire core__GEN_9 ; 
    wire[63:0] core_ll_wdata ; 
    wire[32:0] core__mem_reg_wdata_32to0 ; 
    wire[32:0] core__ibuf_io_pc_32to0 ; 
    wire[63:0] core__io_ptw_customCSRs_csrs_0_value_output ; 
    wire[4:0] core__GEN_10 ; 
    wire[4:0] core__GEN_11 ; 
    wire core__GEN_12 ; 
    wire[4:0] core_id_waddr ; 
    wire[4:0] core_id_raddr2 ; 
    wire[4:0] core_id_raddr3 ; 
    wire core__div_io_req_ready ; 
    wire core__div_io_resp_valid ; 
    wire[4:0] core__div_io_resp_bits_tag ; 
    wire[63:0] core__alu_io_out ; 
    wire[63:0] core__alu_io_adder_out ; 
    wire core__alu_io_cmp_out ; 
    wire core__bpu_io_xcpt_if ; 
    wire core__bpu_io_xcpt_ld ; 
    wire core__bpu_io_xcpt_st ; 
    wire core__bpu_io_debug_if ; 
    wire core__bpu_io_debug_ld ; 
    wire core__bpu_io_debug_st ; 
    wire core__bpu_io_bpwatch_0_rvalid_0 ; 
    wire core__bpu_io_bpwatch_0_wvalid_0 ; 
    wire core__bpu_io_bpwatch_0_ivalid_0 ; 
    wire[63:0] core__csr_io_rw_rdata ; 
    wire core__csr_io_decode_0_fp_illegal ; 
    wire core__csr_io_decode_0_fp_csr ; 
    wire core__csr_io_decode_0_rocc_illegal ; 
    wire core__csr_io_decode_0_read_illegal ; 
    wire core__csr_io_decode_0_write_illegal ; 
    wire core__csr_io_decode_0_write_flush ; 
    wire core__csr_io_decode_0_system_illegal ; 
    wire core__csr_io_decode_0_virtual_access_illegal ; 
    wire core__csr_io_decode_0_virtual_system_illegal ; 
    wire core__csr_io_csr_stall ; 
    wire core__csr_io_rw_stall ; 
    wire core__csr_io_eret ; 
    wire core__csr_io_singleStep ; 
    wire core__csr_io_status_debug ; 
    wire core__csr_io_status_cease ; 
    wire core__csr_io_status_wfi ; 
    wire[31:0] core__csr_io_status_isa ; 
    wire[1:0] core__csr_io_status_dprv ; 
    wire core__csr_io_status_dv ; 
    wire[1:0] core__csr_io_status_prv ; 
    wire core__csr_io_status_v ; 
    wire core__csr_io_status_sd ; 
    wire[22:0] core__csr_io_status_zero2 ; 
    wire core__csr_io_status_mpv ; 
    wire core__csr_io_status_gva ; 
    wire core__csr_io_status_mbe ; 
    wire core__csr_io_status_sbe ; 
    wire[1:0] core__csr_io_status_sxl ; 
    wire[1:0] core__csr_io_status_uxl ; 
    wire core__csr_io_status_sd_rv32 ; 
    wire[7:0] core__csr_io_status_zero1 ; 
    wire core__csr_io_status_tsr ; 
    wire core__csr_io_status_tw ; 
    wire core__csr_io_status_tvm ; 
    wire core__csr_io_status_mxr ; 
    wire core__csr_io_status_sum ; 
    wire core__csr_io_status_mprv ; 
    wire[1:0] core__csr_io_status_xs ; 
    wire[1:0] core__csr_io_status_fs ; 
    wire[1:0] core__csr_io_status_mpp ; 
    wire[1:0] core__csr_io_status_vs ; 
    wire core__csr_io_status_spp ; 
    wire core__csr_io_status_mpie ; 
    wire core__csr_io_status_ube ; 
    wire core__csr_io_status_spie ; 
    wire core__csr_io_status_upie ; 
    wire core__csr_io_status_mie ; 
    wire core__csr_io_status_hie ; 
    wire core__csr_io_status_sie ; 
    wire core__csr_io_status_uie ; 
    wire core__csr_io_hstatus_spvp ; 
    wire[33:0] core__csr_io_evec ; 
    wire[63:0] core__csr_io_time ; 
    wire core__csr_io_interrupt ; 
    wire[63:0] core__csr_io_interrupt_cause ; 
    wire[3:0] core__csr_io_bp_0_control_ttype ; 
    wire core__csr_io_bp_0_control_dmode ; 
    wire[5:0] core__csr_io_bp_0_control_maskmax ; 
    wire[39:0] core__csr_io_bp_0_control_reserved ; 
    wire core__csr_io_bp_0_control_action ; 
    wire core__csr_io_bp_0_control_chain ; 
    wire[1:0] core__csr_io_bp_0_control_zero ; 
    wire[1:0] core__csr_io_bp_0_control_tmatch ; 
    wire core__csr_io_bp_0_control_m ; 
    wire core__csr_io_bp_0_control_h ; 
    wire core__csr_io_bp_0_control_s ; 
    wire core__csr_io_bp_0_control_u ; 
    wire core__csr_io_bp_0_control_x ; 
    wire core__csr_io_bp_0_control_w ; 
    wire core__csr_io_bp_0_control_r ; 
    wire[32:0] core__csr_io_bp_0_address ; 
    wire core__csr_io_bp_0_textra_mselect ; 
    wire[47:0] core__csr_io_bp_0_textra_pad2 ; 
    wire core__csr_io_bp_0_textra_pad1 ; 
    wire core__csr_io_bp_0_textra_sselect ; 
    wire core__csr_io_inhibit_cycle ; 
    wire core__csr_io_trace_0_valid ; 
    wire[33:0] core__csr_io_trace_0_iaddr ; 
    wire[31:0] core__csr_io_trace_0_insn ; 
    wire[2:0] core__csr_io_trace_0_priv ; 
    wire core__csr_io_trace_0_exception ; 
    wire[63:0] core__rf_ext_R0_data ; 
    wire[63:0] core__rf_ext_R1_data ; 
    wire[33:0] core__ibuf_io_pc ; 
    wire[1:0] core__ibuf_io_btb_resp_cfiType ; 
    wire core__ibuf_io_btb_resp_taken ; 
    wire[1:0] core__ibuf_io_btb_resp_mask ; 
    wire core__ibuf_io_btb_resp_bridx ; 
    wire[32:0] core__ibuf_io_btb_resp_target ; 
    wire core__ibuf_io_btb_resp_entry ; 
    wire[7:0] core__ibuf_io_btb_resp_bht_history ; 
    wire core__ibuf_io_btb_resp_bht_value ; 
    wire core__ibuf_io_inst_0_valid ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_pf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_gf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt0_ae_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_pf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_gf_inst ; 
    wire core__ibuf_io_inst_0_bits_xcpt1_ae_inst ; 
    wire core__ibuf_io_inst_0_bits_replay ; 
    wire core__ibuf_io_inst_0_bits_rvc ; 
    wire[31:0] core__ibuf_io_inst_0_bits_inst_bits ; 
    wire[4:0] core__ibuf_io_inst_0_bits_inst_rs1 ; 
    wire[31:0] core__ibuf_io_inst_0_bits_raw ; 
    wire[63:0] core_dcache_bypass_data = core_io_dmem_resp_bits_data_word_bypass ; 
    wire core_coreMonitorBundle_clock = core_clock ; 
    wire core_coreMonitorBundle_reset = core_reset ; 
    wire core_xrfWriteBundle_clock = core_clock ; 
    wire core_xrfWriteBundle_reset = core_reset ; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_lo =2'h0; 
    wire core__hits_WIRE_0 =1'h0; 
    wire core__hits_WIRE_1 =1'h0; 
    wire core__hits_WIRE_2 =1'h0; 
    wire core__hits_WIRE_3 =1'h0; 
    wire core__hits_WIRE_4 =1'h0; 
    wire core__hits_WIRE_5 =1'h0; 
    wire core__hits_WIRE_6 =1'h0; 
    wire core__hits_WIRE_7 =1'h0; 
    wire core__hits_WIRE_8 =1'h0; 
    wire core__hits_WIRE_9 =1'h0; 
    wire core__hits_WIRE_10 =1'h0; 
    wire core__hits_WIRE_1_0 =1'h0; 
    wire core__hits_WIRE_1_1 =1'h0; 
    wire core__hits_WIRE_1_2 =1'h0; 
    wire core__hits_WIRE_1_3 =1'h0; 
    wire core__hits_WIRE_1_4 =1'h0; 
    wire core__hits_WIRE_1_5 =1'h0; 
    wire core__hits_WIRE_1_6 =1'h0; 
    wire core__hits_WIRE_1_7 =1'h0; 
    wire core__hits_WIRE_1_8 =1'h0; 
    wire core__hits_WIRE_1_9 =1'h0; 
    wire core__hits_WIRE_2_0 =1'h0; 
    wire core__hits_WIRE_2_1 =1'h0; 
    wire core__hits_WIRE_2_2 =1'h0; 
    wire core__hits_WIRE_2_3 =1'h0; 
    wire core__hits_WIRE_2_4 =1'h0; 
    wire core__hits_WIRE_2_5 =1'h0; 
    wire core_id_npc_b0 =1'h0; 
    wire core_id_rocc_busy =1'h0; 
    wire core_ex_sfence =1'h0; 
    wire core_mem_br_target_b0 =1'h0; 
    wire core_mem_br_target_b0_1 =1'h0; 
    wire core_coreMonitorBundle_wrenf =1'h0; 
    wire core_xrfWriteBundle_excpt =1'h0; 
    wire core_xrfWriteBundle_valid =1'h0; 
    wire core_xrfWriteBundle_wrenf =1'h0; 
    wire core_clock_en =1'h1; 
    reg core_clock_en_reg ; 
    reg core_long_latency_stall ; 
    reg core_id_reg_pause ; 
    reg core_imem_might_request_reg ; 
    wire core_hits_0 = core__hits_WIRE_0 ; 
    wire core_hits_1 = core__hits_WIRE_1 ; 
    wire core_hits_2 = core__hits_WIRE_2 ; 
    wire core_hits_3 = core__hits_WIRE_3 ; 
    wire core_hits_4 = core__hits_WIRE_4 ; 
    wire core_hits_5 = core__hits_WIRE_5 ; 
    wire core_hits_6 = core__hits_WIRE_6 ; 
    wire core_hits_7 = core__hits_WIRE_7 ; 
    wire core_hits_8 = core__hits_WIRE_8 ; 
    wire core_hits_9 = core__hits_WIRE_9 ; 
    wire core_hits_10 = core__hits_WIRE_10 ; 
    wire core_hits_1_0 = core__hits_WIRE_1_0 ; 
    wire core_hits_1_1 = core__hits_WIRE_1_1 ; 
    wire core_hits_1_2 = core__hits_WIRE_1_2 ; 
    wire core_hits_1_3 = core__hits_WIRE_1_3 ; 
    wire core_hits_1_4 = core__hits_WIRE_1_4 ; 
    wire core_hits_1_5 = core__hits_WIRE_1_5 ; 
    wire core_hits_1_6 = core__hits_WIRE_1_6 ; 
    wire core_hits_1_7 = core__hits_WIRE_1_7 ; 
    wire core_hits_1_8 = core__hits_WIRE_1_8 ; 
    wire core_hits_1_9 = core__hits_WIRE_1_9 ; 
    wire core_hits_2_0 = core__hits_WIRE_2_0 ; 
    wire core_hits_2_1 = core__hits_WIRE_2_1 ; 
    wire core_hits_2_2 = core__hits_WIRE_2_2 ; 
    wire core_hits_2_3 = core__hits_WIRE_2_3 ; 
    wire core_hits_2_4 = core__hits_WIRE_2_4 ; 
    wire core_hits_2_5 = core__hits_WIRE_2_5 ; 
    reg core_ex_ctrl_legal ; 
    reg core_ex_ctrl_fp ; 
    reg core_ex_ctrl_rocc ; 
    reg core_ex_ctrl_branch ; 
    reg core_ex_ctrl_jal ; 
    reg core_ex_ctrl_jalr ; 
    reg core_ex_ctrl_rxs2 ; 
    reg core_ex_ctrl_rxs1 ; reg[1:0] core_ex_ctrl_sel_alu2 ; reg[1:0] core_ex_ctrl_sel_alu1 ; reg[2:0] core_ex_ctrl_sel_imm ; 
    reg core_ex_ctrl_alu_dw ; reg[3:0] core_ex_ctrl_alu_fn ; 
    reg core_ex_ctrl_mem ; reg[4:0] core_ex_ctrl_mem_cmd ; 
    reg core_ex_ctrl_rfs1 ; 
    reg core_ex_ctrl_rfs2 ; 
    reg core_ex_ctrl_rfs3 ; 
    reg core_ex_ctrl_wfd ; 
    reg core_ex_ctrl_mul ; 
    reg core_ex_ctrl_div ; 
    reg core_ex_ctrl_wxd ; reg[2:0] core_ex_ctrl_csr ; 
    reg core_ex_ctrl_fence_i ; 
    reg core_ex_ctrl_fence ; 
    reg core_ex_ctrl_amo ; 
    reg core_ex_ctrl_dp ; 
    reg core_mem_ctrl_legal ; 
    reg core_mem_ctrl_fp ; 
    reg core_mem_ctrl_rocc ; 
    reg core_mem_ctrl_branch ; 
    reg core_mem_ctrl_jal ; 
    reg core_mem_ctrl_jalr ; 
    reg core_mem_ctrl_rxs2 ; 
    reg core_mem_ctrl_rxs1 ; reg[1:0] core_mem_ctrl_sel_alu2 ; reg[1:0] core_mem_ctrl_sel_alu1 ; reg[2:0] core_mem_ctrl_sel_imm ; 
    reg core_mem_ctrl_alu_dw ; reg[3:0] core_mem_ctrl_alu_fn ; 
    reg core_mem_ctrl_mem ; reg[4:0] core_mem_ctrl_mem_cmd ; 
    reg core_mem_ctrl_rfs1 ; 
    reg core_mem_ctrl_rfs2 ; 
    reg core_mem_ctrl_rfs3 ; 
    reg core_mem_ctrl_wfd ; 
    reg core_mem_ctrl_mul ; 
    reg core_mem_ctrl_div ; 
    reg core_mem_ctrl_wxd ; reg[2:0] core_mem_ctrl_csr ; 
    reg core_mem_ctrl_fence_i ; 
    reg core_mem_ctrl_fence ; 
    reg core_mem_ctrl_amo ; 
    reg core_mem_ctrl_dp ; 
    reg core_wb_ctrl_legal ; 
    reg core_wb_ctrl_fp ; 
    reg core_wb_ctrl_rocc ; 
    reg core_wb_ctrl_branch ; 
    reg core_wb_ctrl_jal ; 
    reg core_wb_ctrl_jalr ; 
    reg core_wb_ctrl_rxs2 ; 
    reg core_wb_ctrl_rxs1 ; reg[1:0] core_wb_ctrl_sel_alu2 ; reg[1:0] core_wb_ctrl_sel_alu1 ; reg[2:0] core_wb_ctrl_sel_imm ; 
    reg core_wb_ctrl_alu_dw ; reg[3:0] core_wb_ctrl_alu_fn ; 
    reg core_wb_ctrl_mem ; reg[4:0] core_wb_ctrl_mem_cmd ; 
    reg core_wb_ctrl_rfs1 ; 
    reg core_wb_ctrl_rfs2 ; 
    reg core_wb_ctrl_rfs3 ; 
    reg core_wb_ctrl_wfd ; 
    reg core_wb_ctrl_mul ; 
    reg core_wb_ctrl_div ; 
    reg core_wb_ctrl_wxd ; reg[2:0] core_wb_ctrl_csr ; 
    reg core_wb_ctrl_fence_i ; 
    reg core_wb_ctrl_fence ; 
    reg core_wb_ctrl_amo ; 
    reg core_wb_ctrl_dp ; 
    reg core_ex_reg_xcpt_interrupt ; 
    reg core_ex_reg_valid ; 
    reg core_ex_reg_rvc ; reg[1:0] core_ex_reg_btb_resp_cfiType ; 
    reg core_ex_reg_btb_resp_taken ; reg[1:0] core_ex_reg_btb_resp_mask ; 
    reg core_ex_reg_btb_resp_bridx ; reg[32:0] core_ex_reg_btb_resp_target ; 
    reg core_ex_reg_btb_resp_entry ; reg[7:0] core_ex_reg_btb_resp_bht_history ; 
    reg core_ex_reg_btb_resp_bht_value ; 
    reg core_ex_reg_xcpt ; 
    reg core_ex_reg_flush_pipe ; 
    reg core_ex_reg_load_use ; reg[63:0] core_ex_reg_cause ; 
    reg core_ex_reg_replay ; reg[33:0] core_ex_reg_pc ; reg[1:0] core_ex_reg_mem_size ; 
    reg core_ex_reg_hls ; reg[31:0] core_ex_reg_inst ; reg[31:0] core_ex_reg_raw_inst ; 
    reg core_ex_reg_wphit_0 ; 
    reg core_mem_reg_xcpt_interrupt ; 
    reg core_mem_reg_valid ; 
    reg core_mem_reg_rvc ; reg[1:0] core_mem_reg_btb_resp_cfiType ; 
    reg core_mem_reg_btb_resp_taken ; reg[1:0] core_mem_reg_btb_resp_mask ; 
    reg core_mem_reg_btb_resp_bridx ; reg[32:0] core_mem_reg_btb_resp_target ; 
    reg core_mem_reg_btb_resp_entry ; reg[7:0] core_mem_reg_btb_resp_bht_history ; 
    reg core_mem_reg_btb_resp_bht_value ; 
    reg core_mem_reg_xcpt ; 
    reg core_mem_reg_replay ; 
    reg core_mem_reg_flush_pipe ; reg[63:0] core_mem_reg_cause ; 
    reg core_mem_reg_slow_bypass ; 
    reg core_mem_reg_load ; 
    reg core_mem_reg_store ; 
    reg core_mem_reg_sfence ; reg[33:0] core_mem_reg_pc ; reg[31:0] core_mem_reg_inst ; reg[1:0] core_mem_reg_mem_size ; 
    reg core_mem_reg_hls_or_dv ; reg[31:0] core_mem_reg_raw_inst ; reg[63:0] core_mem_reg_wdata ; reg[63:0] core_mem_reg_rs2 ; 
    reg core_mem_br_taken ; 
    reg core_mem_reg_wphit_0 ; 
    reg core_wb_reg_valid ; 
    reg core_wb_reg_xcpt ; 
    reg core_wb_reg_replay ; 
    reg core_wb_reg_flush_pipe ; reg[63:0] core_wb_reg_cause ; 
    reg core_wb_reg_sfence ; reg[33:0] core_wb_reg_pc ; reg[1:0] core_wb_reg_mem_size ; 
    reg core_wb_reg_hls_or_dv ; 
    reg core_wb_reg_hfence_v ; 
    wire core__io_imem_sfence_bits_hv_output = core_wb_reg_hfence_v ; 
    reg core_wb_reg_hfence_g ; 
    wire core__io_imem_sfence_bits_hg_output = core_wb_reg_hfence_g ; reg[31:0] core_wb_reg_inst ; 
    wire[31:0] core__io_rocc_cmd_bits_inst_WIRE_1 = core_wb_reg_inst ; reg[31:0] core_wb_reg_raw_inst ; reg[63:0] core_wb_reg_wdata ; reg[63:0] core_wb_reg_rs2 ; 
    reg core_wb_reg_wphit_0 ; 
    wire core_take_pc_mem ; 
    wire core_take_pc_wb ; 
    wire core_take_pc_mem_wb = core_take_pc_wb | core_take_pc_mem ;  
    wire core_ibuf_clock;
    wire core_ibuf_reset;
    wire core_ibuf_io_imem_ready;
    wire core_ibuf_io_imem_valid;
    wire[1:0] core_ibuf_io_imem_bits_btb_cfiType;
    wire core_ibuf_io_imem_bits_btb_taken;
    wire[1:0] core_ibuf_io_imem_bits_btb_mask;
    wire core_ibuf_io_imem_bits_btb_bridx;
    wire[32:0] core_ibuf_io_imem_bits_btb_target;
    wire core_ibuf_io_imem_bits_btb_entry;
    wire[7:0] core_ibuf_io_imem_bits_btb_bht_history;
    wire core_ibuf_io_imem_bits_btb_bht_value;
    wire[33:0] core_ibuf_io_imem_bits_pc;
    wire[31:0] core_ibuf_io_imem_bits_data;
    wire[1:0] core_ibuf_io_imem_bits_mask;
    wire core_ibuf_io_imem_bits_xcpt_pf_inst;
    wire core_ibuf_io_imem_bits_xcpt_gf_inst;
    wire core_ibuf_io_imem_bits_xcpt_ae_inst;
    wire core_ibuf_io_imem_bits_replay;
    wire core_ibuf_io_kill;
    wire[33:0] core_ibuf_io_pc;
    wire[1:0] core_ibuf_io_btb_resp_cfiType;
    wire core_ibuf_io_btb_resp_taken;
    wire[1:0] core_ibuf_io_btb_resp_mask;
    wire core_ibuf_io_btb_resp_bridx;
    wire[32:0] core_ibuf_io_btb_resp_target;
    wire core_ibuf_io_btb_resp_entry;
    wire[7:0] core_ibuf_io_btb_resp_bht_history;
    wire core_ibuf_io_btb_resp_bht_value;
    wire core_ibuf_io_inst_0_ready;
    wire core_ibuf_io_inst_0_valid;
    wire core_ibuf_io_inst_0_bits_xcpt0_pf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt0_gf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt0_ae_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_pf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_gf_inst;
    wire core_ibuf_io_inst_0_bits_xcpt1_ae_inst;
    wire core_ibuf_io_inst_0_bits_replay;
    wire core_ibuf_io_inst_0_bits_rvc;
    wire[31:0] core_ibuf_io_inst_0_bits_inst_bits;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rd;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs1;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs2;
    wire[4:0] core_ibuf_io_inst_0_bits_inst_rs3;
    wire[31:0] core_ibuf_io_inst_0_bits_raw;

    wire core_ibuf__exp_io_rvc ; 
    reg core_ibuf_nBufValid ; reg[1:0] core_ibuf_buf_btb_cfiType ; 
    reg core_ibuf_buf_btb_taken ; reg[1:0] core_ibuf_buf_btb_mask ; 
    reg core_ibuf_buf_btb_bridx ; reg[32:0] core_ibuf_buf_btb_target ; 
    reg core_ibuf_buf_btb_entry ; reg[7:0] core_ibuf_buf_btb_bht_history ; 
    reg core_ibuf_buf_btb_bht_value ; reg[33:0] core_ibuf_buf_pc ; reg[31:0] core_ibuf_buf_data ; reg[1:0] core_ibuf_buf_mask ; 
    reg core_ibuf_buf_xcpt_pf_inst ; 
    reg core_ibuf_buf_xcpt_gf_inst ; 
    reg core_ibuf_buf_xcpt_ae_inst ; 
    reg core_ibuf_buf_replay ; reg[1:0] core_ibuf_ibufBTBResp_cfiType ; 
    reg core_ibuf_ibufBTBResp_taken ; reg[1:0] core_ibuf_ibufBTBResp_mask ; 
    reg core_ibuf_ibufBTBResp_bridx ; reg[32:0] core_ibuf_ibufBTBResp_target ; 
    reg core_ibuf_ibufBTBResp_entry ; reg[7:0] core_ibuf_ibufBTBResp_bht_history ; 
    reg core_ibuf_ibufBTBResp_bht_value ; 
    wire core_ibuf_pcWordBits = core_ibuf_io_imem_bits_pc [1]; 
    wire[2:0] core_ibuf__GEN ={1'h0, core_ibuf_io_imem_bits_btb_taken  ? {1'h0, core_ibuf_io_imem_bits_btb_bridx }+2'h1:2'h2}-{2'h0, core_ibuf_pcWordBits }; 
    wire[1:0] core_ibuf_nIC = core_ibuf__GEN [1:0]; 
    wire[1:0] core_ibuf_nReady ; 
    wire[2:0] core_ibuf__GEN_0 ={1'h0, core_ibuf_nReady }-{2'h0, core_ibuf_nBufValid }; 
    wire[1:0] core_ibuf_nICReady = core_ibuf__GEN_0 [1:0]; 
    wire[2:0] core_ibuf__GEN_1 ={1'h0, core_ibuf_io_imem_valid  ?  core_ibuf_nIC :2'h0}+{2'h0, core_ibuf_nBufValid }; 
    wire[1:0] core_ibuf_nValid = core_ibuf__GEN_1 [1:0]; 
    wire[2:0] core_ibuf__GEN_2 ={1'h0, core_ibuf_nIC }-{1'h0, core_ibuf_nICReady }; 
    wire[2:0] core_ibuf__GEN_3 ={2'h0, core_ibuf_nBufValid }-{1'h0, core_ibuf_nReady }; 
    wire[1:0] core_ibuf__GEN_4 = core_ibuf_nReady >={1'h0, core_ibuf_nBufValid }| core_ibuf_nBufValid ==1'h0 ? 2'h0: core_ibuf__GEN_3 [1:0]; 
    wire[2:0] core_ibuf__GEN_5 ={1'h0, core_ibuf_nIC }-{1'h0, core_ibuf_nICReady }; 
    wire core_ibuf__GEN_6 = core_ibuf_io_imem_valid & core_ibuf_nReady >={1'h0, core_ibuf_nBufValid }& core_ibuf_nICReady < core_ibuf_nIC &2'h1>= core_ibuf__GEN_5 [1:0]; 
    wire[2:0] core_ibuf__GEN_7 ={2'h0, core_ibuf_pcWordBits }+{1'h0, core_ibuf_nICReady }; 
    wire[1:0] core_ibuf_shamt = core_ibuf__GEN_7 [1:0]; 
    wire[2:0] core_ibuf__GEN_8 ={1'h0, core_ibuf_nIC }-{1'h0, core_ibuf_nICReady }; 
    wire[1:0] core_ibuf__GEN_9 = core_ibuf__GEN_8 [1:0]; 
    wire[63:0] core_ibuf_buf_data_data ={{ core_ibuf_io_imem_bits_data [31:16], core_ibuf_io_imem_bits_data [31:16]}, core_ibuf_io_imem_bits_data }; 
    wire[63:0] core_ibuf__GEN_10 = core_ibuf_buf_data_data >>{ core_ibuf_shamt ,4'h0}; 
    wire[31:0] core_ibuf__GEN_11 ={16'h0, core_ibuf__GEN_10 [15:0]}; 
    wire[34:0] core_ibuf__GEN_12 ={1'h0, core_ibuf_io_imem_bits_pc }+{32'h0,{ core_ibuf_nICReady ,1'h0}}; 
    wire[33:0] core_ibuf__GEN_13 = core_ibuf_io_imem_bits_pc &34'h3FFFFFFFC| core_ibuf__GEN_12 [33:0]&34'h3; 
    wire[2:0] core_ibuf__GEN_14 ={2'h0, core_ibuf_nBufValid }+3'h2; 
    wire[2:0] core_ibuf__GEN_15 ={1'h0, core_ibuf__GEN_14 [1:0]}-{2'h0, core_ibuf_pcWordBits }; 
    wire[1:0] core_ibuf_icShiftAmt = core_ibuf__GEN_15 [1:0]; 
    wire[63:0] core_ibuf__GEN_16 ={ core_ibuf_io_imem_bits_data ,{ core_ibuf_io_imem_bits_data [15:0], core_ibuf_io_imem_bits_data [15:0]}}; 
    wire[31:0] core_ibuf__GEN_17 ={ core_ibuf__GEN_16 [63:48], core_ibuf__GEN_16 [63:48]}; 
    wire[127:0] core_ibuf_icData_data ={{ core_ibuf__GEN_17 , core_ibuf__GEN_17 }, core_ibuf__GEN_16 }; 
    wire[190:0] core_ibuf__GEN_18 ={63'h0, core_ibuf_icData_data }<<{ core_ibuf_icShiftAmt ,4'h0}; 
    wire[31:0] core_ibuf_icData = core_ibuf__GEN_18 [95:64]; 
    wire[62:0] core_ibuf__GEN_19 =63'hFFFFFFFF<<{ core_ibuf_nBufValid ,4'h0}; 
    wire[31:0] core_ibuf_icMask = core_ibuf__GEN_19 [31:0]; 
    wire[31:0] core_ibuf_inst = core_ibuf_icData & core_ibuf_icMask | core_ibuf_buf_data &~ core_ibuf_icMask ; 
    wire[4:0] core_ibuf__GEN_20 ={1'h0,4'h1<< core_ibuf_nValid }-5'h1; 
    wire[3:0] core_ibuf__GEN_21 = core_ibuf__GEN_20 [3:0]; 
    wire[1:0] core_ibuf_valid = core_ibuf__GEN_21 [1:0]; 
    wire[2:0] core_ibuf__GEN_22 ={1'h0,2'h1<< core_ibuf_nBufValid }-3'h1; 
    wire[1:0] core_ibuf_bufMask = core_ibuf__GEN_22 [1:0]; 
    wire core_ibuf_xcpt_0_pf_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_pf_inst : core_ibuf_io_imem_bits_xcpt_pf_inst ; 
    wire core_ibuf_xcpt_0_gf_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_gf_inst : core_ibuf_io_imem_bits_xcpt_gf_inst ; 
    wire core_ibuf_xcpt_0_ae_inst = core_ibuf_bufMask [0] ?  core_ibuf_buf_xcpt_ae_inst : core_ibuf_io_imem_bits_xcpt_ae_inst ; 
    wire core_ibuf_xcpt_1_pf_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_pf_inst : core_ibuf_io_imem_bits_xcpt_pf_inst ; 
    wire core_ibuf_xcpt_1_gf_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_gf_inst : core_ibuf_io_imem_bits_xcpt_gf_inst ; 
    wire core_ibuf_xcpt_1_ae_inst = core_ibuf_bufMask [1] ?  core_ibuf_buf_xcpt_ae_inst : core_ibuf_io_imem_bits_xcpt_ae_inst ; 
    wire[1:0] core_ibuf_buf_replay_0 = core_ibuf_buf_replay  ?  core_ibuf_bufMask :2'h0; 
    wire[1:0] core_ibuf_ic_replay = core_ibuf_buf_replay_0 |( core_ibuf_io_imem_bits_replay  ?  core_ibuf_valid &~ core_ibuf_bufMask :2'h0); 
    wire core_ibuf__GEN_23 =( core_ibuf_io_imem_valid ==1'h0| core_ibuf_io_imem_bits_btb_taken ==1'h0| core_ibuf_io_imem_bits_btb_bridx >= core_ibuf_pcWordBits )==1'h0; 
  always @( posedge  core_ibuf_clock )
         begin 
             if ( core_ibuf_reset ==1'h0& core_ibuf__GEN_23 )
                 begin 
                     if (1)$error("Assertion failed\n    at IBuf.scala:79 assert(!io.imem.valid || !io.imem.bits.btb.taken || io.imem.bits.btb.bridx >= pcWordBits)\n");
                     if (1)$fatal;
                 end 
         end
    wire core_ibuf_exp_clock;
    wire core_ibuf_exp_reset;
    wire[31:0] core_ibuf_exp_io_in;
    wire[31:0] core_ibuf_exp_io_out_bits;
    wire[4:0] core_ibuf_exp_io_out_rd;
    wire[4:0] core_ibuf_exp_io_out_rs1;
    wire[4:0] core_ibuf_exp_io_out_rs2;
    wire[4:0] core_ibuf_exp_io_out_rs3;
    wire core_ibuf_exp_io_rvc;

    wire[31:0] core_ibuf_exp_io_out_s_24_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_25_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_26_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_27_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_28_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_29_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_30_bits = core_ibuf_exp_io_in ; 
    wire[31:0] core_ibuf_exp_io_out_s_31_bits = core_ibuf_exp_io_in ; 
    wire[11:0] core_ibuf_exp_io_out_s_jalr_lo =12'hE7; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rd =5'h1; 
    wire[11:0] core_ibuf_exp_io_out_s_jr_lo =12'h67; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs1 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rd =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs2 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rd =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs2 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs1 =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rd =5'h0; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs1 =5'h2; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs1 =5'h2; 
    wire[6:0] core_ibuf_exp_io_out_s_opc =(|( core_ibuf_exp_io_in [12:5])) ? 7'h13:7'h1F; 
    wire[2:0] core_ibuf_exp_io_out_s_lo ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_hi ={ core_ibuf_exp_io_in [10:7], core_ibuf_exp_io_in [12:11]}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi ={ core_ibuf_exp_io_out_s_hi_hi , core_ibuf_exp_io_in [5]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_1 ={{2'h1, core_ibuf_exp_io_in [4:2]}, core_ibuf_exp_io_out_s_opc }; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_hi_1 ={{ core_ibuf_exp_io_out_s_hi , core_ibuf_exp_io_out_s_lo },5'h2}; 
    wire[17:0] core_ibuf_exp_io_out_s_hi_1 ={ core_ibuf_exp_io_out_s_hi_hi_1 ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_0_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_0_bits ={2'h0,{ core_ibuf_exp_io_out_s_hi_1 , core_ibuf_exp_io_out_s_lo_1 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_2 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_2 ={{2'h1, core_ibuf_exp_io_in [4:2]},7'h7}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_2 ={{ core_ibuf_exp_io_out_s_hi_2 ,3'h0},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_3 ={ core_ibuf_exp_io_out_s_hi_hi_2 ,3'h3}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_1_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_1_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_3 , core_ibuf_exp_io_out_s_lo_2 }}; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_3 ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_4 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_4 ={{2'h1, core_ibuf_exp_io_in [4:2]},7'h3}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_hi_3 ={{ core_ibuf_exp_io_out_s_hi_4 , core_ibuf_exp_io_out_s_lo_3 },{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_5 ={ core_ibuf_exp_io_out_s_hi_hi_3 ,3'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_2_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_2_bits ={5'h0,{ core_ibuf_exp_io_out_s_hi_5 , core_ibuf_exp_io_out_s_lo_4 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_6 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_5 ={{2'h1, core_ibuf_exp_io_in [4:2]},7'h3}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_4 ={{ core_ibuf_exp_io_out_s_hi_6 ,3'h0},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_7 ={ core_ibuf_exp_io_out_s_hi_hi_4 ,3'h3}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_3_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_3_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_7 , core_ibuf_exp_io_out_s_lo_5 }}; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_6 ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_8 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[6:0] core_ibuf_exp__GEN ={ core_ibuf_exp_io_out_s_hi_8 , core_ibuf_exp_io_out_s_lo_6 }; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_7 ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_9 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[6:0] core_ibuf_exp__GEN_0 ={ core_ibuf_exp_io_out_s_hi_9 , core_ibuf_exp_io_out_s_lo_7 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi ={3'h2, core_ibuf_exp__GEN_0 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_8 ={ core_ibuf_exp_io_out_s_lo_hi ,7'h3F}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_5 ={ core_ibuf_exp__GEN [6:5],{2'h1, core_ibuf_exp_io_in [4:2]}}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_10 ={ core_ibuf_exp_io_out_s_hi_hi_5 ,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_4_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_4_bits ={5'h0,{ core_ibuf_exp_io_out_s_hi_10 , core_ibuf_exp_io_out_s_lo_8 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_11 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[7:0] core_ibuf_exp__GEN_1 ={ core_ibuf_exp_io_out_s_hi_11 ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_12 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[7:0] core_ibuf_exp__GEN_2 ={ core_ibuf_exp_io_out_s_hi_12 ,3'h0}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_1 ={3'h3, core_ibuf_exp__GEN_2 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_9 ={ core_ibuf_exp_io_out_s_lo_hi_1 ,7'h27}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_6 ={ core_ibuf_exp__GEN_1 [7:5],{2'h1, core_ibuf_exp_io_in [4:2]}}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_13 ={ core_ibuf_exp_io_out_s_hi_hi_6 ,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_5_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_5_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_13 , core_ibuf_exp_io_out_s_lo_9 }}; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_10 ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_14 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[6:0] core_ibuf_exp__GEN_3 ={ core_ibuf_exp_io_out_s_hi_14 , core_ibuf_exp_io_out_s_lo_10 }; 
    wire[2:0] core_ibuf_exp_io_out_s_lo_11 ={ core_ibuf_exp_io_in [6],2'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_15 ={ core_ibuf_exp_io_in [5], core_ibuf_exp_io_in [12:10]}; 
    wire[6:0] core_ibuf_exp__GEN_4 ={ core_ibuf_exp_io_out_s_hi_15 , core_ibuf_exp_io_out_s_lo_11 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_2 ={3'h2, core_ibuf_exp__GEN_4 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_12 ={ core_ibuf_exp_io_out_s_lo_hi_2 ,7'h23}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_7 ={ core_ibuf_exp__GEN_3 [6:5],{2'h1, core_ibuf_exp_io_in [4:2]}}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_16 ={ core_ibuf_exp_io_out_s_hi_hi_7 ,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_6_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_6_bits ={5'h0,{ core_ibuf_exp_io_out_s_hi_16 , core_ibuf_exp_io_out_s_lo_12 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_17 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[7:0] core_ibuf_exp__GEN_5 ={ core_ibuf_exp_io_out_s_hi_17 ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_18 ={ core_ibuf_exp_io_in [6:5], core_ibuf_exp_io_in [12:10]}; 
    wire[7:0] core_ibuf_exp__GEN_6 ={ core_ibuf_exp_io_out_s_hi_18 ,3'h0}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_3 ={3'h3, core_ibuf_exp__GEN_6 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_13 ={ core_ibuf_exp_io_out_s_lo_hi_3 ,7'h23}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_8 ={ core_ibuf_exp__GEN_5 [7:5],{2'h1, core_ibuf_exp_io_in [4:2]}}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_19 ={ core_ibuf_exp_io_out_s_hi_hi_8 ,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rd ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_7_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_7_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_19 , core_ibuf_exp_io_out_s_lo_13 }}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_14 ={ core_ibuf_exp_io_in [11:7],7'h13}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_9 ={{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]}, core_ibuf_exp_io_in [11:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_20 ={ core_ibuf_exp_io_out_s_hi_hi_9 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_8_bits ={ core_ibuf_exp_io_out_s_hi_20 , core_ibuf_exp_io_out_s_lo_14 }; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_8_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_1 =(|( core_ibuf_exp_io_in [11:7])) ? 7'h1B:7'h1F; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_15 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_opc_1 }; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_10 ={{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]}, core_ibuf_exp_io_in [11:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_21 ={ core_ibuf_exp_io_out_s_hi_hi_10 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_9_bits ={ core_ibuf_exp_io_out_s_hi_21 , core_ibuf_exp_io_out_s_lo_15 }; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_9_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_16 ={ core_ibuf_exp_io_in [11:7],7'h13}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_11 ={{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]},5'h0}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_22 ={ core_ibuf_exp_io_out_s_hi_hi_11 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_10_bits ={ core_ibuf_exp_io_out_s_hi_22 , core_ibuf_exp_io_out_s_lo_16 }; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_10_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_2 =(|{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]}) ? 7'h37:7'h3F; 
    wire[19:0] core_ibuf_exp_io_out_s_me_hi ={ core_ibuf_exp_io_in [12] ? 15'h7FFF:15'h0, core_ibuf_exp_io_in [6:2]}; 
    wire[31:0] core_ibuf_exp__GEN_7 ={ core_ibuf_exp_io_out_s_me_hi ,12'h0}; 
    wire[24:0] core_ibuf_exp_io_out_s_me_hi_1 ={ core_ibuf_exp__GEN_7 [31:12], core_ibuf_exp_io_in [11:7]}; 
    wire[31:0] core_ibuf_exp_io_out_s_me_bits ={ core_ibuf_exp_io_out_s_me_hi_1 , core_ibuf_exp_io_out_s_opc_2 }; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_me_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire core_ibuf_exp__GEN_8 = core_ibuf_exp_io_in [11:7]==5'h0| core_ibuf_exp_io_in [11:7]==5'h2; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_3 =(|{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]}) ? 7'h13:7'h1F; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_4 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [6]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_17 ={ core_ibuf_exp_io_out_s_lo_hi_4 ,4'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_hi_hi_12 ={ core_ibuf_exp_io_in [12] ? 3'h7:3'h0, core_ibuf_exp_io_in [4:3]}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_23 ={ core_ibuf_exp_io_out_s_hi_hi_12 , core_ibuf_exp_io_in [5]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_18 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_opc_3 }; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_13 ={{ core_ibuf_exp_io_out_s_hi_23 , core_ibuf_exp_io_out_s_lo_17 }, core_ibuf_exp_io_in [11:7]}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_24 ={ core_ibuf_exp_io_out_s_hi_hi_13 ,3'h0}; 
    wire[31:0] core_ibuf_exp_io_out_s_res_bits ={ core_ibuf_exp_io_out_s_hi_24 , core_ibuf_exp_io_out_s_lo_18 }; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_res_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_11_bits = core_ibuf_exp__GEN_8  ?  core_ibuf_exp_io_out_s_res_bits : core_ibuf_exp_io_out_s_me_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rd = core_ibuf_exp__GEN_8  ?  core_ibuf_exp_io_out_s_res_rd : core_ibuf_exp_io_out_s_me_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs1 = core_ibuf_exp__GEN_8  ?  core_ibuf_exp_io_out_s_res_rs1 : core_ibuf_exp_io_out_s_me_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs2 = core_ibuf_exp__GEN_8  ?  core_ibuf_exp_io_out_s_res_rs2 : core_ibuf_exp_io_out_s_me_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_11_rs3 = core_ibuf_exp__GEN_8  ?  core_ibuf_exp_io_out_s_res_rs3 : core_ibuf_exp_io_out_s_me_rs3 ; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_19 ={{2'h1, core_ibuf_exp_io_in [9:7]},7'h13}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_14 ={{ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:2]},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_25 ={ core_ibuf_exp_io_out_s_hi_hi_14 ,3'h5}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_20 ={{2'h1, core_ibuf_exp_io_in [9:7]},7'h13}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_15 ={{ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:2]},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_26 ={ core_ibuf_exp_io_out_s_hi_hi_15 ,3'h5}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_21 ={{2'h1, core_ibuf_exp_io_in [9:7]},7'h13}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_hi_16 ={{ core_ibuf_exp_io_in [12] ? 7'h7F:7'h0, core_ibuf_exp_io_in [6:2]},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[19:0] core_ibuf_exp_io_out_s_hi_27 ={ core_ibuf_exp_io_out_s_hi_hi_16 ,3'h7}; 
    wire[2:0] core_ibuf_exp__GEN_9 ={ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:5]}; 
    wire[2:0] core_ibuf_exp_io_out_s_funct =(& core_ibuf_exp__GEN_9 ) ? 3'h3: core_ibuf_exp__GEN_9 ==3'h6 ? 3'h2: core_ibuf_exp__GEN_9 ==3'h5 ? 3'h0: core_ibuf_exp__GEN_9 ==3'h4 ? 3'h0: core_ibuf_exp__GEN_9 ==3'h3 ? 3'h7: core_ibuf_exp__GEN_9 ==3'h2 ? 3'h6: core_ibuf_exp__GEN_9 ==3'h1 ? 3'h4:3'h0; 
    wire[30:0] core_ibuf_exp_io_out_s_sub = core_ibuf_exp_io_in [6:5]==2'h0 ? 31'h40000000:31'h0; 
    wire[6:0] core_ibuf_exp_io_out_s_opc_4 = core_ibuf_exp_io_in [12] ? 7'h3B:7'h33; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_22 ={{2'h1, core_ibuf_exp_io_in [9:7]}, core_ibuf_exp_io_out_s_opc_4 }; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_hi_17 ={{2'h1, core_ibuf_exp_io_in [4:2]},{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_28 ={ core_ibuf_exp_io_out_s_hi_hi_17 , core_ibuf_exp_io_out_s_funct }; 
    wire[31:0] core_ibuf_exp_io_out_s_12_bits =(&( core_ibuf_exp_io_in [11:10])) ? {1'h0,{6'h0,{ core_ibuf_exp_io_out_s_hi_28 , core_ibuf_exp_io_out_s_lo_22 }}| core_ibuf_exp_io_out_s_sub }: core_ibuf_exp_io_in [11:10]==2'h2 ? { core_ibuf_exp_io_out_s_hi_27 , core_ibuf_exp_io_out_s_lo_21 }:{1'h0, core_ibuf_exp_io_in [11:10]==2'h1 ? {5'h0,{ core_ibuf_exp_io_out_s_hi_26 , core_ibuf_exp_io_out_s_lo_20 }}|31'h40000000:{5'h0,{ core_ibuf_exp_io_out_s_hi_25 , core_ibuf_exp_io_out_s_lo_19 }}}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rd ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_12_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo ={ core_ibuf_exp_io_in [5:3],1'h0}; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_5 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [11]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_23 ={ core_ibuf_exp_io_out_s_lo_hi_5 , core_ibuf_exp_io_out_s_lo_lo }; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo ={ core_ibuf_exp_io_in [6], core_ibuf_exp_io_in [7]}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi ={ core_ibuf_exp_io_in [12] ? 10'h3FF:10'h0, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_18 ={ core_ibuf_exp_io_out_s_hi_hi_hi , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_29 ={ core_ibuf_exp_io_out_s_hi_hi_18 , core_ibuf_exp_io_out_s_hi_lo }; 
    wire[20:0] core_ibuf_exp__GEN_10 ={ core_ibuf_exp_io_out_s_hi_29 , core_ibuf_exp_io_out_s_lo_23 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_1 ={ core_ibuf_exp_io_in [5:3],1'h0}; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_6 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [11]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_24 ={ core_ibuf_exp_io_out_s_lo_hi_6 , core_ibuf_exp_io_out_s_lo_lo_1 }; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_1 ={ core_ibuf_exp_io_in [6], core_ibuf_exp_io_in [7]}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_1 ={ core_ibuf_exp_io_in [12] ? 10'h3FF:10'h0, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_19 ={ core_ibuf_exp_io_out_s_hi_hi_hi_1 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_30 ={ core_ibuf_exp_io_out_s_hi_hi_19 , core_ibuf_exp_io_out_s_hi_lo_1 }; 
    wire[20:0] core_ibuf_exp__GEN_11 ={ core_ibuf_exp_io_out_s_hi_30 , core_ibuf_exp_io_out_s_lo_24 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_2 ={ core_ibuf_exp_io_in [5:3],1'h0}; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_7 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [11]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_25 ={ core_ibuf_exp_io_out_s_lo_hi_7 , core_ibuf_exp_io_out_s_lo_lo_2 }; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_2 ={ core_ibuf_exp_io_in [6], core_ibuf_exp_io_in [7]}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_2 ={ core_ibuf_exp_io_in [12] ? 10'h3FF:10'h0, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_20 ={ core_ibuf_exp_io_out_s_hi_hi_hi_2 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_31 ={ core_ibuf_exp_io_out_s_hi_hi_20 , core_ibuf_exp_io_out_s_hi_lo_2 }; 
    wire[20:0] core_ibuf_exp__GEN_12 ={ core_ibuf_exp_io_out_s_hi_31 , core_ibuf_exp_io_out_s_lo_25 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_lo_3 ={ core_ibuf_exp_io_in [5:3],1'h0}; 
    wire[1:0] core_ibuf_exp_io_out_s_lo_hi_8 ={ core_ibuf_exp_io_in [2], core_ibuf_exp_io_in [11]}; 
    wire[5:0] core_ibuf_exp_io_out_s_lo_26 ={ core_ibuf_exp_io_out_s_lo_hi_8 , core_ibuf_exp_io_out_s_lo_lo_3 }; 
    wire[1:0] core_ibuf_exp_io_out_s_hi_lo_3 ={ core_ibuf_exp_io_in [6], core_ibuf_exp_io_in [7]}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_hi_3 ={ core_ibuf_exp_io_in [12] ? 10'h3FF:10'h0, core_ibuf_exp_io_in [8]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_21 ={ core_ibuf_exp_io_out_s_hi_hi_hi_3 , core_ibuf_exp_io_in [10:9]}; 
    wire[14:0] core_ibuf_exp_io_out_s_hi_32 ={ core_ibuf_exp_io_out_s_hi_hi_21 , core_ibuf_exp_io_out_s_hi_lo_3 }; 
    wire[20:0] core_ibuf_exp__GEN_13 ={ core_ibuf_exp_io_out_s_hi_32 , core_ibuf_exp_io_out_s_lo_26 }; 
    wire[12:0] core_ibuf_exp_io_out_s_lo_hi_9 ={ core_ibuf_exp__GEN_13 [19:12],5'h0}; 
    wire[19:0] core_ibuf_exp_io_out_s_lo_27 ={ core_ibuf_exp_io_out_s_lo_hi_9 ,7'h6F}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_22 ={ core_ibuf_exp__GEN_10 [20], core_ibuf_exp__GEN_11 [10:1]}; 
    wire[11:0] core_ibuf_exp_io_out_s_hi_33 ={ core_ibuf_exp_io_out_s_hi_hi_22 , core_ibuf_exp__GEN_12 [11]}; 
    wire[31:0] core_ibuf_exp_io_out_s_13_bits ={ core_ibuf_exp_io_out_s_hi_33 , core_ibuf_exp_io_out_s_lo_27 }; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs2 ={2'h1, core_ibuf_exp_io_in [4:2]}; 
    wire[4:0] core_ibuf_exp_io_out_s_13_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_10 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_28 ={ core_ibuf_exp_io_out_s_lo_hi_10 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_23 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_34 ={ core_ibuf_exp_io_out_s_hi_hi_23 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_14 ={ core_ibuf_exp_io_out_s_hi_34 , core_ibuf_exp_io_out_s_lo_28 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_11 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_29 ={ core_ibuf_exp_io_out_s_lo_hi_11 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_24 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_35 ={ core_ibuf_exp_io_out_s_hi_hi_24 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_15 ={ core_ibuf_exp_io_out_s_hi_35 , core_ibuf_exp_io_out_s_lo_29 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_12 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_30 ={ core_ibuf_exp_io_out_s_lo_hi_12 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_25 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_36 ={ core_ibuf_exp_io_out_s_hi_hi_25 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_16 ={ core_ibuf_exp_io_out_s_hi_36 , core_ibuf_exp_io_out_s_lo_30 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_13 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_31 ={ core_ibuf_exp_io_out_s_lo_hi_13 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_26 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_37 ={ core_ibuf_exp_io_out_s_hi_hi_26 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_17 ={ core_ibuf_exp_io_out_s_hi_37 , core_ibuf_exp_io_out_s_lo_31 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_lo_4 ={ core_ibuf_exp__GEN_17 [11],7'h63}; 
    wire[6:0] core_ibuf_exp_io_out_s_lo_hi_14 ={3'h0, core_ibuf_exp__GEN_16 [4:1]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_32 ={ core_ibuf_exp_io_out_s_lo_hi_14 , core_ibuf_exp_io_out_s_lo_lo_4 }; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_lo_4 ={5'h0,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_27 ={ core_ibuf_exp__GEN_14 [12], core_ibuf_exp__GEN_15 [10:5]}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_38 ={ core_ibuf_exp_io_out_s_hi_hi_27 , core_ibuf_exp_io_out_s_hi_lo_4 }; 
    wire[31:0] core_ibuf_exp_io_out_s_14_bits ={ core_ibuf_exp_io_out_s_hi_38 , core_ibuf_exp_io_out_s_lo_32 }; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rd ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_14_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_15 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_33 ={ core_ibuf_exp_io_out_s_lo_hi_15 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_28 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_39 ={ core_ibuf_exp_io_out_s_hi_hi_28 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_18 ={ core_ibuf_exp_io_out_s_hi_39 , core_ibuf_exp_io_out_s_lo_33 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_16 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_34 ={ core_ibuf_exp_io_out_s_lo_hi_16 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_29 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_40 ={ core_ibuf_exp_io_out_s_hi_hi_29 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_19 ={ core_ibuf_exp_io_out_s_hi_40 , core_ibuf_exp_io_out_s_lo_34 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_17 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_35 ={ core_ibuf_exp_io_out_s_lo_hi_17 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_30 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_41 ={ core_ibuf_exp_io_out_s_hi_hi_30 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_20 ={ core_ibuf_exp_io_out_s_hi_41 , core_ibuf_exp_io_out_s_lo_35 }; 
    wire[3:0] core_ibuf_exp_io_out_s_lo_hi_18 ={ core_ibuf_exp_io_in [11:10], core_ibuf_exp_io_in [4:3]}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_36 ={ core_ibuf_exp_io_out_s_lo_hi_18 ,1'h0}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_31 ={ core_ibuf_exp_io_in [12] ? 5'h1F:5'h0, core_ibuf_exp_io_in [6:5]}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_42 ={ core_ibuf_exp_io_out_s_hi_hi_31 , core_ibuf_exp_io_in [2]}; 
    wire[12:0] core_ibuf_exp__GEN_21 ={ core_ibuf_exp_io_out_s_hi_42 , core_ibuf_exp_io_out_s_lo_36 }; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_lo_5 ={ core_ibuf_exp__GEN_21 [11],7'h63}; 
    wire[6:0] core_ibuf_exp_io_out_s_lo_hi_19 ={3'h1, core_ibuf_exp__GEN_20 [4:1]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_37 ={ core_ibuf_exp_io_out_s_lo_hi_19 , core_ibuf_exp_io_out_s_lo_lo_5 }; 
    wire[9:0] core_ibuf_exp_io_out_s_hi_lo_5 ={5'h0,{2'h1, core_ibuf_exp_io_in [9:7]}}; 
    wire[6:0] core_ibuf_exp_io_out_s_hi_hi_32 ={ core_ibuf_exp__GEN_18 [12], core_ibuf_exp__GEN_19 [10:5]}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_43 ={ core_ibuf_exp_io_out_s_hi_hi_32 , core_ibuf_exp_io_out_s_hi_lo_5 }; 
    wire[31:0] core_ibuf_exp_io_out_s_15_bits ={ core_ibuf_exp_io_out_s_hi_43 , core_ibuf_exp_io_out_s_lo_37 }; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs1 ={2'h1, core_ibuf_exp_io_in [9:7]}; 
    wire[4:0] core_ibuf_exp_io_out_s_15_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[6:0] core_ibuf_exp_io_out_s_load_opc =(|( core_ibuf_exp_io_in [11:7])) ? 7'h3:7'h1F; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_38 ={ core_ibuf_exp_io_in [11:7],7'h13}; 
    wire[10:0] core_ibuf_exp_io_out_s_hi_hi_33 ={{ core_ibuf_exp_io_in [12], core_ibuf_exp_io_in [6:2]}, core_ibuf_exp_io_in [11:7]}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_44 ={ core_ibuf_exp_io_out_s_hi_hi_33 ,3'h1}; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_16_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_16_bits ={6'h0,{ core_ibuf_exp_io_out_s_hi_44 , core_ibuf_exp_io_out_s_lo_38 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_39 ={ core_ibuf_exp_io_in [6:5],3'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_45 ={ core_ibuf_exp_io_in [4:2], core_ibuf_exp_io_in [12]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_40 ={ core_ibuf_exp_io_in [11:7],7'h7}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_hi_34 ={{ core_ibuf_exp_io_out_s_hi_45 , core_ibuf_exp_io_out_s_lo_39 },5'h2}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_46 ={ core_ibuf_exp_io_out_s_hi_hi_34 ,3'h3}; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_17_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_17_bits ={3'h0,{ core_ibuf_exp_io_out_s_hi_46 , core_ibuf_exp_io_out_s_lo_40 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_41 ={ core_ibuf_exp_io_in [6:4],2'h0}; 
    wire[2:0] core_ibuf_exp_io_out_s_hi_47 ={ core_ibuf_exp_io_in [3:2], core_ibuf_exp_io_in [12]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_42 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_load_opc }; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_hi_35 ={{ core_ibuf_exp_io_out_s_hi_47 , core_ibuf_exp_io_out_s_lo_41 },5'h2}; 
    wire[15:0] core_ibuf_exp_io_out_s_hi_48 ={ core_ibuf_exp_io_out_s_hi_hi_35 ,3'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_18_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_18_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_48 , core_ibuf_exp_io_out_s_lo_42 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_lo_43 ={ core_ibuf_exp_io_in [6:5],3'h0}; 
    wire[3:0] core_ibuf_exp_io_out_s_hi_49 ={ core_ibuf_exp_io_in [4:2], core_ibuf_exp_io_in [12]}; 
    wire[11:0] core_ibuf_exp_io_out_s_lo_44 ={ core_ibuf_exp_io_in [11:7], core_ibuf_exp_io_out_s_load_opc }; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_hi_36 ={{ core_ibuf_exp_io_out_s_hi_49 , core_ibuf_exp_io_out_s_lo_43 },5'h2}; 
    wire[16:0] core_ibuf_exp_io_out_s_hi_50 ={ core_ibuf_exp_io_out_s_hi_hi_36 ,3'h3}; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_19_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_19_bits ={3'h0,{ core_ibuf_exp_io_out_s_hi_50 , core_ibuf_exp_io_out_s_lo_44 }}; 
    wire[11:0] core_ibuf_exp_io_out_s_mv_lo ={ core_ibuf_exp_io_in [11:7],7'h33}; 
    wire[9:0] core_ibuf_exp_io_out_s_mv_hi_hi ={ core_ibuf_exp_io_in [6:2],5'h0}; 
    wire[12:0] core_ibuf_exp_io_out_s_mv_hi ={ core_ibuf_exp_io_out_s_mv_hi_hi ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_mv_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_mv_bits ={7'h0,{ core_ibuf_exp_io_out_s_mv_hi , core_ibuf_exp_io_out_s_mv_lo }}; 
    wire[11:0] core_ibuf_exp_io_out_s_add_lo ={ core_ibuf_exp_io_in [11:7],7'h33}; 
    wire[9:0] core_ibuf_exp_io_out_s_add_hi_hi ={ core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[12:0] core_ibuf_exp_io_out_s_add_hi ={ core_ibuf_exp_io_out_s_add_hi_hi ,3'h0}; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_add_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_add_bits ={7'h0,{ core_ibuf_exp_io_out_s_add_hi , core_ibuf_exp_io_out_s_add_lo }}; 
    wire[9:0] core_ibuf_exp_io_out_s_jr_hi_hi ={ core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[12:0] core_ibuf_exp_io_out_s_jr_hi ={ core_ibuf_exp_io_out_s_jr_hi_hi ,3'h0}; 
    wire[24:0] core_ibuf_exp_io_out_s_jr ={ core_ibuf_exp_io_out_s_jr_hi , core_ibuf_exp_io_out_s_jr_lo }; 
    wire[24:0] core_ibuf_exp_io_out_s_reserved ={ core_ibuf_exp_io_out_s_jr [24:7],7'h1F}; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_reserved_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_jr_reserved_bits ={7'h0,(|( core_ibuf_exp_io_in [11:7])) ?  core_ibuf_exp_io_out_s_jr : core_ibuf_exp_io_out_s_reserved }; 
    wire core_ibuf_exp__GEN_22 =|( core_ibuf_exp_io_in [6:2]); 
    wire[31:0] core_ibuf_exp_io_out_s_jr_mv_bits = core_ibuf_exp__GEN_22  ?  core_ibuf_exp_io_out_s_mv_bits : core_ibuf_exp_io_out_s_jr_reserved_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rd = core_ibuf_exp__GEN_22  ?  core_ibuf_exp_io_out_s_mv_rd : core_ibuf_exp_io_out_s_jr_reserved_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs1 = core_ibuf_exp__GEN_22  ?  core_ibuf_exp_io_out_s_mv_rs1 : core_ibuf_exp_io_out_s_jr_reserved_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs2 = core_ibuf_exp__GEN_22  ?  core_ibuf_exp_io_out_s_mv_rs2 : core_ibuf_exp_io_out_s_jr_reserved_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jr_mv_rs3 = core_ibuf_exp__GEN_22  ?  core_ibuf_exp_io_out_s_mv_rs3 : core_ibuf_exp_io_out_s_jr_reserved_rs3 ; 
    wire[9:0] core_ibuf_exp_io_out_s_jalr_hi_hi ={ core_ibuf_exp_io_in [6:2], core_ibuf_exp_io_in [11:7]}; 
    wire[12:0] core_ibuf_exp_io_out_s_jalr_hi ={ core_ibuf_exp_io_out_s_jalr_hi_hi ,3'h0}; 
    wire[24:0] core_ibuf_exp_io_out_s_jalr ={ core_ibuf_exp_io_out_s_jalr_hi , core_ibuf_exp_io_out_s_jalr_lo }; 
    wire[24:0] core_ibuf_exp_io_out_s_ebreak ={ core_ibuf_exp_io_out_s_jr [24:7],7'h73}|25'h100000; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs1 = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_ebreak_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_jalr_ebreak_bits ={7'h0,(|( core_ibuf_exp_io_in [11:7])) ?  core_ibuf_exp_io_out_s_jalr : core_ibuf_exp_io_out_s_ebreak }; 
    wire core_ibuf_exp__GEN_23 =|( core_ibuf_exp_io_in [6:2]); 
    wire[31:0] core_ibuf_exp_io_out_s_jalr_add_bits = core_ibuf_exp__GEN_23  ?  core_ibuf_exp_io_out_s_add_bits : core_ibuf_exp_io_out_s_jalr_ebreak_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rd = core_ibuf_exp__GEN_23  ?  core_ibuf_exp_io_out_s_add_rd : core_ibuf_exp_io_out_s_jalr_ebreak_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs1 = core_ibuf_exp__GEN_23  ?  core_ibuf_exp_io_out_s_add_rs1 : core_ibuf_exp_io_out_s_jalr_ebreak_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs2 = core_ibuf_exp__GEN_23  ?  core_ibuf_exp_io_out_s_add_rs2 : core_ibuf_exp_io_out_s_jalr_ebreak_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_jalr_add_rs3 = core_ibuf_exp__GEN_23  ?  core_ibuf_exp_io_out_s_add_rs3 : core_ibuf_exp_io_out_s_jalr_ebreak_rs3 ; 
    wire[31:0] core_ibuf_exp_io_out_s_20_bits = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_bits : core_ibuf_exp_io_out_s_jr_mv_bits ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rd = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rd : core_ibuf_exp_io_out_s_jr_mv_rd ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs1 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs1 : core_ibuf_exp_io_out_s_jr_mv_rs1 ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs2 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs2 : core_ibuf_exp_io_out_s_jr_mv_rs2 ; 
    wire[4:0] core_ibuf_exp_io_out_s_20_rs3 = core_ibuf_exp_io_in [12] ?  core_ibuf_exp_io_out_s_jalr_add_rs3 : core_ibuf_exp_io_out_s_jr_mv_rs3 ; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_51 ={ core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_in [12:10]}; 
    wire[8:0] core_ibuf_exp__GEN_24 ={ core_ibuf_exp_io_out_s_hi_51 ,3'h0}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_52 ={ core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_in [12:10]}; 
    wire[8:0] core_ibuf_exp__GEN_25 ={ core_ibuf_exp_io_out_s_hi_52 ,3'h0}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_20 ={3'h3, core_ibuf_exp__GEN_25 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_45 ={ core_ibuf_exp_io_out_s_lo_hi_20 ,7'h27}; 
    wire[8:0] core_ibuf_exp_io_out_s_hi_hi_37 ={ core_ibuf_exp__GEN_24 [8:5], core_ibuf_exp_io_in [6:2]}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_53 ={ core_ibuf_exp_io_out_s_hi_hi_37 ,5'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_21_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_21_bits ={3'h0,{ core_ibuf_exp_io_out_s_hi_53 , core_ibuf_exp_io_out_s_lo_45 }}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_54 ={ core_ibuf_exp_io_in [8:7], core_ibuf_exp_io_in [12:9]}; 
    wire[7:0] core_ibuf_exp__GEN_26 ={ core_ibuf_exp_io_out_s_hi_54 ,2'h0}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_55 ={ core_ibuf_exp_io_in [8:7], core_ibuf_exp_io_in [12:9]}; 
    wire[7:0] core_ibuf_exp__GEN_27 ={ core_ibuf_exp_io_out_s_hi_55 ,2'h0}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_21 ={3'h2, core_ibuf_exp__GEN_27 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_46 ={ core_ibuf_exp_io_out_s_lo_hi_21 ,7'h23}; 
    wire[7:0] core_ibuf_exp_io_out_s_hi_hi_38 ={ core_ibuf_exp__GEN_26 [7:5], core_ibuf_exp_io_in [6:2]}; 
    wire[12:0] core_ibuf_exp_io_out_s_hi_56 ={ core_ibuf_exp_io_out_s_hi_hi_38 ,5'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_22_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_22_bits ={4'h0,{ core_ibuf_exp_io_out_s_hi_56 , core_ibuf_exp_io_out_s_lo_46 }}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_57 ={ core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_in [12:10]}; 
    wire[8:0] core_ibuf_exp__GEN_28 ={ core_ibuf_exp_io_out_s_hi_57 ,3'h0}; 
    wire[5:0] core_ibuf_exp_io_out_s_hi_58 ={ core_ibuf_exp_io_in [9:7], core_ibuf_exp_io_in [12:10]}; 
    wire[8:0] core_ibuf_exp__GEN_29 ={ core_ibuf_exp_io_out_s_hi_58 ,3'h0}; 
    wire[7:0] core_ibuf_exp_io_out_s_lo_hi_22 ={3'h3, core_ibuf_exp__GEN_29 [4:0]}; 
    wire[14:0] core_ibuf_exp_io_out_s_lo_47 ={ core_ibuf_exp_io_out_s_lo_hi_22 ,7'h23}; 
    wire[8:0] core_ibuf_exp_io_out_s_hi_hi_39 ={ core_ibuf_exp__GEN_28 [8:5], core_ibuf_exp_io_in [6:2]}; 
    wire[13:0] core_ibuf_exp_io_out_s_hi_59 ={ core_ibuf_exp_io_out_s_hi_hi_39 ,5'h2}; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs2 = core_ibuf_exp_io_in [6:2]; 
    wire[4:0] core_ibuf_exp_io_out_s_23_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[31:0] core_ibuf_exp_io_out_s_23_bits ={3'h0,{ core_ibuf_exp_io_out_s_hi_59 , core_ibuf_exp_io_out_s_lo_47 }}; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_24_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_25_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_26_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_27_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_28_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_29_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_30_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rd = core_ibuf_exp_io_in [11:7]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs1 = core_ibuf_exp_io_in [19:15]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs2 = core_ibuf_exp_io_in [24:20]; 
    wire[4:0] core_ibuf_exp_io_out_s_31_rs3 = core_ibuf_exp_io_in [31:27]; 
    wire[4:0] core_ibuf_exp__GEN_30 ={ core_ibuf_exp_io_in [1:0], core_ibuf_exp_io_in [15:13]}; 
    wire core_ibuf_exp__GEN_31 = core_ibuf_exp__GEN_30 ==5'h1; 
    wire core_ibuf_exp__GEN_32 = core_ibuf_exp__GEN_30 ==5'h2; 
    wire core_ibuf_exp__GEN_33 = core_ibuf_exp__GEN_30 ==5'h3; 
    wire core_ibuf_exp__GEN_34 = core_ibuf_exp__GEN_30 ==5'h4; 
    wire core_ibuf_exp__GEN_35 = core_ibuf_exp__GEN_30 ==5'h5; 
    wire core_ibuf_exp__GEN_36 = core_ibuf_exp__GEN_30 ==5'h6; 
    wire core_ibuf_exp__GEN_37 = core_ibuf_exp__GEN_30 ==5'h7; 
    wire core_ibuf_exp__GEN_38 = core_ibuf_exp__GEN_30 ==5'h8; 
    wire core_ibuf_exp__GEN_39 = core_ibuf_exp__GEN_30 ==5'h9; 
    wire core_ibuf_exp__GEN_40 = core_ibuf_exp__GEN_30 ==5'hA; 
    wire core_ibuf_exp__GEN_41 = core_ibuf_exp__GEN_30 ==5'hB; 
    wire core_ibuf_exp__GEN_42 = core_ibuf_exp__GEN_30 ==5'hC; 
    wire core_ibuf_exp__GEN_43 = core_ibuf_exp__GEN_30 ==5'hD; 
    wire core_ibuf_exp__GEN_44 = core_ibuf_exp__GEN_30 ==5'hE; 
    wire core_ibuf_exp__GEN_45 = core_ibuf_exp__GEN_30 ==5'hF; 
    wire core_ibuf_exp__GEN_46 = core_ibuf_exp__GEN_30 ==5'h10; 
    wire core_ibuf_exp__GEN_47 = core_ibuf_exp__GEN_30 ==5'h11; 
    wire core_ibuf_exp__GEN_48 = core_ibuf_exp__GEN_30 ==5'h12; 
    wire core_ibuf_exp__GEN_49 = core_ibuf_exp__GEN_30 ==5'h13; 
    wire core_ibuf_exp__GEN_50 = core_ibuf_exp__GEN_30 ==5'h14; 
    wire core_ibuf_exp__GEN_51 = core_ibuf_exp__GEN_30 ==5'h15; 
    wire core_ibuf_exp__GEN_52 = core_ibuf_exp__GEN_30 ==5'h16; 
    wire core_ibuf_exp__GEN_53 = core_ibuf_exp__GEN_30 ==5'h17; 
    wire core_ibuf_exp__GEN_54 = core_ibuf_exp__GEN_30 ==5'h18; 
    wire core_ibuf_exp__GEN_55 = core_ibuf_exp__GEN_30 ==5'h19; 
    wire core_ibuf_exp__GEN_56 = core_ibuf_exp__GEN_30 ==5'h1A; 
    wire core_ibuf_exp__GEN_57 = core_ibuf_exp__GEN_30 ==5'h1B; 
    wire core_ibuf_exp__GEN_58 = core_ibuf_exp__GEN_30 ==5'h1C; 
    wire core_ibuf_exp__GEN_59 = core_ibuf_exp__GEN_30 ==5'h1D; 
    wire core_ibuf_exp__GEN_60 = core_ibuf_exp__GEN_30 ==5'h1E; 
    wire core_ibuf_exp__GEN_61 =& core_ibuf_exp__GEN_30 ; 
  assign  core_ibuf_exp_io_out_bits = core_ibuf_exp__GEN_61  ?  core_ibuf_exp_io_out_s_31_bits : core_ibuf_exp__GEN_60  ?  core_ibuf_exp_io_out_s_30_bits : core_ibuf_exp__GEN_59  ?  core_ibuf_exp_io_out_s_29_bits : core_ibuf_exp__GEN_58  ?  core_ibuf_exp_io_out_s_28_bits : core_ibuf_exp__GEN_57  ?  core_ibuf_exp_io_out_s_27_bits : core_ibuf_exp__GEN_56  ?  core_ibuf_exp_io_out_s_26_bits : core_ibuf_exp__GEN_55  ?  core_ibuf_exp_io_out_s_25_bits : core_ibuf_exp__GEN_54  ?  core_ibuf_exp_io_out_s_24_bits : core_ibuf_exp__GEN_53  ?  core_ibuf_exp_io_out_s_23_bits : core_ibuf_exp__GEN_52  ?  core_ibuf_exp_io_out_s_22_bits : core_ibuf_exp__GEN_51  ?  core_ibuf_exp_io_out_s_21_bits : core_ibuf_exp__GEN_50  ?  core_ibuf_exp_io_out_s_20_bits : core_ibuf_exp__GEN_49  ?  core_ibuf_exp_io_out_s_19_bits : core_ibuf_exp__GEN_48  ?  core_ibuf_exp_io_out_s_18_bits : core_ibuf_exp__GEN_47  ?  core_ibuf_exp_io_out_s_17_bits : core_ibuf_exp__GEN_46  ?  core_ibuf_exp_io_out_s_16_bits : core_ibuf_exp__GEN_45  ?  core_ibuf_exp_io_out_s_15_bits : core_ibuf_exp__GEN_44  ?  core_ibuf_exp_io_out_s_14_bits : core_ibuf_exp__GEN_43  ?  core_ibuf_exp_io_out_s_13_bits : core_ibuf_exp__GEN_42  ?  core_ibuf_exp_io_out_s_12_bits : core_ibuf_exp__GEN_41  ?  core_ibuf_exp_io_out_s_11_bits : core_ibuf_exp__GEN_40  ?  core_ibuf_exp_io_out_s_10_bits : core_ibuf_exp__GEN_39  ?  core_ibuf_exp_io_out_s_9_bits : core_ibuf_exp__GEN_38  ?  core_ibuf_exp_io_out_s_8_bits : core_ibuf_exp__GEN_37  ?  core_ibuf_exp_io_out_s_7_bits : core_ibuf_exp__GEN_36  ?  core_ibuf_exp_io_out_s_6_bits : core_ibuf_exp__GEN_35  ?  core_ibuf_exp_io_out_s_5_bits : core_ibuf_exp__GEN_34  ?  core_ibuf_exp_io_out_s_4_bits : core_ibuf_exp__GEN_33  ?  core_ibuf_exp_io_out_s_3_bits : core_ibuf_exp__GEN_32  ?  core_ibuf_exp_io_out_s_2_bits : core_ibuf_exp__GEN_31  ?  core_ibuf_exp_io_out_s_1_bits : core_ibuf_exp_io_out_s_0_bits ; 
  assign  core_ibuf_exp_io_out_rd = core_ibuf_exp__GEN_61  ?  core_ibuf_exp_io_out_s_31_rd : core_ibuf_exp__GEN_60  ?  core_ibuf_exp_io_out_s_30_rd : core_ibuf_exp__GEN_59  ?  core_ibuf_exp_io_out_s_29_rd : core_ibuf_exp__GEN_58  ?  core_ibuf_exp_io_out_s_28_rd : core_ibuf_exp__GEN_57  ?  core_ibuf_exp_io_out_s_27_rd : core_ibuf_exp__GEN_56  ?  core_ibuf_exp_io_out_s_26_rd : core_ibuf_exp__GEN_55  ?  core_ibuf_exp_io_out_s_25_rd : core_ibuf_exp__GEN_54  ?  core_ibuf_exp_io_out_s_24_rd : core_ibuf_exp__GEN_53  ?  core_ibuf_exp_io_out_s_23_rd : core_ibuf_exp__GEN_52  ?  core_ibuf_exp_io_out_s_22_rd : core_ibuf_exp__GEN_51  ?  core_ibuf_exp_io_out_s_21_rd : core_ibuf_exp__GEN_50  ?  core_ibuf_exp_io_out_s_20_rd : core_ibuf_exp__GEN_49  ?  core_ibuf_exp_io_out_s_19_rd : core_ibuf_exp__GEN_48  ?  core_ibuf_exp_io_out_s_18_rd : core_ibuf_exp__GEN_47  ?  core_ibuf_exp_io_out_s_17_rd : core_ibuf_exp__GEN_46  ?  core_ibuf_exp_io_out_s_16_rd : core_ibuf_exp__GEN_45  ?  core_ibuf_exp_io_out_s_15_rd : core_ibuf_exp__GEN_44  ?  core_ibuf_exp_io_out_s_14_rd : core_ibuf_exp__GEN_43  ?  core_ibuf_exp_io_out_s_13_rd : core_ibuf_exp__GEN_42  ?  core_ibuf_exp_io_out_s_12_rd : core_ibuf_exp__GEN_41  ?  core_ibuf_exp_io_out_s_11_rd : core_ibuf_exp__GEN_40  ?  core_ibuf_exp_io_out_s_10_rd : core_ibuf_exp__GEN_39  ?  core_ibuf_exp_io_out_s_9_rd : core_ibuf_exp__GEN_38  ?  core_ibuf_exp_io_out_s_8_rd : core_ibuf_exp__GEN_37  ?  core_ibuf_exp_io_out_s_7_rd : core_ibuf_exp__GEN_36  ?  core_ibuf_exp_io_out_s_6_rd : core_ibuf_exp__GEN_35  ?  core_ibuf_exp_io_out_s_5_rd : core_ibuf_exp__GEN_34  ?  core_ibuf_exp_io_out_s_4_rd : core_ibuf_exp__GEN_33  ?  core_ibuf_exp_io_out_s_3_rd : core_ibuf_exp__GEN_32  ?  core_ibuf_exp_io_out_s_2_rd : core_ibuf_exp__GEN_31  ?  core_ibuf_exp_io_out_s_1_rd : core_ibuf_exp_io_out_s_0_rd ; 
  assign  core_ibuf_exp_io_out_rs1 = core_ibuf_exp__GEN_61  ?  core_ibuf_exp_io_out_s_31_rs1 : core_ibuf_exp__GEN_60  ?  core_ibuf_exp_io_out_s_30_rs1 : core_ibuf_exp__GEN_59  ?  core_ibuf_exp_io_out_s_29_rs1 : core_ibuf_exp__GEN_58  ?  core_ibuf_exp_io_out_s_28_rs1 : core_ibuf_exp__GEN_57  ?  core_ibuf_exp_io_out_s_27_rs1 : core_ibuf_exp__GEN_56  ?  core_ibuf_exp_io_out_s_26_rs1 : core_ibuf_exp__GEN_55  ?  core_ibuf_exp_io_out_s_25_rs1 : core_ibuf_exp__GEN_54  ?  core_ibuf_exp_io_out_s_24_rs1 : core_ibuf_exp__GEN_53  ?  core_ibuf_exp_io_out_s_23_rs1 : core_ibuf_exp__GEN_52  ?  core_ibuf_exp_io_out_s_22_rs1 : core_ibuf_exp__GEN_51  ?  core_ibuf_exp_io_out_s_21_rs1 : core_ibuf_exp__GEN_50  ?  core_ibuf_exp_io_out_s_20_rs1 : core_ibuf_exp__GEN_49  ?  core_ibuf_exp_io_out_s_19_rs1 : core_ibuf_exp__GEN_48  ?  core_ibuf_exp_io_out_s_18_rs1 : core_ibuf_exp__GEN_47  ?  core_ibuf_exp_io_out_s_17_rs1 : core_ibuf_exp__GEN_46  ?  core_ibuf_exp_io_out_s_16_rs1 : core_ibuf_exp__GEN_45  ?  core_ibuf_exp_io_out_s_15_rs1 : core_ibuf_exp__GEN_44  ?  core_ibuf_exp_io_out_s_14_rs1 : core_ibuf_exp__GEN_43  ?  core_ibuf_exp_io_out_s_13_rs1 : core_ibuf_exp__GEN_42  ?  core_ibuf_exp_io_out_s_12_rs1 : core_ibuf_exp__GEN_41  ?  core_ibuf_exp_io_out_s_11_rs1 : core_ibuf_exp__GEN_40  ?  core_ibuf_exp_io_out_s_10_rs1 : core_ibuf_exp__GEN_39  ?  core_ibuf_exp_io_out_s_9_rs1 : core_ibuf_exp__GEN_38  ?  core_ibuf_exp_io_out_s_8_rs1 : core_ibuf_exp__GEN_37  ?  core_ibuf_exp_io_out_s_7_rs1 : core_ibuf_exp__GEN_36  ?  core_ibuf_exp_io_out_s_6_rs1 : core_ibuf_exp__GEN_35  ?  core_ibuf_exp_io_out_s_5_rs1 : core_ibuf_exp__GEN_34  ?  core_ibuf_exp_io_out_s_4_rs1 : core_ibuf_exp__GEN_33  ?  core_ibuf_exp_io_out_s_3_rs1 : core_ibuf_exp__GEN_32  ?  core_ibuf_exp_io_out_s_2_rs1 : core_ibuf_exp__GEN_31  ?  core_ibuf_exp_io_out_s_1_rs1 : core_ibuf_exp_io_out_s_0_rs1 ; 
  assign  core_ibuf_exp_io_out_rs2 = core_ibuf_exp__GEN_61  ?  core_ibuf_exp_io_out_s_31_rs2 : core_ibuf_exp__GEN_60  ?  core_ibuf_exp_io_out_s_30_rs2 : core_ibuf_exp__GEN_59  ?  core_ibuf_exp_io_out_s_29_rs2 : core_ibuf_exp__GEN_58  ?  core_ibuf_exp_io_out_s_28_rs2 : core_ibuf_exp__GEN_57  ?  core_ibuf_exp_io_out_s_27_rs2 : core_ibuf_exp__GEN_56  ?  core_ibuf_exp_io_out_s_26_rs2 : core_ibuf_exp__GEN_55  ?  core_ibuf_exp_io_out_s_25_rs2 : core_ibuf_exp__GEN_54  ?  core_ibuf_exp_io_out_s_24_rs2 : core_ibuf_exp__GEN_53  ?  core_ibuf_exp_io_out_s_23_rs2 : core_ibuf_exp__GEN_52  ?  core_ibuf_exp_io_out_s_22_rs2 : core_ibuf_exp__GEN_51  ?  core_ibuf_exp_io_out_s_21_rs2 : core_ibuf_exp__GEN_50  ?  core_ibuf_exp_io_out_s_20_rs2 : core_ibuf_exp__GEN_49  ?  core_ibuf_exp_io_out_s_19_rs2 : core_ibuf_exp__GEN_48  ?  core_ibuf_exp_io_out_s_18_rs2 : core_ibuf_exp__GEN_47  ?  core_ibuf_exp_io_out_s_17_rs2 : core_ibuf_exp__GEN_46  ?  core_ibuf_exp_io_out_s_16_rs2 : core_ibuf_exp__GEN_45  ?  core_ibuf_exp_io_out_s_15_rs2 : core_ibuf_exp__GEN_44  ?  core_ibuf_exp_io_out_s_14_rs2 : core_ibuf_exp__GEN_43  ?  core_ibuf_exp_io_out_s_13_rs2 : core_ibuf_exp__GEN_42  ?  core_ibuf_exp_io_out_s_12_rs2 : core_ibuf_exp__GEN_41  ?  core_ibuf_exp_io_out_s_11_rs2 : core_ibuf_exp__GEN_40  ?  core_ibuf_exp_io_out_s_10_rs2 : core_ibuf_exp__GEN_39  ?  core_ibuf_exp_io_out_s_9_rs2 : core_ibuf_exp__GEN_38  ?  core_ibuf_exp_io_out_s_8_rs2 : core_ibuf_exp__GEN_37  ?  core_ibuf_exp_io_out_s_7_rs2 : core_ibuf_exp__GEN_36  ?  core_ibuf_exp_io_out_s_6_rs2 : core_ibuf_exp__GEN_35  ?  core_ibuf_exp_io_out_s_5_rs2 : core_ibuf_exp__GEN_34  ?  core_ibuf_exp_io_out_s_4_rs2 : core_ibuf_exp__GEN_33  ?  core_ibuf_exp_io_out_s_3_rs2 : core_ibuf_exp__GEN_32  ?  core_ibuf_exp_io_out_s_2_rs2 : core_ibuf_exp__GEN_31  ?  core_ibuf_exp_io_out_s_1_rs2 : core_ibuf_exp_io_out_s_0_rs2 ; 
  assign  core_ibuf_exp_io_out_rs3 = core_ibuf_exp__GEN_61  ?  core_ibuf_exp_io_out_s_31_rs3 : core_ibuf_exp__GEN_60  ?  core_ibuf_exp_io_out_s_30_rs3 : core_ibuf_exp__GEN_59  ?  core_ibuf_exp_io_out_s_29_rs3 : core_ibuf_exp__GEN_58  ?  core_ibuf_exp_io_out_s_28_rs3 : core_ibuf_exp__GEN_57  ?  core_ibuf_exp_io_out_s_27_rs3 : core_ibuf_exp__GEN_56  ?  core_ibuf_exp_io_out_s_26_rs3 : core_ibuf_exp__GEN_55  ?  core_ibuf_exp_io_out_s_25_rs3 : core_ibuf_exp__GEN_54  ?  core_ibuf_exp_io_out_s_24_rs3 : core_ibuf_exp__GEN_53  ?  core_ibuf_exp_io_out_s_23_rs3 : core_ibuf_exp__GEN_52  ?  core_ibuf_exp_io_out_s_22_rs3 : core_ibuf_exp__GEN_51  ?  core_ibuf_exp_io_out_s_21_rs3 : core_ibuf_exp__GEN_50  ?  core_ibuf_exp_io_out_s_20_rs3 : core_ibuf_exp__GEN_49  ?  core_ibuf_exp_io_out_s_19_rs3 : core_ibuf_exp__GEN_48  ?  core_ibuf_exp_io_out_s_18_rs3 : core_ibuf_exp__GEN_47  ?  core_ibuf_exp_io_out_s_17_rs3 : core_ibuf_exp__GEN_46  ?  core_ibuf_exp_io_out_s_16_rs3 : core_ibuf_exp__GEN_45  ?  core_ibuf_exp_io_out_s_15_rs3 : core_ibuf_exp__GEN_44  ?  core_ibuf_exp_io_out_s_14_rs3 : core_ibuf_exp__GEN_43  ?  core_ibuf_exp_io_out_s_13_rs3 : core_ibuf_exp__GEN_42  ?  core_ibuf_exp_io_out_s_12_rs3 : core_ibuf_exp__GEN_41  ?  core_ibuf_exp_io_out_s_11_rs3 : core_ibuf_exp__GEN_40  ?  core_ibuf_exp_io_out_s_10_rs3 : core_ibuf_exp__GEN_39  ?  core_ibuf_exp_io_out_s_9_rs3 : core_ibuf_exp__GEN_38  ?  core_ibuf_exp_io_out_s_8_rs3 : core_ibuf_exp__GEN_37  ?  core_ibuf_exp_io_out_s_7_rs3 : core_ibuf_exp__GEN_36  ?  core_ibuf_exp_io_out_s_6_rs3 : core_ibuf_exp__GEN_35  ?  core_ibuf_exp_io_out_s_5_rs3 : core_ibuf_exp__GEN_34  ?  core_ibuf_exp_io_out_s_4_rs3 : core_ibuf_exp__GEN_33  ?  core_ibuf_exp_io_out_s_3_rs3 : core_ibuf_exp__GEN_32  ?  core_ibuf_exp_io_out_s_2_rs3 : core_ibuf_exp__GEN_31  ?  core_ibuf_exp_io_out_s_1_rs3 : core_ibuf_exp_io_out_s_0_rs3 ; 
  assign  core_ibuf_exp_io_rvc = core_ibuf_exp_io_in [1:0]!=2'h3;
    assign core_ibuf_exp_clock = core_ibuf_clock;
    assign core_ibuf_exp_reset = core_ibuf_reset;
    assign core_ibuf_exp_io_in = core_ibuf_inst;
    assign core_ibuf_io_inst_0_bits_inst_bits = core_ibuf_exp_io_out_bits;
    assign core_ibuf_io_inst_0_bits_inst_rd = core_ibuf_exp_io_out_rd;
    assign core_ibuf_io_inst_0_bits_inst_rs1 = core_ibuf_exp_io_out_rs1;
    assign core_ibuf_io_inst_0_bits_inst_rs2 = core_ibuf_exp_io_out_rs2;
    assign core_ibuf_io_inst_0_bits_inst_rs3 = core_ibuf_exp_io_out_rs3;
    assign core_ibuf__exp_io_rvc = core_ibuf_exp_io_rvc;
     
    wire[1:0] core_ibuf__GEN_24 = core_ibuf_ic_replay >>2'h1; 
    wire core_ibuf_replay = core_ibuf_ic_replay [0]| core_ibuf__exp_io_rvc ==1'h0& core_ibuf__GEN_24 [0]; 
    wire[1:0] core_ibuf__GEN_25 = core_ibuf_valid >>2'h1; 
    wire core_ibuf_full_insn = core_ibuf__exp_io_rvc | core_ibuf__GEN_25 [0]| core_ibuf_buf_replay_0 [0]; 
    wire[1:0] core_ibuf_io_inst_0_bits_xcpt1_hi ={ core_ibuf_xcpt_1_pf_inst , core_ibuf_xcpt_1_gf_inst }; 
    wire[2:0] core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 = core_ibuf__exp_io_rvc  ? 3'h0:{ core_ibuf_io_inst_0_bits_xcpt1_hi , core_ibuf_xcpt_1_ae_inst }; 
    wire core_ibuf__io_inst_0_bits_xcpt1_WIRE_ae_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [0]; 
    wire core_ibuf__io_inst_0_bits_xcpt1_WIRE_gf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [1]; 
    wire core_ibuf__io_inst_0_bits_xcpt1_WIRE_pf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_1 [2]; 
    wire[1:0] core_ibuf__GEN_26 = core_ibuf_bufMask >>2'h1; 
    wire core_ibuf__GEN_27 = core_ibuf_bufMask [0]& core_ibuf__exp_io_rvc | core_ibuf__GEN_26 [0]; 
  assign  core_ibuf_nReady = core_ibuf_full_insn  ? ( core_ibuf__exp_io_rvc  ? 2'h1:2'h2):2'h0; 
  always @( posedge  core_ibuf_clock )
         begin 
             if ( core_ibuf_reset ) 
                 core_ibuf_nBufValid  <=1'h0;
              else 
                 if ( core_ibuf_io_kill ) 
                     core_ibuf_nBufValid  <=1'h0;
                  else 
                     if ( core_ibuf_io_inst_0_ready )
                         begin 
                             if ( core_ibuf__GEN_6 ) 
                                 core_ibuf_nBufValid  <= core_ibuf__GEN_9 [0];
                              else  
                                 core_ibuf_nBufValid  <= core_ibuf__GEN_4 [0];
                         end 
                      else 
                         begin 
                         end 
         end
  always @( posedge  core_ibuf_clock )
         begin 
             if ( core_ibuf_io_inst_0_ready )
                 begin 
                     if ( core_ibuf__GEN_6 )
                         begin  
                             core_ibuf_buf_btb_cfiType  <= core_ibuf_io_imem_bits_btb_cfiType ; 
                             core_ibuf_buf_btb_taken  <= core_ibuf_io_imem_bits_btb_taken ; 
                             core_ibuf_buf_btb_mask  <= core_ibuf_io_imem_bits_btb_mask ; 
                             core_ibuf_buf_btb_bridx  <= core_ibuf_io_imem_bits_btb_bridx ; 
                             core_ibuf_buf_btb_target  <= core_ibuf_io_imem_bits_btb_target ; 
                             core_ibuf_buf_btb_entry  <= core_ibuf_io_imem_bits_btb_entry ; 
                             core_ibuf_buf_btb_bht_history  <= core_ibuf_io_imem_bits_btb_bht_history ; 
                             core_ibuf_buf_btb_bht_value  <= core_ibuf_io_imem_bits_btb_bht_value ; 
                             core_ibuf_buf_pc  <= core_ibuf__GEN_13 ; 
                             core_ibuf_buf_data  <= core_ibuf__GEN_11 ; 
                             core_ibuf_buf_mask  <= core_ibuf_io_imem_bits_mask ; 
                             core_ibuf_buf_xcpt_pf_inst  <= core_ibuf_io_imem_bits_xcpt_pf_inst ; 
                             core_ibuf_buf_xcpt_gf_inst  <= core_ibuf_io_imem_bits_xcpt_gf_inst ; 
                             core_ibuf_buf_xcpt_ae_inst  <= core_ibuf_io_imem_bits_xcpt_ae_inst ; 
                             core_ibuf_buf_replay  <= core_ibuf_io_imem_bits_replay ; 
                             core_ibuf_ibufBTBResp_cfiType  <= core_ibuf_io_imem_bits_btb_cfiType ; 
                             core_ibuf_ibufBTBResp_taken  <= core_ibuf_io_imem_bits_btb_taken ; 
                             core_ibuf_ibufBTBResp_mask  <= core_ibuf_io_imem_bits_btb_mask ; 
                             core_ibuf_ibufBTBResp_bridx  <= core_ibuf_io_imem_bits_btb_bridx ; 
                             core_ibuf_ibufBTBResp_target  <= core_ibuf_io_imem_bits_btb_target ; 
                             core_ibuf_ibufBTBResp_entry  <= core_ibuf_io_imem_bits_btb_entry ; 
                             core_ibuf_ibufBTBResp_bht_history  <= core_ibuf_io_imem_bits_btb_bht_history ; 
                             core_ibuf_ibufBTBResp_bht_value  <= core_ibuf_io_imem_bits_btb_bht_value ;
                         end 
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end 
         end
  assign  core_ibuf_io_imem_ready = core_ibuf_io_inst_0_ready & core_ibuf_nReady >={1'h0, core_ibuf_nBufValid }&( core_ibuf_nICReady >= core_ibuf_nIC |2'h1>= core_ibuf__GEN_2 [1:0]); 
  assign  core_ibuf_io_pc = core_ibuf_nBufValid >1'h0 ?  core_ibuf_buf_pc : core_ibuf_io_imem_bits_pc ; 
  assign  core_ibuf_io_btb_resp_cfiType = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_cfiType : core_ibuf_io_imem_bits_btb_cfiType ; 
  assign  core_ibuf_io_btb_resp_taken = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_taken : core_ibuf_io_imem_bits_btb_taken ; 
  assign  core_ibuf_io_btb_resp_mask = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_mask : core_ibuf_io_imem_bits_btb_mask ; 
  assign  core_ibuf_io_btb_resp_bridx = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_bridx : core_ibuf_io_imem_bits_btb_bridx ; 
  assign  core_ibuf_io_btb_resp_target = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_target : core_ibuf_io_imem_bits_btb_target ; 
  assign  core_ibuf_io_btb_resp_entry = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_entry : core_ibuf_io_imem_bits_btb_entry ; 
  assign  core_ibuf_io_btb_resp_bht_history = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_bht_history : core_ibuf_io_imem_bits_btb_bht_history ; 
  assign  core_ibuf_io_btb_resp_bht_value = core_ibuf__GEN_27  ?  core_ibuf_ibufBTBResp_bht_value : core_ibuf_io_imem_bits_btb_bht_value ; 
  assign  core_ibuf_io_inst_0_valid = core_ibuf_valid [0]& core_ibuf_full_insn ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_pf_inst = core_ibuf_xcpt_0_pf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_gf_inst = core_ibuf_xcpt_0_gf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt0_ae_inst = core_ibuf_xcpt_0_ae_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_pf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_pf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_gf_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_gf_inst ; 
  assign  core_ibuf_io_inst_0_bits_xcpt1_ae_inst = core_ibuf__io_inst_0_bits_xcpt1_WIRE_ae_inst ; 
  assign  core_ibuf_io_inst_0_bits_replay = core_ibuf_replay ; 
  assign  core_ibuf_io_inst_0_bits_rvc = core_ibuf__exp_io_rvc ; 
  assign  core_ibuf_io_inst_0_bits_raw = core_ibuf_inst ;
    assign core_ibuf_clock = core_clock;
    assign core_ibuf_reset = core_reset;
    assign core_io_imem_resp_ready = core_ibuf_io_imem_ready;
    assign core_ibuf_io_imem_valid = core_io_imem_resp_valid;
    assign core_ibuf_io_imem_bits_btb_cfiType = core_io_imem_resp_bits_btb_cfiType;
    assign core_ibuf_io_imem_bits_btb_taken = core_io_imem_resp_bits_btb_taken;
    assign core_ibuf_io_imem_bits_btb_mask = core_io_imem_resp_bits_btb_mask;
    assign core_ibuf_io_imem_bits_btb_bridx = core_io_imem_resp_bits_btb_bridx;
    assign core_ibuf_io_imem_bits_btb_target = core_io_imem_resp_bits_btb_target;
    assign core_ibuf_io_imem_bits_btb_entry = core_io_imem_resp_bits_btb_entry;
    assign core_ibuf_io_imem_bits_btb_bht_history = core_io_imem_resp_bits_btb_bht_history;
    assign core_ibuf_io_imem_bits_btb_bht_value = core_io_imem_resp_bits_btb_bht_value;
    assign core_ibuf_io_imem_bits_pc = core_io_imem_resp_bits_pc;
    assign core_ibuf_io_imem_bits_data = core_io_imem_resp_bits_data;
    assign core_ibuf_io_imem_bits_mask = core_io_imem_resp_bits_mask;
    assign core_ibuf_io_imem_bits_xcpt_pf_inst = core_io_imem_resp_bits_xcpt_pf_inst;
    assign core_ibuf_io_imem_bits_xcpt_gf_inst = core_io_imem_resp_bits_xcpt_gf_inst;
    assign core_ibuf_io_imem_bits_xcpt_ae_inst = core_io_imem_resp_bits_xcpt_ae_inst;
    assign core_ibuf_io_imem_bits_replay = core_io_imem_resp_bits_replay;
    assign core_ibuf_io_kill = core_take_pc_mem_wb;
    assign core__ibuf_io_pc = core_ibuf_io_pc;
    assign core__ibuf_io_btb_resp_cfiType = core_ibuf_io_btb_resp_cfiType;
    assign core__ibuf_io_btb_resp_taken = core_ibuf_io_btb_resp_taken;
    assign core__ibuf_io_btb_resp_mask = core_ibuf_io_btb_resp_mask;
    assign core__ibuf_io_btb_resp_bridx = core_ibuf_io_btb_resp_bridx;
    assign core__ibuf_io_btb_resp_target = core_ibuf_io_btb_resp_target;
    assign core__ibuf_io_btb_resp_entry = core_ibuf_io_btb_resp_entry;
    assign core__ibuf_io_btb_resp_bht_history = core_ibuf_io_btb_resp_bht_history;
    assign core__ibuf_io_btb_resp_bht_value = core_ibuf_io_btb_resp_bht_value;
    assign core_ibuf_io_inst_0_ready = core__GEN;
    assign core__ibuf_io_inst_0_valid = core_ibuf_io_inst_0_valid;
    assign core__ibuf_io_inst_0_bits_xcpt0_pf_inst = core_ibuf_io_inst_0_bits_xcpt0_pf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt0_gf_inst = core_ibuf_io_inst_0_bits_xcpt0_gf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt0_ae_inst = core_ibuf_io_inst_0_bits_xcpt0_ae_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_pf_inst = core_ibuf_io_inst_0_bits_xcpt1_pf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_gf_inst = core_ibuf_io_inst_0_bits_xcpt1_gf_inst;
    assign core__ibuf_io_inst_0_bits_xcpt1_ae_inst = core_ibuf_io_inst_0_bits_xcpt1_ae_inst;
    assign core__ibuf_io_inst_0_bits_replay = core_ibuf_io_inst_0_bits_replay;
    assign core__ibuf_io_inst_0_bits_rvc = core_ibuf_io_inst_0_bits_rvc;
    assign core__ibuf_io_inst_0_bits_inst_bits = core_ibuf_io_inst_0_bits_inst_bits;
    assign core_id_waddr = core_ibuf_io_inst_0_bits_inst_rd;
    assign core__ibuf_io_inst_0_bits_inst_rs1 = core_ibuf_io_inst_0_bits_inst_rs1;
    assign core_id_raddr2 = core_ibuf_io_inst_0_bits_inst_rs2;
    assign core_id_raddr3 = core_ibuf_io_inst_0_bits_inst_rs3;
    assign core__ibuf_io_inst_0_bits_raw = core_ibuf_io_inst_0_bits_raw;
     
    wire[31:0] core_id_ctrl_decoder_decoded_plaInput ; 
  assign  core_id_ctrl_decoder_decoded_plaInput = core__ibuf_io_inst_0_bits_inst_bits ; 
    wire core_id_ctrl_decoder_0 ; 
    wire[4:0] core_id_raddr1 ; 
  assign  core_id_raddr1 = core__ibuf_io_inst_0_bits_inst_rs1 ; 
    wire core_id_ctrl_decoder_1 ; 
    wire core_id_ctrl_decoder_2 ; 
    wire core_id_ctrl_decoder_3 ; 
    wire core_id_ctrl_decoder_4 ; 
    wire core_id_ctrl_decoder_5 ; 
    wire core_id_ctrl_decoder_6 ; 
    wire core_id_ctrl_decoder_7 ; 
    wire[1:0] core_id_ctrl_decoder_8 ; 
    wire[1:0] core_id_ctrl_decoder_9 ; 
    wire[2:0] core_id_ctrl_decoder_10 ; 
    wire core_id_ctrl_decoder_11 ; 
    wire[3:0] core_id_ctrl_decoder_12 ; 
    wire core_id_ctrl_decoder_13 ; 
    wire[4:0] core_id_ctrl_decoder_14 ; 
    wire core_id_ctrl_decoder_15 ; 
    wire core_id_ctrl_decoder_16 ; 
    wire core_id_ctrl_decoder_17 ; 
    wire core_id_ctrl_decoder_18 ; 
    wire core_id_ctrl_decoder_19 ; 
    wire core_id_ctrl_decoder_20 ; 
    wire core_id_ctrl_decoder_21 ; 
    wire[2:0] core_id_ctrl_decoder_22 ; 
    wire core_id_ctrl_decoder_23 ; 
    wire core_id_ctrl_decoder_24 ; 
    wire core_id_ctrl_decoder_25 ; 
    wire core_id_ctrl_decoder_26 ; 
    wire[31:0] core_id_ctrl_decoder_decoded_invInputs =~ core_id_ctrl_decoder_decoded_plaInput ; 
    wire[39:0] core_id_ctrl_decoder_decoded_invMatrixOutputs ; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4 , core_id_ctrl_decoder_decoded_andMatrixInput_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo ={ core_id_ctrl_decoder_decoded_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2 , core_id_ctrl_decoder_decoded_andMatrixInput_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0 , core_id_ctrl_decoder_decoded_andMatrixInput_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi ={ core_id_ctrl_decoder_decoded_hi_hi , core_id_ctrl_decoder_decoded_hi_lo }; 
    wire core__GEN_13 =&{ core_id_ctrl_decoder_decoded_hi , core_id_ctrl_decoder_decoded_lo }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_1 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_1 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_1 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_1 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_1 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_1 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_1 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_1 , core_id_ctrl_decoder_decoded_andMatrixInput_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_1 , core_id_ctrl_decoder_decoded_andMatrixInput_5_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_1 ={ core_id_ctrl_decoder_decoded_lo_hi_1 , core_id_ctrl_decoder_decoded_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_1 , core_id_ctrl_decoder_decoded_andMatrixInput_3_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_1 , core_id_ctrl_decoder_decoded_andMatrixInput_1_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_1 ={ core_id_ctrl_decoder_decoded_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_1 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_2 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_2 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_2 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_2 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_2 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_2 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_2 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_1 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_2 , core_id_ctrl_decoder_decoded_andMatrixInput_7_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_2 , core_id_ctrl_decoder_decoded_andMatrixInput_5_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_2 ={ core_id_ctrl_decoder_decoded_lo_hi_2 , core_id_ctrl_decoder_decoded_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_2 , core_id_ctrl_decoder_decoded_andMatrixInput_3_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_2 , core_id_ctrl_decoder_decoded_andMatrixInput_1_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_2 ={ core_id_ctrl_decoder_decoded_hi_hi_2 , core_id_ctrl_decoder_decoded_hi_lo_2 }; 
    wire core__GEN_14 =&{ core_id_ctrl_decoder_decoded_hi_2 , core_id_ctrl_decoder_decoded_lo_2 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_3 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_3 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_3 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_3 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_3 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_3 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_3 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_3 , core_id_ctrl_decoder_decoded_andMatrixInput_5_3 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_3 ={ core_id_ctrl_decoder_decoded_lo_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_6_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_3 , core_id_ctrl_decoder_decoded_andMatrixInput_3_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_3 , core_id_ctrl_decoder_decoded_andMatrixInput_1_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_3 ={ core_id_ctrl_decoder_decoded_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_3 }; 
    wire core__GEN_15 =&{ core_id_ctrl_decoder_decoded_hi_3 , core_id_ctrl_decoder_decoded_lo_3 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_4 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_4 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_4 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_4 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_4 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_4 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_4 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_4 , core_id_ctrl_decoder_decoded_andMatrixInput_7_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_4 , core_id_ctrl_decoder_decoded_andMatrixInput_5_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_4 ={ core_id_ctrl_decoder_decoded_lo_hi_4 , core_id_ctrl_decoder_decoded_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_4 , core_id_ctrl_decoder_decoded_andMatrixInput_3_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_4 , core_id_ctrl_decoder_decoded_andMatrixInput_1_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_4 ={ core_id_ctrl_decoder_decoded_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_4 }; 
    wire core__GEN_16 =&{ core_id_ctrl_decoder_decoded_hi_4 , core_id_ctrl_decoder_decoded_lo_4 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_5 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_5 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_5 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_5 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_5 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_5 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_5 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_3 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_3 , core_id_ctrl_decoder_decoded_andMatrixInput_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_5 , core_id_ctrl_decoder_decoded_andMatrixInput_6_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_5 ={ core_id_ctrl_decoder_decoded_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_5 , core_id_ctrl_decoder_decoded_andMatrixInput_4_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_5 , core_id_ctrl_decoder_decoded_andMatrixInput_1_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_5 ={ core_id_ctrl_decoder_decoded_hi_hi_hi , core_id_ctrl_decoder_decoded_andMatrixInput_2_5 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_5 ={ core_id_ctrl_decoder_decoded_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_5 }; 
    wire core__GEN_17 =&{ core_id_ctrl_decoder_decoded_hi_5 , core_id_ctrl_decoder_decoded_lo_5 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_6 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_6 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_6 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_6 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_6 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_6 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_6 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_4 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_1 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_4 , core_id_ctrl_decoder_decoded_andMatrixInput_8_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_6 , core_id_ctrl_decoder_decoded_andMatrixInput_6_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_6 ={ core_id_ctrl_decoder_decoded_lo_hi_6 , core_id_ctrl_decoder_decoded_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_6 , core_id_ctrl_decoder_decoded_andMatrixInput_4_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_6 , core_id_ctrl_decoder_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_6 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_2_6 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_6 ={ core_id_ctrl_decoder_decoded_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_lo_6 }; 
    wire core__GEN_18 =&{ core_id_ctrl_decoder_decoded_hi_6 , core_id_ctrl_decoder_decoded_lo_6 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_7 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_7 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_7 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_7 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_7 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_7 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_7 , core_id_ctrl_decoder_decoded_andMatrixInput_4_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_7 ={ core_id_ctrl_decoder_decoded_lo_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_5_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_7 , core_id_ctrl_decoder_decoded_andMatrixInput_1_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_7 ={ core_id_ctrl_decoder_decoded_hi_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_2_7 }; 
    wire core__GEN_19 =&{ core_id_ctrl_decoder_decoded_hi_7 , core_id_ctrl_decoder_decoded_lo_7 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_8 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_8 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_8 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_8 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_8 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_8 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_7 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_8 , core_id_ctrl_decoder_decoded_andMatrixInput_5_8 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_8 ={ core_id_ctrl_decoder_decoded_lo_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_6_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_8 , core_id_ctrl_decoder_decoded_andMatrixInput_3_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_8 , core_id_ctrl_decoder_decoded_andMatrixInput_1_8 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_8 ={ core_id_ctrl_decoder_decoded_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_7 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_9 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_9 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_9 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_9 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_9 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_9 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_8 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_8 , core_id_ctrl_decoder_decoded_andMatrixInput_7_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_9 , core_id_ctrl_decoder_decoded_andMatrixInput_5_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_9 ={ core_id_ctrl_decoder_decoded_lo_hi_9 , core_id_ctrl_decoder_decoded_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_9 , core_id_ctrl_decoder_decoded_andMatrixInput_3_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_9 , core_id_ctrl_decoder_decoded_andMatrixInput_1_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_9 ={ core_id_ctrl_decoder_decoded_hi_hi_9 , core_id_ctrl_decoder_decoded_hi_lo_8 }; 
    wire core__GEN_20 =&{ core_id_ctrl_decoder_decoded_hi_9 , core_id_ctrl_decoder_decoded_lo_9 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_10 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_10 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_10 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_10 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_10 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_10 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_9 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_6 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_9 , core_id_ctrl_decoder_decoded_andMatrixInput_7_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_10 , core_id_ctrl_decoder_decoded_andMatrixInput_5_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_10 ={ core_id_ctrl_decoder_decoded_lo_hi_10 , core_id_ctrl_decoder_decoded_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_10 , core_id_ctrl_decoder_decoded_andMatrixInput_3_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_10 , core_id_ctrl_decoder_decoded_andMatrixInput_1_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_10 ={ core_id_ctrl_decoder_decoded_hi_hi_10 , core_id_ctrl_decoder_decoded_hi_lo_9 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_11 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_11 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_11 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_11 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_11 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_11 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_10 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_7 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_2 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_12 , core_id_ctrl_decoder_decoded_andMatrixInput_13 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_7 ={ core_id_ctrl_decoder_decoded_lo_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_10 , core_id_ctrl_decoder_decoded_andMatrixInput_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_2 , core_id_ctrl_decoder_decoded_andMatrixInput_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_11 ={ core_id_ctrl_decoder_decoded_lo_hi_hi , core_id_ctrl_decoder_decoded_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_11 ={ core_id_ctrl_decoder_decoded_lo_hi_11 , core_id_ctrl_decoder_decoded_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_10 , core_id_ctrl_decoder_decoded_andMatrixInput_7_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_11 , core_id_ctrl_decoder_decoded_andMatrixInput_5_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_10 ={ core_id_ctrl_decoder_decoded_hi_lo_hi , core_id_ctrl_decoder_decoded_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_11 , core_id_ctrl_decoder_decoded_andMatrixInput_3_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_11 , core_id_ctrl_decoder_decoded_andMatrixInput_1_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_11 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_hi_hi_lo }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_11 ={ core_id_ctrl_decoder_decoded_hi_hi_11 , core_id_ctrl_decoder_decoded_hi_lo_10 }; 
    wire core__GEN_21 =&{ core_id_ctrl_decoder_decoded_hi_11 , core_id_ctrl_decoder_decoded_lo_11 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_12 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_12 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_12 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_12 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_12 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_12 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_11 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_8 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_3 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_1 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_1 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_1 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_1 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_1 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_1 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_1 , core_id_ctrl_decoder_decoded_andMatrixInput_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_1 , core_id_ctrl_decoder_decoded_andMatrixInput_13_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_8 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_1 , core_id_ctrl_decoder_decoded_andMatrixInput_11_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_3 , core_id_ctrl_decoder_decoded_andMatrixInput_9_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_12 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_lo_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_12 ={ core_id_ctrl_decoder_decoded_lo_hi_12 , core_id_ctrl_decoder_decoded_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_11 , core_id_ctrl_decoder_decoded_andMatrixInput_7_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_12 , core_id_ctrl_decoder_decoded_andMatrixInput_5_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_11 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_12 , core_id_ctrl_decoder_decoded_andMatrixInput_3_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_12 , core_id_ctrl_decoder_decoded_andMatrixInput_1_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_12 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_12 ={ core_id_ctrl_decoder_decoded_hi_hi_12 , core_id_ctrl_decoder_decoded_hi_lo_11 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_13 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_13 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_13 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_13 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_13 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_13 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_12 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_9 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_2 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_2 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_2 , core_id_ctrl_decoder_decoded_andMatrixInput_11_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_9 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_12_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_9 , core_id_ctrl_decoder_decoded_andMatrixInput_8_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_13 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_9_2 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_13 ={ core_id_ctrl_decoder_decoded_lo_hi_13 , core_id_ctrl_decoder_decoded_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_13 , core_id_ctrl_decoder_decoded_andMatrixInput_5_13 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_12 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_6_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_13 , core_id_ctrl_decoder_decoded_andMatrixInput_3_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_13 , core_id_ctrl_decoder_decoded_andMatrixInput_1_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_13 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_13 ={ core_id_ctrl_decoder_decoded_hi_hi_13 , core_id_ctrl_decoder_decoded_hi_lo_12 }; 
    wire core__GEN_22 =&{ core_id_ctrl_decoder_decoded_hi_13 , core_id_ctrl_decoder_decoded_lo_13 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_14 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_14 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_14 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_14 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_14 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_14 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_13 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_10 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_3 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_3 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_3 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_3 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_3 , core_id_ctrl_decoder_decoded_andMatrixInput_13_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_10 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_14_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_3 , core_id_ctrl_decoder_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_5 , core_id_ctrl_decoder_decoded_andMatrixInput_9_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_14 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_14 ={ core_id_ctrl_decoder_decoded_lo_hi_14 , core_id_ctrl_decoder_decoded_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_13 , core_id_ctrl_decoder_decoded_andMatrixInput_7_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_14 , core_id_ctrl_decoder_decoded_andMatrixInput_5_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_13 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_14 , core_id_ctrl_decoder_decoded_andMatrixInput_3_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_14 , core_id_ctrl_decoder_decoded_andMatrixInput_1_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_14 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_14 ={ core_id_ctrl_decoder_decoded_hi_hi_14 , core_id_ctrl_decoder_decoded_hi_lo_13 }; 
    wire core__GEN_23 =&{ core_id_ctrl_decoder_decoded_hi_14 , core_id_ctrl_decoder_decoded_lo_14 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_15 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_15 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_15 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_15 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_15 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_15 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_14 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_11 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_6 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_4 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_4 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_4 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_3 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_3 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_4 , core_id_ctrl_decoder_decoded_andMatrixInput_13_3 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_11 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_14_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_4 , core_id_ctrl_decoder_decoded_andMatrixInput_11_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_6 , core_id_ctrl_decoder_decoded_andMatrixInput_9_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_15 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_15 ={ core_id_ctrl_decoder_decoded_lo_hi_15 , core_id_ctrl_decoder_decoded_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_14 , core_id_ctrl_decoder_decoded_andMatrixInput_7_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_15 , core_id_ctrl_decoder_decoded_andMatrixInput_5_15 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_14 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_15 , core_id_ctrl_decoder_decoded_andMatrixInput_3_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_15 , core_id_ctrl_decoder_decoded_andMatrixInput_1_15 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_15 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_hi_lo_4 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_15 ={ core_id_ctrl_decoder_decoded_hi_hi_15 , core_id_ctrl_decoder_decoded_hi_lo_14 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_16 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_16 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_16 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_16 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_16 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_16 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_15 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_12 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_15 , core_id_ctrl_decoder_decoded_andMatrixInput_7_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_16 , core_id_ctrl_decoder_decoded_andMatrixInput_5_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_16 ={ core_id_ctrl_decoder_decoded_lo_hi_16 , core_id_ctrl_decoder_decoded_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_16 , core_id_ctrl_decoder_decoded_andMatrixInput_3_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_16 , core_id_ctrl_decoder_decoded_andMatrixInput_1_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_16 ={ core_id_ctrl_decoder_decoded_hi_hi_16 , core_id_ctrl_decoder_decoded_hi_lo_15 }; 
    wire core__GEN_24 =&{ core_id_ctrl_decoder_decoded_hi_16 , core_id_ctrl_decoder_decoded_lo_16 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_17 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_17 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_17 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_17 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_17 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_17 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_16 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_13 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_7 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_13 , core_id_ctrl_decoder_decoded_andMatrixInput_8_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_17 , core_id_ctrl_decoder_decoded_andMatrixInput_6_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_17 ={ core_id_ctrl_decoder_decoded_lo_hi_17 , core_id_ctrl_decoder_decoded_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_17 , core_id_ctrl_decoder_decoded_andMatrixInput_4_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_17 , core_id_ctrl_decoder_decoded_andMatrixInput_1_17 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_17 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_2_17 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_17 ={ core_id_ctrl_decoder_decoded_hi_hi_17 , core_id_ctrl_decoder_decoded_hi_lo_16 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_18 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_18 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_18 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_18 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_18 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_18 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_17 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_14 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_8 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_14 , core_id_ctrl_decoder_decoded_andMatrixInput_8_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_18 , core_id_ctrl_decoder_decoded_andMatrixInput_6_17 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_18 ={ core_id_ctrl_decoder_decoded_lo_hi_18 , core_id_ctrl_decoder_decoded_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_18 , core_id_ctrl_decoder_decoded_andMatrixInput_4_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_18 , core_id_ctrl_decoder_decoded_andMatrixInput_1_18 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_18 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_2_18 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_18 ={ core_id_ctrl_decoder_decoded_hi_hi_18 , core_id_ctrl_decoder_decoded_hi_lo_17 }; 
    wire core__GEN_25 =&{ core_id_ctrl_decoder_decoded_hi_18 , core_id_ctrl_decoder_decoded_lo_18 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_19 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_19 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_19 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_19 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_19 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_19 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_18 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_15 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_9 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_9 , core_id_ctrl_decoder_decoded_andMatrixInput_9_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_19 , core_id_ctrl_decoder_decoded_andMatrixInput_6_18 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_19 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_andMatrixInput_7_15 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_19 ={ core_id_ctrl_decoder_decoded_lo_hi_19 , core_id_ctrl_decoder_decoded_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_19 , core_id_ctrl_decoder_decoded_andMatrixInput_4_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_19 , core_id_ctrl_decoder_decoded_andMatrixInput_1_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_19 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_9 , core_id_ctrl_decoder_decoded_andMatrixInput_2_19 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_19 ={ core_id_ctrl_decoder_decoded_hi_hi_19 , core_id_ctrl_decoder_decoded_hi_lo_18 }; 
    wire core__GEN_26 =&{ core_id_ctrl_decoder_decoded_hi_19 , core_id_ctrl_decoder_decoded_lo_19 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_20 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_20 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_20 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_20 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_20 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_20 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_19 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_20 , core_id_ctrl_decoder_decoded_andMatrixInput_5_20 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_20 ={ core_id_ctrl_decoder_decoded_lo_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_6_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_20 , core_id_ctrl_decoder_decoded_andMatrixInput_3_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_20 , core_id_ctrl_decoder_decoded_andMatrixInput_1_20 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_20 ={ core_id_ctrl_decoder_decoded_hi_hi_20 , core_id_ctrl_decoder_decoded_hi_lo_19 }; 
    wire core__GEN_27 =&{ core_id_ctrl_decoder_decoded_hi_20 , core_id_ctrl_decoder_decoded_lo_20 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_21 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_21 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_21 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_21 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_21 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_21 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_20 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_16 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_10 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_6 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_5 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_5 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_4 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_4 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_1 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_25 , core_id_ctrl_decoder_decoded_andMatrixInput_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_23 , core_id_ctrl_decoder_decoded_andMatrixInput_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_21 , core_id_ctrl_decoder_decoded_andMatrixInput_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_lo_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_16 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_18 , core_id_ctrl_decoder_decoded_andMatrixInput_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_16 , core_id_ctrl_decoder_decoded_andMatrixInput_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_4 , core_id_ctrl_decoder_decoded_andMatrixInput_15_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_lo_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_21 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_hi_lo_4 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_21 ={ core_id_ctrl_decoder_decoded_lo_hi_21 , core_id_ctrl_decoder_decoded_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_5 , core_id_ctrl_decoder_decoded_andMatrixInput_12_5 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_4 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_13_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_6 , core_id_ctrl_decoder_decoded_andMatrixInput_10_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_16 , core_id_ctrl_decoder_decoded_andMatrixInput_8_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_hi_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_20 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_21 , core_id_ctrl_decoder_decoded_andMatrixInput_5_21 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi , core_id_ctrl_decoder_decoded_andMatrixInput_6_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_21 , core_id_ctrl_decoder_decoded_andMatrixInput_3_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_21 , core_id_ctrl_decoder_decoded_andMatrixInput_1_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_10 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_hi_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_21 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_10 , core_id_ctrl_decoder_decoded_hi_hi_lo_5 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_21 ={ core_id_ctrl_decoder_decoded_hi_hi_21 , core_id_ctrl_decoder_decoded_hi_lo_20 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_22 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_22 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_22 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_22 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_22 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_22 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_21 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_17 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_11 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_7 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_6 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_6 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_6 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_5 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_5 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_2 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_1 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_1 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_1 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_1 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_1 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_1 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_1 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_1 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_1 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_1 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_1 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_1 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28 , core_id_ctrl_decoder_decoded_andMatrixInput_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_2 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_andMatrixInput_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_1 , core_id_ctrl_decoder_decoded_andMatrixInput_27_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_1 , core_id_ctrl_decoder_decoded_andMatrixInput_25_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_1 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_17 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_lo_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_1 , core_id_ctrl_decoder_decoded_andMatrixInput_23_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_1 , core_id_ctrl_decoder_decoded_andMatrixInput_21_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_1 , core_id_ctrl_decoder_decoded_andMatrixInput_19_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_1 , core_id_ctrl_decoder_decoded_andMatrixInput_17_1 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_22 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_lo_5 }; 
    wire[14:0] core_id_ctrl_decoder_decoded_lo_22 ={ core_id_ctrl_decoder_decoded_lo_hi_22 , core_id_ctrl_decoder_decoded_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_5 , core_id_ctrl_decoder_decoded_andMatrixInput_15_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_6 , core_id_ctrl_decoder_decoded_andMatrixInput_13_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_5 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_6 , core_id_ctrl_decoder_decoded_andMatrixInput_11_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_11 , core_id_ctrl_decoder_decoded_andMatrixInput_9_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_21 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_hi_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_21 , core_id_ctrl_decoder_decoded_andMatrixInput_7_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_22 , core_id_ctrl_decoder_decoded_andMatrixInput_5_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_1 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_22 , core_id_ctrl_decoder_decoded_andMatrixInput_3_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_22 , core_id_ctrl_decoder_decoded_andMatrixInput_1_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_11 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_1 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_1 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_22 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_11 , core_id_ctrl_decoder_decoded_hi_hi_lo_6 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_22 ={ core_id_ctrl_decoder_decoded_hi_hi_22 , core_id_ctrl_decoder_decoded_hi_lo_21 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_23 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_23 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_23 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_23 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_23 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_23 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_22 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_18 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_12 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_8 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_12 , core_id_ctrl_decoder_decoded_andMatrixInput_9_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_23 , core_id_ctrl_decoder_decoded_andMatrixInput_6_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_23 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_7_18 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_23 ={ core_id_ctrl_decoder_decoded_lo_hi_23 , core_id_ctrl_decoder_decoded_lo_lo_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_23 , core_id_ctrl_decoder_decoded_andMatrixInput_4_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_23 , core_id_ctrl_decoder_decoded_andMatrixInput_1_23 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_23 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_12 , core_id_ctrl_decoder_decoded_andMatrixInput_2_23 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_23 ={ core_id_ctrl_decoder_decoded_hi_hi_23 , core_id_ctrl_decoder_decoded_hi_lo_22 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_24 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_24 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_24 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_24 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_24 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_24 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_23 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_19 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_13 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_9 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_7 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_7 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_7 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_7 , core_id_ctrl_decoder_decoded_andMatrixInput_12_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_19 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_13_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_9 , core_id_ctrl_decoder_decoded_andMatrixInput_10_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_19 , core_id_ctrl_decoder_decoded_andMatrixInput_8_13 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_24 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_9 , core_id_ctrl_decoder_decoded_lo_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_24 ={ core_id_ctrl_decoder_decoded_lo_hi_24 , core_id_ctrl_decoder_decoded_lo_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_24 , core_id_ctrl_decoder_decoded_andMatrixInput_5_24 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_23 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_andMatrixInput_6_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_24 , core_id_ctrl_decoder_decoded_andMatrixInput_3_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_24 , core_id_ctrl_decoder_decoded_andMatrixInput_1_24 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_24 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_13 , core_id_ctrl_decoder_decoded_hi_hi_lo_7 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_24 ={ core_id_ctrl_decoder_decoded_hi_hi_24 , core_id_ctrl_decoder_decoded_hi_lo_23 }; 
    wire core__GEN_28 =&{ core_id_ctrl_decoder_decoded_hi_24 , core_id_ctrl_decoder_decoded_lo_24 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_25 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_25 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_25 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_25 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_25 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_25 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_24 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_20 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_14 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_10 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_8 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_8 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_8 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_7 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_8 , core_id_ctrl_decoder_decoded_andMatrixInput_13_7 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_20 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_8 , core_id_ctrl_decoder_decoded_andMatrixInput_14_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_8 , core_id_ctrl_decoder_decoded_andMatrixInput_11_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_14 , core_id_ctrl_decoder_decoded_andMatrixInput_9_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_25 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_10 , core_id_ctrl_decoder_decoded_lo_hi_lo_7 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_25 ={ core_id_ctrl_decoder_decoded_lo_hi_25 , core_id_ctrl_decoder_decoded_lo_lo_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_24 , core_id_ctrl_decoder_decoded_andMatrixInput_7_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_25 , core_id_ctrl_decoder_decoded_andMatrixInput_5_25 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_24 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_25 , core_id_ctrl_decoder_decoded_andMatrixInput_3_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_25 , core_id_ctrl_decoder_decoded_andMatrixInput_1_25 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_25 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_14 , core_id_ctrl_decoder_decoded_hi_hi_lo_8 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_25 ={ core_id_ctrl_decoder_decoded_hi_hi_25 , core_id_ctrl_decoder_decoded_hi_lo_24 }; 
    wire core__GEN_29 =&{ core_id_ctrl_decoder_decoded_hi_25 , core_id_ctrl_decoder_decoded_lo_25 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_26 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_26 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_26 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_26 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_26 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_26 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_25 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_21 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_15 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_11 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_9 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_9 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_9 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_8 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_7 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_9 , core_id_ctrl_decoder_decoded_andMatrixInput_13_8 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_21 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_9 , core_id_ctrl_decoder_decoded_andMatrixInput_14_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_9 , core_id_ctrl_decoder_decoded_andMatrixInput_11_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_15 , core_id_ctrl_decoder_decoded_andMatrixInput_9_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_26 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_11 , core_id_ctrl_decoder_decoded_lo_hi_lo_8 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_26 ={ core_id_ctrl_decoder_decoded_lo_hi_26 , core_id_ctrl_decoder_decoded_lo_lo_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_25 , core_id_ctrl_decoder_decoded_andMatrixInput_7_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_26 , core_id_ctrl_decoder_decoded_andMatrixInput_5_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_25 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_9 , core_id_ctrl_decoder_decoded_hi_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_26 , core_id_ctrl_decoder_decoded_andMatrixInput_3_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_26 , core_id_ctrl_decoder_decoded_andMatrixInput_1_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_26 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_15 , core_id_ctrl_decoder_decoded_hi_hi_lo_9 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_26 ={ core_id_ctrl_decoder_decoded_hi_hi_26 , core_id_ctrl_decoder_decoded_hi_lo_25 }; 
    wire core__GEN_30 =&{ core_id_ctrl_decoder_decoded_hi_26 , core_id_ctrl_decoder_decoded_lo_26 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_27 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_27 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_27 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_27 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_27 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_27 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_26 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_22 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_16 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_12 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_10 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_10 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_10 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_9 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_8 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_3 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_8 , core_id_ctrl_decoder_decoded_andMatrixInput_15_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_10 , core_id_ctrl_decoder_decoded_andMatrixInput_13_9 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_22 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_10 , core_id_ctrl_decoder_decoded_lo_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_10 , core_id_ctrl_decoder_decoded_andMatrixInput_11_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_16 , core_id_ctrl_decoder_decoded_andMatrixInput_9_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_27 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_12 , core_id_ctrl_decoder_decoded_lo_hi_lo_9 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_27 ={ core_id_ctrl_decoder_decoded_lo_hi_27 , core_id_ctrl_decoder_decoded_lo_lo_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_26 , core_id_ctrl_decoder_decoded_andMatrixInput_7_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_27 , core_id_ctrl_decoder_decoded_andMatrixInput_5_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_26 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_10 , core_id_ctrl_decoder_decoded_hi_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_27 , core_id_ctrl_decoder_decoded_andMatrixInput_3_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_27 , core_id_ctrl_decoder_decoded_andMatrixInput_1_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_27 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_16 , core_id_ctrl_decoder_decoded_hi_hi_lo_10 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_27 ={ core_id_ctrl_decoder_decoded_hi_hi_27 , core_id_ctrl_decoder_decoded_hi_lo_26 }; 
    wire core__GEN_31 =&{ core_id_ctrl_decoder_decoded_hi_27 , core_id_ctrl_decoder_decoded_lo_27 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_28 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_28 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_28 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_28 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_28 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_28 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_27 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_23 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_27 , core_id_ctrl_decoder_decoded_andMatrixInput_7_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_28 , core_id_ctrl_decoder_decoded_andMatrixInput_5_28 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_28 ={ core_id_ctrl_decoder_decoded_lo_hi_28 , core_id_ctrl_decoder_decoded_lo_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_28 , core_id_ctrl_decoder_decoded_andMatrixInput_3_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_28 , core_id_ctrl_decoder_decoded_andMatrixInput_1_28 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_28 ={ core_id_ctrl_decoder_decoded_hi_hi_28 , core_id_ctrl_decoder_decoded_hi_lo_27 }; 
    wire core__GEN_32 =&{ core_id_ctrl_decoder_decoded_hi_28 , core_id_ctrl_decoder_decoded_lo_28 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_29 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_29 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_29 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_29 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_29 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_29 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_28 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_24 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_17 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_24 , core_id_ctrl_decoder_decoded_andMatrixInput_8_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_29 , core_id_ctrl_decoder_decoded_andMatrixInput_6_28 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_29 ={ core_id_ctrl_decoder_decoded_lo_hi_29 , core_id_ctrl_decoder_decoded_lo_lo_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_29 , core_id_ctrl_decoder_decoded_andMatrixInput_4_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_29 , core_id_ctrl_decoder_decoded_andMatrixInput_1_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_29 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_17 , core_id_ctrl_decoder_decoded_andMatrixInput_2_29 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_29 ={ core_id_ctrl_decoder_decoded_hi_hi_29 , core_id_ctrl_decoder_decoded_hi_lo_28 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_30 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_30 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_30 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_30 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_30 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_30 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_29 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_25 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_18 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_25 , core_id_ctrl_decoder_decoded_andMatrixInput_8_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_30 , core_id_ctrl_decoder_decoded_andMatrixInput_6_29 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_30 ={ core_id_ctrl_decoder_decoded_lo_hi_30 , core_id_ctrl_decoder_decoded_lo_lo_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_30 , core_id_ctrl_decoder_decoded_andMatrixInput_4_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_30 , core_id_ctrl_decoder_decoded_andMatrixInput_1_30 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_30 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_18 , core_id_ctrl_decoder_decoded_andMatrixInput_2_30 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_30 ={ core_id_ctrl_decoder_decoded_hi_hi_30 , core_id_ctrl_decoder_decoded_hi_lo_29 }; 
    wire core__GEN_33 =&{ core_id_ctrl_decoder_decoded_hi_30 , core_id_ctrl_decoder_decoded_lo_30 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_31 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_31 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_31 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_31 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_31 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_31 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_30 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_26 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_30 , core_id_ctrl_decoder_decoded_andMatrixInput_7_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_31 , core_id_ctrl_decoder_decoded_andMatrixInput_5_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_31 ={ core_id_ctrl_decoder_decoded_lo_hi_31 , core_id_ctrl_decoder_decoded_lo_lo_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_31 , core_id_ctrl_decoder_decoded_andMatrixInput_3_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_31 , core_id_ctrl_decoder_decoded_andMatrixInput_1_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_31 ={ core_id_ctrl_decoder_decoded_hi_hi_31 , core_id_ctrl_decoder_decoded_hi_lo_30 }; 
    wire core__GEN_34 =&{ core_id_ctrl_decoder_decoded_hi_31 , core_id_ctrl_decoder_decoded_lo_31 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_32 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_32 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_32 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_32 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_32 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_32 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_31 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_27 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_31 , core_id_ctrl_decoder_decoded_andMatrixInput_7_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_32 , core_id_ctrl_decoder_decoded_andMatrixInput_5_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_32 ={ core_id_ctrl_decoder_decoded_lo_hi_32 , core_id_ctrl_decoder_decoded_lo_lo_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_32 , core_id_ctrl_decoder_decoded_andMatrixInput_3_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_32 , core_id_ctrl_decoder_decoded_andMatrixInput_1_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_32 ={ core_id_ctrl_decoder_decoded_hi_hi_32 , core_id_ctrl_decoder_decoded_hi_lo_31 }; 
    wire core__GEN_35 =&{ core_id_ctrl_decoder_decoded_hi_32 , core_id_ctrl_decoder_decoded_lo_32 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_33 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_33 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_33 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_33 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_33 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_33 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_32 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_28 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_19 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_28 , core_id_ctrl_decoder_decoded_andMatrixInput_8_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_33 , core_id_ctrl_decoder_decoded_andMatrixInput_6_32 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_33 ={ core_id_ctrl_decoder_decoded_lo_hi_33 , core_id_ctrl_decoder_decoded_lo_lo_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_33 , core_id_ctrl_decoder_decoded_andMatrixInput_4_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_33 , core_id_ctrl_decoder_decoded_andMatrixInput_1_33 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_33 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_19 , core_id_ctrl_decoder_decoded_andMatrixInput_2_33 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_33 ={ core_id_ctrl_decoder_decoded_hi_hi_33 , core_id_ctrl_decoder_decoded_hi_lo_32 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_34 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_34 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_34 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_34 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_34 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_34 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_33 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_29 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_20 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_13 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_11 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_13 , core_id_ctrl_decoder_decoded_andMatrixInput_10_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_33 , core_id_ctrl_decoder_decoded_andMatrixInput_7_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_34 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_13 , core_id_ctrl_decoder_decoded_andMatrixInput_8_20 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_34 ={ core_id_ctrl_decoder_decoded_lo_hi_34 , core_id_ctrl_decoder_decoded_lo_lo_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_34 , core_id_ctrl_decoder_decoded_andMatrixInput_4_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_33 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_11 , core_id_ctrl_decoder_decoded_andMatrixInput_5_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_34 , core_id_ctrl_decoder_decoded_andMatrixInput_1_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_34 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_2_34 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_hi_34 ={ core_id_ctrl_decoder_decoded_hi_hi_34 , core_id_ctrl_decoder_decoded_hi_lo_33 }; 
    wire core__GEN_36 =&{ core_id_ctrl_decoder_decoded_hi_34 , core_id_ctrl_decoder_decoded_lo_34 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_35 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_35 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_35 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_35 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_35 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_35 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_34 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_30 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_21 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_14 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_12 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_11 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_11 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_10 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_9 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_11 , core_id_ctrl_decoder_decoded_andMatrixInput_13_10 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_30 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_11 , core_id_ctrl_decoder_decoded_andMatrixInput_14_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_12 , core_id_ctrl_decoder_decoded_andMatrixInput_11_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_21 , core_id_ctrl_decoder_decoded_andMatrixInput_9_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_35 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_14 , core_id_ctrl_decoder_decoded_lo_hi_lo_10 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_35 ={ core_id_ctrl_decoder_decoded_lo_hi_35 , core_id_ctrl_decoder_decoded_lo_lo_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_34 , core_id_ctrl_decoder_decoded_andMatrixInput_7_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_35 , core_id_ctrl_decoder_decoded_andMatrixInput_5_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_34 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_12 , core_id_ctrl_decoder_decoded_hi_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_35 , core_id_ctrl_decoder_decoded_andMatrixInput_3_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_35 , core_id_ctrl_decoder_decoded_andMatrixInput_1_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_35 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_21 , core_id_ctrl_decoder_decoded_hi_hi_lo_11 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_35 ={ core_id_ctrl_decoder_decoded_hi_hi_35 , core_id_ctrl_decoder_decoded_hi_lo_34 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_36 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_36 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_36 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_36 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_36 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_36 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_35 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_31 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_22 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_15 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_13 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_12 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_12 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_11 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_10 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_4 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_10 , core_id_ctrl_decoder_decoded_andMatrixInput_15_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_12 , core_id_ctrl_decoder_decoded_andMatrixInput_13_11 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_31 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_12 , core_id_ctrl_decoder_decoded_lo_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_13 , core_id_ctrl_decoder_decoded_andMatrixInput_11_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_22 , core_id_ctrl_decoder_decoded_andMatrixInput_9_15 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_36 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_15 , core_id_ctrl_decoder_decoded_lo_hi_lo_11 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_36 ={ core_id_ctrl_decoder_decoded_lo_hi_36 , core_id_ctrl_decoder_decoded_lo_lo_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_10 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_35 , core_id_ctrl_decoder_decoded_andMatrixInput_7_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_36 , core_id_ctrl_decoder_decoded_andMatrixInput_5_36 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_35 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_13 , core_id_ctrl_decoder_decoded_hi_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_36 , core_id_ctrl_decoder_decoded_andMatrixInput_3_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_36 , core_id_ctrl_decoder_decoded_andMatrixInput_1_36 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_36 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_22 , core_id_ctrl_decoder_decoded_hi_hi_lo_12 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_36 ={ core_id_ctrl_decoder_decoded_hi_hi_36 , core_id_ctrl_decoder_decoded_hi_lo_35 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_37 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_37 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_37 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_37 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_37 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_37 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_36 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_32 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_36 , core_id_ctrl_decoder_decoded_andMatrixInput_7_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_37 , core_id_ctrl_decoder_decoded_andMatrixInput_5_37 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_37 ={ core_id_ctrl_decoder_decoded_lo_hi_37 , core_id_ctrl_decoder_decoded_lo_lo_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_37 , core_id_ctrl_decoder_decoded_andMatrixInput_3_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_37 , core_id_ctrl_decoder_decoded_andMatrixInput_1_37 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_37 ={ core_id_ctrl_decoder_decoded_hi_hi_37 , core_id_ctrl_decoder_decoded_hi_lo_36 }; 
    wire core__GEN_37 =&{ core_id_ctrl_decoder_decoded_hi_37 , core_id_ctrl_decoder_decoded_lo_37 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_38 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_38 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_38 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_38 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_38 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_38 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_37 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_33 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_23 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_33 , core_id_ctrl_decoder_decoded_andMatrixInput_8_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_38 , core_id_ctrl_decoder_decoded_andMatrixInput_6_37 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_38 ={ core_id_ctrl_decoder_decoded_lo_hi_38 , core_id_ctrl_decoder_decoded_lo_lo_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_38 , core_id_ctrl_decoder_decoded_andMatrixInput_4_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_38 , core_id_ctrl_decoder_decoded_andMatrixInput_1_38 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_38 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_23 , core_id_ctrl_decoder_decoded_andMatrixInput_2_38 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_38 ={ core_id_ctrl_decoder_decoded_hi_hi_38 , core_id_ctrl_decoder_decoded_hi_lo_37 }; 
    wire core__GEN_38 =&{ core_id_ctrl_decoder_decoded_hi_38 , core_id_ctrl_decoder_decoded_lo_38 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_39 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_39 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_39 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_39 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_39 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_39 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_38 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_34 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_24 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_34 , core_id_ctrl_decoder_decoded_andMatrixInput_8_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_39 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_39 , core_id_ctrl_decoder_decoded_andMatrixInput_6_38 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_39 ={ core_id_ctrl_decoder_decoded_lo_hi_39 , core_id_ctrl_decoder_decoded_lo_lo_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_39 , core_id_ctrl_decoder_decoded_andMatrixInput_4_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_39 , core_id_ctrl_decoder_decoded_andMatrixInput_1_39 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_39 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_24 , core_id_ctrl_decoder_decoded_andMatrixInput_2_39 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_39 ={ core_id_ctrl_decoder_decoded_hi_hi_39 , core_id_ctrl_decoder_decoded_hi_lo_38 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_40 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_40 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_40 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_40 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_40 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_40 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_39 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_35 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_25 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_16 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_14 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_13 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_13 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_12 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_11 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_13 , core_id_ctrl_decoder_decoded_andMatrixInput_13_12 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_35 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_13 , core_id_ctrl_decoder_decoded_andMatrixInput_14_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_14 , core_id_ctrl_decoder_decoded_andMatrixInput_11_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_25 , core_id_ctrl_decoder_decoded_andMatrixInput_9_16 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_40 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_16 , core_id_ctrl_decoder_decoded_lo_hi_lo_12 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_40 ={ core_id_ctrl_decoder_decoded_lo_hi_40 , core_id_ctrl_decoder_decoded_lo_lo_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_11 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_39 , core_id_ctrl_decoder_decoded_andMatrixInput_7_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_40 , core_id_ctrl_decoder_decoded_andMatrixInput_5_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_39 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_14 , core_id_ctrl_decoder_decoded_hi_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_40 , core_id_ctrl_decoder_decoded_andMatrixInput_3_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_40 , core_id_ctrl_decoder_decoded_andMatrixInput_1_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_40 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_25 , core_id_ctrl_decoder_decoded_hi_hi_lo_13 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_40 ={ core_id_ctrl_decoder_decoded_hi_hi_40 , core_id_ctrl_decoder_decoded_hi_lo_39 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_41 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_41 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_41 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_41 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_41 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_41 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_40 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_36 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_26 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_36 , core_id_ctrl_decoder_decoded_andMatrixInput_8_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_41 , core_id_ctrl_decoder_decoded_andMatrixInput_6_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_41 ={ core_id_ctrl_decoder_decoded_lo_hi_41 , core_id_ctrl_decoder_decoded_lo_lo_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_41 , core_id_ctrl_decoder_decoded_andMatrixInput_4_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_41 , core_id_ctrl_decoder_decoded_andMatrixInput_1_41 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_41 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_26 , core_id_ctrl_decoder_decoded_andMatrixInput_2_41 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_41 ={ core_id_ctrl_decoder_decoded_hi_hi_41 , core_id_ctrl_decoder_decoded_hi_lo_40 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_42 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_42 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_42 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_42 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_42 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_42 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_41 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_37 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_27 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_17 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_15 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_14 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_14 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_13 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_14 , core_id_ctrl_decoder_decoded_andMatrixInput_12_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_37 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_14 , core_id_ctrl_decoder_decoded_andMatrixInput_13_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_17 , core_id_ctrl_decoder_decoded_andMatrixInput_10_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_37 , core_id_ctrl_decoder_decoded_andMatrixInput_8_27 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_42 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_17 , core_id_ctrl_decoder_decoded_lo_hi_lo_13 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_42 ={ core_id_ctrl_decoder_decoded_lo_hi_42 , core_id_ctrl_decoder_decoded_lo_lo_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_42 , core_id_ctrl_decoder_decoded_andMatrixInput_5_42 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_41 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_15 , core_id_ctrl_decoder_decoded_andMatrixInput_6_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_42 , core_id_ctrl_decoder_decoded_andMatrixInput_3_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_42 , core_id_ctrl_decoder_decoded_andMatrixInput_1_42 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_42 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_27 , core_id_ctrl_decoder_decoded_hi_hi_lo_14 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_42 ={ core_id_ctrl_decoder_decoded_hi_hi_42 , core_id_ctrl_decoder_decoded_hi_lo_41 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_43 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_43 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_43 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_43 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_43 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_43 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_42 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_38 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_42 , core_id_ctrl_decoder_decoded_andMatrixInput_7_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_43 , core_id_ctrl_decoder_decoded_andMatrixInput_5_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_43 ={ core_id_ctrl_decoder_decoded_lo_hi_43 , core_id_ctrl_decoder_decoded_lo_lo_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_43 , core_id_ctrl_decoder_decoded_andMatrixInput_3_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_43 , core_id_ctrl_decoder_decoded_andMatrixInput_1_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_43 ={ core_id_ctrl_decoder_decoded_hi_hi_43 , core_id_ctrl_decoder_decoded_hi_lo_42 }; 
    wire core__GEN_39 =&{ core_id_ctrl_decoder_decoded_hi_43 , core_id_ctrl_decoder_decoded_lo_43 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_44 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_44 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_44 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_44 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_44 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_44 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_43 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_39 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_28 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_18 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_16 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_15 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_15 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_14 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_12 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_15 , core_id_ctrl_decoder_decoded_andMatrixInput_13_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_39 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_15 , core_id_ctrl_decoder_decoded_andMatrixInput_14_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_16 , core_id_ctrl_decoder_decoded_andMatrixInput_11_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_28 , core_id_ctrl_decoder_decoded_andMatrixInput_9_18 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_44 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_18 , core_id_ctrl_decoder_decoded_lo_hi_lo_14 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_44 ={ core_id_ctrl_decoder_decoded_lo_hi_44 , core_id_ctrl_decoder_decoded_lo_lo_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_12 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_43 , core_id_ctrl_decoder_decoded_andMatrixInput_7_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_44 , core_id_ctrl_decoder_decoded_andMatrixInput_5_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_43 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_16 , core_id_ctrl_decoder_decoded_hi_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_44 , core_id_ctrl_decoder_decoded_andMatrixInput_3_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_44 , core_id_ctrl_decoder_decoded_andMatrixInput_1_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_44 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_28 , core_id_ctrl_decoder_decoded_hi_hi_lo_15 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_44 ={ core_id_ctrl_decoder_decoded_hi_hi_44 , core_id_ctrl_decoder_decoded_hi_lo_43 }; 
    wire core__GEN_40 =&{ core_id_ctrl_decoder_decoded_hi_44 , core_id_ctrl_decoder_decoded_lo_44 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_45 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_45 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_45 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_45 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_45 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_45 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_44 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_40 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_29 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_19 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_17 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_16 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_16 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_15 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_13 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_16 , core_id_ctrl_decoder_decoded_andMatrixInput_13_15 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_40 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_16 , core_id_ctrl_decoder_decoded_andMatrixInput_14_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_17 , core_id_ctrl_decoder_decoded_andMatrixInput_11_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_29 , core_id_ctrl_decoder_decoded_andMatrixInput_9_19 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_45 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_19 , core_id_ctrl_decoder_decoded_lo_hi_lo_15 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_45 ={ core_id_ctrl_decoder_decoded_lo_hi_45 , core_id_ctrl_decoder_decoded_lo_lo_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_13 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_44 , core_id_ctrl_decoder_decoded_andMatrixInput_7_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_45 , core_id_ctrl_decoder_decoded_andMatrixInput_5_45 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_44 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_17 , core_id_ctrl_decoder_decoded_hi_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_45 , core_id_ctrl_decoder_decoded_andMatrixInput_3_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_45 , core_id_ctrl_decoder_decoded_andMatrixInput_1_45 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_45 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_29 , core_id_ctrl_decoder_decoded_hi_hi_lo_16 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_45 ={ core_id_ctrl_decoder_decoded_hi_hi_45 , core_id_ctrl_decoder_decoded_hi_lo_44 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_46 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_46 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_46 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_46 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_46 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_46 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_45 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_41 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_30 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_20 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_18 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_17 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_17 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_16 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_14 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_17 , core_id_ctrl_decoder_decoded_andMatrixInput_13_16 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_41 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_17 , core_id_ctrl_decoder_decoded_andMatrixInput_14_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_18 , core_id_ctrl_decoder_decoded_andMatrixInput_11_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_30 , core_id_ctrl_decoder_decoded_andMatrixInput_9_20 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_46 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_20 , core_id_ctrl_decoder_decoded_lo_hi_lo_16 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_46 ={ core_id_ctrl_decoder_decoded_lo_hi_46 , core_id_ctrl_decoder_decoded_lo_lo_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_45 , core_id_ctrl_decoder_decoded_andMatrixInput_7_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_46 , core_id_ctrl_decoder_decoded_andMatrixInput_5_46 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_45 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_18 , core_id_ctrl_decoder_decoded_hi_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_46 , core_id_ctrl_decoder_decoded_andMatrixInput_3_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_46 , core_id_ctrl_decoder_decoded_andMatrixInput_1_46 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_46 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_30 , core_id_ctrl_decoder_decoded_hi_hi_lo_17 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_46 ={ core_id_ctrl_decoder_decoded_hi_hi_46 , core_id_ctrl_decoder_decoded_hi_lo_45 }; 
    wire core__GEN_41 =&{ core_id_ctrl_decoder_decoded_hi_46 , core_id_ctrl_decoder_decoded_lo_46 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_47 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_47 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_47 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_47 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_47 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_47 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_46 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_42 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_31 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_21 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_19 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_18 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_18 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_17 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_15 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_5 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_15 , core_id_ctrl_decoder_decoded_andMatrixInput_15_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_18 , core_id_ctrl_decoder_decoded_andMatrixInput_13_17 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_42 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_18 , core_id_ctrl_decoder_decoded_lo_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_19 , core_id_ctrl_decoder_decoded_andMatrixInput_11_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_31 , core_id_ctrl_decoder_decoded_andMatrixInput_9_21 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_47 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_21 , core_id_ctrl_decoder_decoded_lo_hi_lo_17 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_47 ={ core_id_ctrl_decoder_decoded_lo_hi_47 , core_id_ctrl_decoder_decoded_lo_lo_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_46 , core_id_ctrl_decoder_decoded_andMatrixInput_7_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_47 , core_id_ctrl_decoder_decoded_andMatrixInput_5_47 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_46 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_19 , core_id_ctrl_decoder_decoded_hi_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_47 , core_id_ctrl_decoder_decoded_andMatrixInput_3_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_47 , core_id_ctrl_decoder_decoded_andMatrixInput_1_47 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_47 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_31 , core_id_ctrl_decoder_decoded_hi_hi_lo_18 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_47 ={ core_id_ctrl_decoder_decoded_hi_hi_47 , core_id_ctrl_decoder_decoded_hi_lo_46 }; 
    wire core__GEN_42 =&{ core_id_ctrl_decoder_decoded_hi_47 , core_id_ctrl_decoder_decoded_lo_47 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_48 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_48 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_48 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_48 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_48 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_48 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_47 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_43 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_32 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_22 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_20 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_19 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_19 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_18 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_16 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_16 , core_id_ctrl_decoder_decoded_andMatrixInput_15_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_19 , core_id_ctrl_decoder_decoded_andMatrixInput_13_18 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_43 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_19 , core_id_ctrl_decoder_decoded_lo_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_20 , core_id_ctrl_decoder_decoded_andMatrixInput_11_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_32 , core_id_ctrl_decoder_decoded_andMatrixInput_9_22 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_48 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_22 , core_id_ctrl_decoder_decoded_lo_hi_lo_18 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_48 ={ core_id_ctrl_decoder_decoded_lo_hi_48 , core_id_ctrl_decoder_decoded_lo_lo_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_47 , core_id_ctrl_decoder_decoded_andMatrixInput_7_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_48 , core_id_ctrl_decoder_decoded_andMatrixInput_5_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_47 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_20 , core_id_ctrl_decoder_decoded_hi_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_48 , core_id_ctrl_decoder_decoded_andMatrixInput_3_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_48 , core_id_ctrl_decoder_decoded_andMatrixInput_1_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_48 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_32 , core_id_ctrl_decoder_decoded_hi_hi_lo_19 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_48 ={ core_id_ctrl_decoder_decoded_hi_hi_48 , core_id_ctrl_decoder_decoded_hi_lo_47 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_49 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_49 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_49 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_49 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_49 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_49 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_48 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_44 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_33 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_23 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_21 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_20 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_20 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_19 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_17 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_20 , core_id_ctrl_decoder_decoded_andMatrixInput_13_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_44 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_20 , core_id_ctrl_decoder_decoded_andMatrixInput_14_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_21 , core_id_ctrl_decoder_decoded_andMatrixInput_11_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_33 , core_id_ctrl_decoder_decoded_andMatrixInput_9_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_49 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_23 , core_id_ctrl_decoder_decoded_lo_hi_lo_19 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_49 ={ core_id_ctrl_decoder_decoded_lo_hi_49 , core_id_ctrl_decoder_decoded_lo_lo_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_48 , core_id_ctrl_decoder_decoded_andMatrixInput_7_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_49 , core_id_ctrl_decoder_decoded_andMatrixInput_5_49 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_48 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_21 , core_id_ctrl_decoder_decoded_hi_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_49 , core_id_ctrl_decoder_decoded_andMatrixInput_3_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_49 , core_id_ctrl_decoder_decoded_andMatrixInput_1_49 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_49 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_33 , core_id_ctrl_decoder_decoded_hi_hi_lo_20 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_49 ={ core_id_ctrl_decoder_decoded_hi_hi_49 , core_id_ctrl_decoder_decoded_hi_lo_48 }; 
    wire core__GEN_43 =&{ core_id_ctrl_decoder_decoded_hi_49 , core_id_ctrl_decoder_decoded_lo_49 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_50 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_50 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_50 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_50 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_50 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_50 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_49 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_45 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_34 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_24 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_22 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_21 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_21 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_20 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_18 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_7 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_18 , core_id_ctrl_decoder_decoded_andMatrixInput_15_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_21 , core_id_ctrl_decoder_decoded_andMatrixInput_13_20 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_45 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_21 , core_id_ctrl_decoder_decoded_lo_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_22 , core_id_ctrl_decoder_decoded_andMatrixInput_11_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_34 , core_id_ctrl_decoder_decoded_andMatrixInput_9_24 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_50 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_24 , core_id_ctrl_decoder_decoded_lo_hi_lo_20 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_50 ={ core_id_ctrl_decoder_decoded_lo_hi_50 , core_id_ctrl_decoder_decoded_lo_lo_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_18 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_49 , core_id_ctrl_decoder_decoded_andMatrixInput_7_45 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_50 , core_id_ctrl_decoder_decoded_andMatrixInput_5_50 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_49 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_22 , core_id_ctrl_decoder_decoded_hi_lo_lo_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_50 , core_id_ctrl_decoder_decoded_andMatrixInput_3_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_50 , core_id_ctrl_decoder_decoded_andMatrixInput_1_50 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_50 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_34 , core_id_ctrl_decoder_decoded_hi_hi_lo_21 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_50 ={ core_id_ctrl_decoder_decoded_hi_hi_50 , core_id_ctrl_decoder_decoded_hi_lo_49 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_51 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_51 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_51 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_51 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_51 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_51 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_50 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_46 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_35 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_25 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_23 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_22 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_22 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_21 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_19 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_22 , core_id_ctrl_decoder_decoded_andMatrixInput_13_21 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_46 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_22 , core_id_ctrl_decoder_decoded_andMatrixInput_14_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_23 , core_id_ctrl_decoder_decoded_andMatrixInput_11_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_35 , core_id_ctrl_decoder_decoded_andMatrixInput_9_25 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_51 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_25 , core_id_ctrl_decoder_decoded_lo_hi_lo_21 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_51 ={ core_id_ctrl_decoder_decoded_lo_hi_51 , core_id_ctrl_decoder_decoded_lo_lo_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_19 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_50 , core_id_ctrl_decoder_decoded_andMatrixInput_7_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_51 , core_id_ctrl_decoder_decoded_andMatrixInput_5_51 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_50 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_23 , core_id_ctrl_decoder_decoded_hi_lo_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_51 , core_id_ctrl_decoder_decoded_andMatrixInput_3_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_51 , core_id_ctrl_decoder_decoded_andMatrixInput_1_51 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_35 , core_id_ctrl_decoder_decoded_hi_hi_lo_22 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_51 , core_id_ctrl_decoder_decoded_hi_lo_50 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_52 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_52 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_52 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_52 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_52 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_52 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_51 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_47 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_51 , core_id_ctrl_decoder_decoded_andMatrixInput_7_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_52 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_52 , core_id_ctrl_decoder_decoded_andMatrixInput_5_52 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_52 ={ core_id_ctrl_decoder_decoded_lo_hi_52 , core_id_ctrl_decoder_decoded_lo_lo_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_51 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_52 , core_id_ctrl_decoder_decoded_andMatrixInput_3_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_52 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_52 , core_id_ctrl_decoder_decoded_andMatrixInput_1_52 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_52 ={ core_id_ctrl_decoder_decoded_hi_hi_52 , core_id_ctrl_decoder_decoded_hi_lo_51 }; 
    wire core__GEN_44 =&{ core_id_ctrl_decoder_decoded_hi_52 , core_id_ctrl_decoder_decoded_lo_52 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_53 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_53 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_53 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_53 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_53 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_53 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_52 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_48 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_36 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_48 , core_id_ctrl_decoder_decoded_andMatrixInput_8_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_53 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_53 , core_id_ctrl_decoder_decoded_andMatrixInput_6_52 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_53 ={ core_id_ctrl_decoder_decoded_lo_hi_53 , core_id_ctrl_decoder_decoded_lo_lo_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_52 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_53 , core_id_ctrl_decoder_decoded_andMatrixInput_4_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_53 , core_id_ctrl_decoder_decoded_andMatrixInput_1_53 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_53 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_36 , core_id_ctrl_decoder_decoded_andMatrixInput_2_53 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_53 ={ core_id_ctrl_decoder_decoded_hi_hi_53 , core_id_ctrl_decoder_decoded_hi_lo_52 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_54 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_54 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_54 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_54 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_54 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_54 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_53 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_49 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_37 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_49 , core_id_ctrl_decoder_decoded_andMatrixInput_8_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_54 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_54 , core_id_ctrl_decoder_decoded_andMatrixInput_6_53 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_54 ={ core_id_ctrl_decoder_decoded_lo_hi_54 , core_id_ctrl_decoder_decoded_lo_lo_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_53 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_54 , core_id_ctrl_decoder_decoded_andMatrixInput_4_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_54 , core_id_ctrl_decoder_decoded_andMatrixInput_1_54 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_54 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_37 , core_id_ctrl_decoder_decoded_andMatrixInput_2_54 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_54 ={ core_id_ctrl_decoder_decoded_hi_hi_54 , core_id_ctrl_decoder_decoded_hi_lo_53 }; 
    wire core__GEN_45 =&{ core_id_ctrl_decoder_decoded_hi_54 , core_id_ctrl_decoder_decoded_lo_54 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_55 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_55 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_55 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_55 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_55 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_55 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_54 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_50 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_38 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_50 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_50 , core_id_ctrl_decoder_decoded_andMatrixInput_8_38 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_55 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_55 , core_id_ctrl_decoder_decoded_andMatrixInput_6_54 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_55 ={ core_id_ctrl_decoder_decoded_lo_hi_55 , core_id_ctrl_decoder_decoded_lo_lo_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_54 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_55 , core_id_ctrl_decoder_decoded_andMatrixInput_4_55 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_55 , core_id_ctrl_decoder_decoded_andMatrixInput_1_55 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_55 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_38 , core_id_ctrl_decoder_decoded_andMatrixInput_2_55 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_55 ={ core_id_ctrl_decoder_decoded_hi_hi_55 , core_id_ctrl_decoder_decoded_hi_lo_54 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_56 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_56 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_56 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_56 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_56 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_56 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_55 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_51 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_39 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_26 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_24 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_23 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_23 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_22 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_20 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_23 , core_id_ctrl_decoder_decoded_andMatrixInput_13_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_51 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_23 , core_id_ctrl_decoder_decoded_andMatrixInput_14_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_24 , core_id_ctrl_decoder_decoded_andMatrixInput_11_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_39 , core_id_ctrl_decoder_decoded_andMatrixInput_9_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_56 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_26 , core_id_ctrl_decoder_decoded_lo_hi_lo_22 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_56 ={ core_id_ctrl_decoder_decoded_lo_hi_56 , core_id_ctrl_decoder_decoded_lo_lo_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_20 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_55 , core_id_ctrl_decoder_decoded_andMatrixInput_7_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_56 , core_id_ctrl_decoder_decoded_andMatrixInput_5_56 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_55 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_24 , core_id_ctrl_decoder_decoded_hi_lo_lo_20 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_56 , core_id_ctrl_decoder_decoded_andMatrixInput_3_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_39 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_56 , core_id_ctrl_decoder_decoded_andMatrixInput_1_56 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_56 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_39 , core_id_ctrl_decoder_decoded_hi_hi_lo_23 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_56 ={ core_id_ctrl_decoder_decoded_hi_hi_56 , core_id_ctrl_decoder_decoded_hi_lo_55 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_57 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_57 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_57 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_57 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_57 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_57 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_56 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_52 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_52 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_56 , core_id_ctrl_decoder_decoded_andMatrixInput_7_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_57 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_57 , core_id_ctrl_decoder_decoded_andMatrixInput_5_57 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_57 ={ core_id_ctrl_decoder_decoded_lo_hi_57 , core_id_ctrl_decoder_decoded_lo_lo_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_56 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_57 , core_id_ctrl_decoder_decoded_andMatrixInput_3_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_57 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_57 , core_id_ctrl_decoder_decoded_andMatrixInput_1_57 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_57 ={ core_id_ctrl_decoder_decoded_hi_hi_57 , core_id_ctrl_decoder_decoded_hi_lo_56 }; 
    wire core__GEN_46 =&{ core_id_ctrl_decoder_decoded_hi_57 , core_id_ctrl_decoder_decoded_lo_57 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_58 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_58 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_58 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_58 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_58 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_58 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_57 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_53 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_40 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_53 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_53 , core_id_ctrl_decoder_decoded_andMatrixInput_8_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_58 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_58 , core_id_ctrl_decoder_decoded_andMatrixInput_6_57 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_58 ={ core_id_ctrl_decoder_decoded_lo_hi_58 , core_id_ctrl_decoder_decoded_lo_lo_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_57 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_58 , core_id_ctrl_decoder_decoded_andMatrixInput_4_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_58 , core_id_ctrl_decoder_decoded_andMatrixInput_1_58 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_58 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_40 , core_id_ctrl_decoder_decoded_andMatrixInput_2_58 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_58 ={ core_id_ctrl_decoder_decoded_hi_hi_58 , core_id_ctrl_decoder_decoded_hi_lo_57 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_59 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_59 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_59 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_59 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_59 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_59 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_58 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_54 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_41 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_54 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_54 , core_id_ctrl_decoder_decoded_andMatrixInput_8_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_59 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_59 , core_id_ctrl_decoder_decoded_andMatrixInput_6_58 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_59 ={ core_id_ctrl_decoder_decoded_lo_hi_59 , core_id_ctrl_decoder_decoded_lo_lo_54 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_58 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_59 , core_id_ctrl_decoder_decoded_andMatrixInput_4_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_59 , core_id_ctrl_decoder_decoded_andMatrixInput_1_59 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_59 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_41 , core_id_ctrl_decoder_decoded_andMatrixInput_2_59 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_59 ={ core_id_ctrl_decoder_decoded_hi_hi_59 , core_id_ctrl_decoder_decoded_hi_lo_58 }; 
    wire core__GEN_47 =&{ core_id_ctrl_decoder_decoded_hi_59 , core_id_ctrl_decoder_decoded_lo_59 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_60 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_60 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_60 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_60 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_60 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_60 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_59 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_55 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_42 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_27 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_55 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_42 , core_id_ctrl_decoder_decoded_andMatrixInput_9_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_60 , core_id_ctrl_decoder_decoded_andMatrixInput_6_59 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_60 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_27 , core_id_ctrl_decoder_decoded_andMatrixInput_7_55 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_60 ={ core_id_ctrl_decoder_decoded_lo_hi_60 , core_id_ctrl_decoder_decoded_lo_lo_55 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_59 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_60 , core_id_ctrl_decoder_decoded_andMatrixInput_4_60 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_60 , core_id_ctrl_decoder_decoded_andMatrixInput_1_60 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_60 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_42 , core_id_ctrl_decoder_decoded_andMatrixInput_2_60 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_60 ={ core_id_ctrl_decoder_decoded_hi_hi_60 , core_id_ctrl_decoder_decoded_hi_lo_59 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_61 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_61 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_61 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_61 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_61 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_61 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_60 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_56 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_43 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_28 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_25 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_24 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_24 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_23 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_24 , core_id_ctrl_decoder_decoded_andMatrixInput_12_24 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_56 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_24 , core_id_ctrl_decoder_decoded_andMatrixInput_13_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_28 , core_id_ctrl_decoder_decoded_andMatrixInput_10_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_56 , core_id_ctrl_decoder_decoded_andMatrixInput_8_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_61 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_28 , core_id_ctrl_decoder_decoded_lo_hi_lo_23 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_61 ={ core_id_ctrl_decoder_decoded_lo_hi_61 , core_id_ctrl_decoder_decoded_lo_lo_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_61 , core_id_ctrl_decoder_decoded_andMatrixInput_5_61 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_60 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_25 , core_id_ctrl_decoder_decoded_andMatrixInput_6_60 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_61 , core_id_ctrl_decoder_decoded_andMatrixInput_3_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_61 , core_id_ctrl_decoder_decoded_andMatrixInput_1_61 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_61 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_43 , core_id_ctrl_decoder_decoded_hi_hi_lo_24 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_61 ={ core_id_ctrl_decoder_decoded_hi_hi_61 , core_id_ctrl_decoder_decoded_hi_lo_60 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_62 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_62 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_62 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_62 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_62 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_62 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_61 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_57 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_44 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_29 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_26 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_25 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_25 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_24 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_21 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_25 , core_id_ctrl_decoder_decoded_andMatrixInput_13_24 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_57 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_25 , core_id_ctrl_decoder_decoded_andMatrixInput_14_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_26 , core_id_ctrl_decoder_decoded_andMatrixInput_11_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_44 , core_id_ctrl_decoder_decoded_andMatrixInput_9_29 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_62 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_29 , core_id_ctrl_decoder_decoded_lo_hi_lo_24 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_62 ={ core_id_ctrl_decoder_decoded_lo_hi_62 , core_id_ctrl_decoder_decoded_lo_lo_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_21 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_61 , core_id_ctrl_decoder_decoded_andMatrixInput_7_57 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_62 , core_id_ctrl_decoder_decoded_andMatrixInput_5_62 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_61 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_26 , core_id_ctrl_decoder_decoded_hi_lo_lo_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_62 , core_id_ctrl_decoder_decoded_andMatrixInput_3_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_62 , core_id_ctrl_decoder_decoded_andMatrixInput_1_62 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_62 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_44 , core_id_ctrl_decoder_decoded_hi_hi_lo_25 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_62 ={ core_id_ctrl_decoder_decoded_hi_hi_62 , core_id_ctrl_decoder_decoded_hi_lo_61 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_63 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_63 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_63 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_63 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_63 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_63 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_62 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_58 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_45 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_30 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_27 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_26 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_26 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_25 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_22 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_26 , core_id_ctrl_decoder_decoded_andMatrixInput_13_25 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_58 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_26 , core_id_ctrl_decoder_decoded_andMatrixInput_14_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_27 , core_id_ctrl_decoder_decoded_andMatrixInput_11_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_45 , core_id_ctrl_decoder_decoded_andMatrixInput_9_30 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_63 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_30 , core_id_ctrl_decoder_decoded_lo_hi_lo_25 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_63 ={ core_id_ctrl_decoder_decoded_lo_hi_63 , core_id_ctrl_decoder_decoded_lo_lo_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_22 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_62 , core_id_ctrl_decoder_decoded_andMatrixInput_7_58 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_63 , core_id_ctrl_decoder_decoded_andMatrixInput_5_63 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_62 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_27 , core_id_ctrl_decoder_decoded_hi_lo_lo_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_63 , core_id_ctrl_decoder_decoded_andMatrixInput_3_63 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_63 , core_id_ctrl_decoder_decoded_andMatrixInput_1_63 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_63 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_45 , core_id_ctrl_decoder_decoded_hi_hi_lo_26 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_63 ={ core_id_ctrl_decoder_decoded_hi_hi_63 , core_id_ctrl_decoder_decoded_hi_lo_62 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_64 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_64 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_64 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_64 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_64 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_64 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_63 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_59 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_46 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_31 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_28 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_27 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_27 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_26 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_23 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_27 , core_id_ctrl_decoder_decoded_andMatrixInput_13_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_59 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_27 , core_id_ctrl_decoder_decoded_andMatrixInput_14_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_28 , core_id_ctrl_decoder_decoded_andMatrixInput_11_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_46 , core_id_ctrl_decoder_decoded_andMatrixInput_9_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_64 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_31 , core_id_ctrl_decoder_decoded_lo_hi_lo_26 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_64 ={ core_id_ctrl_decoder_decoded_lo_hi_64 , core_id_ctrl_decoder_decoded_lo_lo_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_23 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_63 , core_id_ctrl_decoder_decoded_andMatrixInput_7_59 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_64 , core_id_ctrl_decoder_decoded_andMatrixInput_5_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_63 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_28 , core_id_ctrl_decoder_decoded_hi_lo_lo_23 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_64 , core_id_ctrl_decoder_decoded_andMatrixInput_3_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_46 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_64 , core_id_ctrl_decoder_decoded_andMatrixInput_1_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_64 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_46 , core_id_ctrl_decoder_decoded_hi_hi_lo_27 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_64 ={ core_id_ctrl_decoder_decoded_hi_hi_64 , core_id_ctrl_decoder_decoded_hi_lo_63 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_65 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_65 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_65 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_65 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_65 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_65 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_64 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_60 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_47 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_32 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_29 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_28 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_28 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_27 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_28 , core_id_ctrl_decoder_decoded_andMatrixInput_12_28 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_60 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_28 , core_id_ctrl_decoder_decoded_andMatrixInput_13_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_32 , core_id_ctrl_decoder_decoded_andMatrixInput_10_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_60 , core_id_ctrl_decoder_decoded_andMatrixInput_8_47 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_65 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_32 , core_id_ctrl_decoder_decoded_lo_hi_lo_27 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_65 ={ core_id_ctrl_decoder_decoded_lo_hi_65 , core_id_ctrl_decoder_decoded_lo_lo_60 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_65 , core_id_ctrl_decoder_decoded_andMatrixInput_5_65 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_64 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_29 , core_id_ctrl_decoder_decoded_andMatrixInput_6_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_65 , core_id_ctrl_decoder_decoded_andMatrixInput_3_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_65 , core_id_ctrl_decoder_decoded_andMatrixInput_1_65 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_65 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_47 , core_id_ctrl_decoder_decoded_hi_hi_lo_28 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_65 ={ core_id_ctrl_decoder_decoded_hi_hi_65 , core_id_ctrl_decoder_decoded_hi_lo_64 }; 
    wire core__GEN_48 =&{ core_id_ctrl_decoder_decoded_hi_65 , core_id_ctrl_decoder_decoded_lo_65 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_66 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_66 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_66 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_66 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_66 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_66 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_65 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_61 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_48 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_33 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_30 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_29 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_29 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_28 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_24 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_29 , core_id_ctrl_decoder_decoded_andMatrixInput_13_28 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_61 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_29 , core_id_ctrl_decoder_decoded_andMatrixInput_14_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_28 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_30 , core_id_ctrl_decoder_decoded_andMatrixInput_11_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_48 , core_id_ctrl_decoder_decoded_andMatrixInput_9_33 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_66 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_33 , core_id_ctrl_decoder_decoded_lo_hi_lo_28 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_66 ={ core_id_ctrl_decoder_decoded_lo_hi_66 , core_id_ctrl_decoder_decoded_lo_lo_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_24 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_65 , core_id_ctrl_decoder_decoded_andMatrixInput_7_61 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_66 , core_id_ctrl_decoder_decoded_andMatrixInput_5_66 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_65 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_30 , core_id_ctrl_decoder_decoded_hi_lo_lo_24 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_66 , core_id_ctrl_decoder_decoded_andMatrixInput_3_66 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_66 , core_id_ctrl_decoder_decoded_andMatrixInput_1_66 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_66 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_48 , core_id_ctrl_decoder_decoded_hi_hi_lo_29 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_66 ={ core_id_ctrl_decoder_decoded_hi_hi_66 , core_id_ctrl_decoder_decoded_hi_lo_65 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_67 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_67 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_67 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_67 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_67 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_67 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_66 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_62 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_49 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_34 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_31 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_30 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_30 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_29 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_25 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_30 , core_id_ctrl_decoder_decoded_andMatrixInput_13_29 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_62 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_30 , core_id_ctrl_decoder_decoded_andMatrixInput_14_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_29 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_31 , core_id_ctrl_decoder_decoded_andMatrixInput_11_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_49 , core_id_ctrl_decoder_decoded_andMatrixInput_9_34 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_67 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_34 , core_id_ctrl_decoder_decoded_lo_hi_lo_29 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_67 ={ core_id_ctrl_decoder_decoded_lo_hi_67 , core_id_ctrl_decoder_decoded_lo_lo_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_25 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_66 , core_id_ctrl_decoder_decoded_andMatrixInput_7_62 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_67 , core_id_ctrl_decoder_decoded_andMatrixInput_5_67 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_66 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_31 , core_id_ctrl_decoder_decoded_hi_lo_lo_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_67 , core_id_ctrl_decoder_decoded_andMatrixInput_3_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_49 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_67 , core_id_ctrl_decoder_decoded_andMatrixInput_1_67 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_67 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_49 , core_id_ctrl_decoder_decoded_hi_hi_lo_30 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_67 ={ core_id_ctrl_decoder_decoded_hi_hi_67 , core_id_ctrl_decoder_decoded_hi_lo_66 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_68 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_68 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_68 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_68 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_68 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_68 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_67 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_63 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_50 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_35 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_32 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_31 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_31 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_32 , core_id_ctrl_decoder_decoded_andMatrixInput_11_31 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_63 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_31 , core_id_ctrl_decoder_decoded_andMatrixInput_12_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_63 , core_id_ctrl_decoder_decoded_andMatrixInput_8_50 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_68 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_35 , core_id_ctrl_decoder_decoded_andMatrixInput_9_35 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_68 ={ core_id_ctrl_decoder_decoded_lo_hi_68 , core_id_ctrl_decoder_decoded_lo_lo_63 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_68 , core_id_ctrl_decoder_decoded_andMatrixInput_5_68 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_67 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_32 , core_id_ctrl_decoder_decoded_andMatrixInput_6_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_68 , core_id_ctrl_decoder_decoded_andMatrixInput_3_68 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_50 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_68 , core_id_ctrl_decoder_decoded_andMatrixInput_1_68 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_68 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_50 , core_id_ctrl_decoder_decoded_hi_hi_lo_31 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_68 ={ core_id_ctrl_decoder_decoded_hi_hi_68 , core_id_ctrl_decoder_decoded_hi_lo_67 }; 
    wire core__GEN_49 =&{ core_id_ctrl_decoder_decoded_hi_68 , core_id_ctrl_decoder_decoded_lo_68 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_69 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_69 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_69 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_69 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_69 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_69 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_68 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_64 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_51 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_36 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_33 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_32 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_32 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_30 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_26 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_8 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_15_8 , core_id_ctrl_decoder_decoded_andMatrixInput_16_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_13_30 , core_id_ctrl_decoder_decoded_andMatrixInput_14_26 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_64 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_32 , core_id_ctrl_decoder_decoded_lo_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_30 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_32 , core_id_ctrl_decoder_decoded_andMatrixInput_12_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_36 , core_id_ctrl_decoder_decoded_andMatrixInput_10_33 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_69 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_36 , core_id_ctrl_decoder_decoded_lo_hi_lo_30 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_69 ={ core_id_ctrl_decoder_decoded_lo_hi_69 , core_id_ctrl_decoder_decoded_lo_lo_64 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_26 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_64 , core_id_ctrl_decoder_decoded_andMatrixInput_8_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_69 , core_id_ctrl_decoder_decoded_andMatrixInput_6_68 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_68 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_33 , core_id_ctrl_decoder_decoded_hi_lo_lo_26 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_69 , core_id_ctrl_decoder_decoded_andMatrixInput_4_69 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_69 , core_id_ctrl_decoder_decoded_andMatrixInput_1_69 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_hi_51 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_2_69 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_hi_69 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_51 , core_id_ctrl_decoder_decoded_hi_hi_lo_32 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_hi_69 ={ core_id_ctrl_decoder_decoded_hi_hi_69 , core_id_ctrl_decoder_decoded_hi_lo_68 }; 
    wire core__GEN_50 =&{ core_id_ctrl_decoder_decoded_hi_69 , core_id_ctrl_decoder_decoded_lo_69 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_70 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_70 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_70 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_70 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_70 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_70 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_69 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_65 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_52 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_37 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_34 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_33 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_33 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_31 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_27 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_9 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_3 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_17_2 , core_id_ctrl_decoder_decoded_andMatrixInput_18_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_15_9 , core_id_ctrl_decoder_decoded_andMatrixInput_16_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_65 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_33 , core_id_ctrl_decoder_decoded_lo_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_31 ={ core_id_ctrl_decoder_decoded_andMatrixInput_13_31 , core_id_ctrl_decoder_decoded_andMatrixInput_14_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_34 , core_id_ctrl_decoder_decoded_andMatrixInput_11_33 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_hi_37 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_12_33 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_lo_hi_70 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_37 , core_id_ctrl_decoder_decoded_lo_hi_lo_31 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_lo_70 ={ core_id_ctrl_decoder_decoded_lo_hi_70 , core_id_ctrl_decoder_decoded_lo_lo_65 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_27 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_52 , core_id_ctrl_decoder_decoded_andMatrixInput_9_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_5_70 , core_id_ctrl_decoder_decoded_andMatrixInput_6_69 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_hi_34 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_7_65 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_lo_69 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_34 , core_id_ctrl_decoder_decoded_hi_lo_lo_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_70 , core_id_ctrl_decoder_decoded_andMatrixInput_4_70 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_70 , core_id_ctrl_decoder_decoded_andMatrixInput_1_70 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_hi_52 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_2_70 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_hi_hi_70 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_52 , core_id_ctrl_decoder_decoded_hi_hi_lo_33 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_hi_70 ={ core_id_ctrl_decoder_decoded_hi_hi_70 , core_id_ctrl_decoder_decoded_hi_lo_69 }; 
    wire core__GEN_51 =&{ core_id_ctrl_decoder_decoded_hi_70 , core_id_ctrl_decoder_decoded_lo_70 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_71 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_71 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_71 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_71 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_71 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_71 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_70 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_66 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_53 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_38 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_35 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_34 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_34 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_32 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_28 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_10 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_4 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_3 = core_id_ctrl_decoder_decoded_plaInput [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_3 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_2 = core_id_ctrl_decoder_decoded_plaInput [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_2 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_2 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_2 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_2 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_2 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_2 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_2 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_2 , core_id_ctrl_decoder_decoded_andMatrixInput_26_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_10 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_27_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_2 , core_id_ctrl_decoder_decoded_andMatrixInput_24_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_2 , core_id_ctrl_decoder_decoded_andMatrixInput_22_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_34 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_2 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_66 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_34 , core_id_ctrl_decoder_decoded_lo_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_3 , core_id_ctrl_decoder_decoded_andMatrixInput_19_2 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_32 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_20_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_4 , core_id_ctrl_decoder_decoded_andMatrixInput_17_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_28 , core_id_ctrl_decoder_decoded_andMatrixInput_15_10 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_38 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_71 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_38 , core_id_ctrl_decoder_decoded_lo_hi_lo_32 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_71 ={ core_id_ctrl_decoder_decoded_lo_hi_71 , core_id_ctrl_decoder_decoded_lo_lo_66 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_34 , core_id_ctrl_decoder_decoded_andMatrixInput_12_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_28 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_13_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_38 , core_id_ctrl_decoder_decoded_andMatrixInput_10_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_66 , core_id_ctrl_decoder_decoded_andMatrixInput_8_53 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_35 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_70 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_35 , core_id_ctrl_decoder_decoded_hi_lo_lo_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_71 , core_id_ctrl_decoder_decoded_andMatrixInput_5_71 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_34 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_andMatrixInput_6_70 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_71 , core_id_ctrl_decoder_decoded_andMatrixInput_3_71 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_71 , core_id_ctrl_decoder_decoded_andMatrixInput_1_71 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_53 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_2 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_71 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_53 , core_id_ctrl_decoder_decoded_hi_hi_lo_34 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_71 ={ core_id_ctrl_decoder_decoded_hi_hi_71 , core_id_ctrl_decoder_decoded_hi_lo_70 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_72 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_72 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_72 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_72 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_72 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_72 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_71 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_67 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_54 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_39 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_36 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_35 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_35 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_33 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_29 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_11 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_5 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_4 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_4 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_3 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_3 = core_id_ctrl_decoder_decoded_plaInput [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_3 = core_id_ctrl_decoder_decoded_invInputs [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_3 = core_id_ctrl_decoder_decoded_plaInput [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_3 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_3 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_3 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_3 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_3 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_1 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_1 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_1 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_1 , core_id_ctrl_decoder_decoded_andMatrixInput_29_1 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_11 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_andMatrixInput_30_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_3 , core_id_ctrl_decoder_decoded_andMatrixInput_27_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_3 , core_id_ctrl_decoder_decoded_andMatrixInput_25_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_35 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_67 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_35 , core_id_ctrl_decoder_decoded_lo_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_3 , core_id_ctrl_decoder_decoded_andMatrixInput_23_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_3 , core_id_ctrl_decoder_decoded_andMatrixInput_21_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_33 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_4 , core_id_ctrl_decoder_decoded_andMatrixInput_19_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_5 , core_id_ctrl_decoder_decoded_andMatrixInput_17_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_39 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_72 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_39 , core_id_ctrl_decoder_decoded_lo_hi_lo_33 }; 
    wire[14:0] core_id_ctrl_decoder_decoded_lo_72 ={ core_id_ctrl_decoder_decoded_lo_hi_72 , core_id_ctrl_decoder_decoded_lo_lo_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_29 , core_id_ctrl_decoder_decoded_andMatrixInput_15_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_35 , core_id_ctrl_decoder_decoded_andMatrixInput_13_33 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_29 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_36 , core_id_ctrl_decoder_decoded_andMatrixInput_11_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_54 , core_id_ctrl_decoder_decoded_andMatrixInput_9_39 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_36 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_71 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_36 , core_id_ctrl_decoder_decoded_hi_lo_lo_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_71 , core_id_ctrl_decoder_decoded_andMatrixInput_7_67 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_72 , core_id_ctrl_decoder_decoded_andMatrixInput_5_72 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_35 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_72 , core_id_ctrl_decoder_decoded_andMatrixInput_3_72 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_72 , core_id_ctrl_decoder_decoded_andMatrixInput_1_72 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_54 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_3 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_72 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_54 , core_id_ctrl_decoder_decoded_hi_hi_lo_35 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_72 ={ core_id_ctrl_decoder_decoded_hi_hi_72 , core_id_ctrl_decoder_decoded_hi_lo_71 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_73 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_73 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_73 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_73 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_73 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_73 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_72 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_68 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_55 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_40 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_37 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_36 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_36 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_34 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_36 , core_id_ctrl_decoder_decoded_andMatrixInput_12_36 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_68 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_36 , core_id_ctrl_decoder_decoded_andMatrixInput_13_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_40 , core_id_ctrl_decoder_decoded_andMatrixInput_10_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_68 , core_id_ctrl_decoder_decoded_andMatrixInput_8_55 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_73 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_40 , core_id_ctrl_decoder_decoded_lo_hi_lo_34 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_73 ={ core_id_ctrl_decoder_decoded_lo_hi_73 , core_id_ctrl_decoder_decoded_lo_lo_68 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_73 , core_id_ctrl_decoder_decoded_andMatrixInput_5_73 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_72 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_37 , core_id_ctrl_decoder_decoded_andMatrixInput_6_72 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_36 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_73 , core_id_ctrl_decoder_decoded_andMatrixInput_3_73 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_55 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_73 , core_id_ctrl_decoder_decoded_andMatrixInput_1_73 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_73 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_55 , core_id_ctrl_decoder_decoded_hi_hi_lo_36 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_73 ={ core_id_ctrl_decoder_decoded_hi_hi_73 , core_id_ctrl_decoder_decoded_hi_lo_72 }; 
    wire core__GEN_52 =&{ core_id_ctrl_decoder_decoded_hi_73 , core_id_ctrl_decoder_decoded_lo_73 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_74 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_74 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_74 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_74 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_74 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_74 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_73 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_69 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_56 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_41 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_38 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_37 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_41 , core_id_ctrl_decoder_decoded_andMatrixInput_10_38 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_69 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_37 , core_id_ctrl_decoder_decoded_andMatrixInput_11_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_73 , core_id_ctrl_decoder_decoded_andMatrixInput_7_69 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_74 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_41 , core_id_ctrl_decoder_decoded_andMatrixInput_8_56 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_74 ={ core_id_ctrl_decoder_decoded_lo_hi_74 , core_id_ctrl_decoder_decoded_lo_lo_69 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_74 , core_id_ctrl_decoder_decoded_andMatrixInput_4_74 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_73 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_38 , core_id_ctrl_decoder_decoded_andMatrixInput_5_74 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_56 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_74 , core_id_ctrl_decoder_decoded_andMatrixInput_1_74 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_74 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_56 , core_id_ctrl_decoder_decoded_andMatrixInput_2_74 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_hi_74 ={ core_id_ctrl_decoder_decoded_hi_hi_74 , core_id_ctrl_decoder_decoded_hi_lo_73 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_75 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_75 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_75 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_75 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_75 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_75 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_74 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_70 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_57 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_42 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_39 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_38 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_37 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_35 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_30 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_12 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_6 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_5 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_5 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_4 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_4 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_4 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_4 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_4 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_4 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_4 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_4 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_4 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_4 , core_id_ctrl_decoder_decoded_andMatrixInput_26_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_12 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_27_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_4 , core_id_ctrl_decoder_decoded_andMatrixInput_24_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_4 , core_id_ctrl_decoder_decoded_andMatrixInput_22_4 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_38 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_70 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_38 , core_id_ctrl_decoder_decoded_lo_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_5 , core_id_ctrl_decoder_decoded_andMatrixInput_19_4 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_35 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_20_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_6 , core_id_ctrl_decoder_decoded_andMatrixInput_17_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_30 , core_id_ctrl_decoder_decoded_andMatrixInput_15_12 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_42 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_75 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_42 , core_id_ctrl_decoder_decoded_lo_hi_lo_35 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_75 ={ core_id_ctrl_decoder_decoded_lo_hi_75 , core_id_ctrl_decoder_decoded_lo_lo_70 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_38 , core_id_ctrl_decoder_decoded_andMatrixInput_12_37 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_30 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_13_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_42 , core_id_ctrl_decoder_decoded_andMatrixInput_10_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_70 , core_id_ctrl_decoder_decoded_andMatrixInput_8_57 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_39 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_74 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_39 , core_id_ctrl_decoder_decoded_hi_lo_lo_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_75 , core_id_ctrl_decoder_decoded_andMatrixInput_5_75 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_37 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_andMatrixInput_6_74 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_4 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_75 , core_id_ctrl_decoder_decoded_andMatrixInput_3_75 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_75 , core_id_ctrl_decoder_decoded_andMatrixInput_1_75 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_57 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_4 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_75 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_57 , core_id_ctrl_decoder_decoded_hi_hi_lo_37 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_75 ={ core_id_ctrl_decoder_decoded_hi_hi_75 , core_id_ctrl_decoder_decoded_hi_lo_74 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_76 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_76 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_76 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_76 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_76 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_76 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_75 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_71 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_58 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_43 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_40 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_39 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_38 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_36 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_31 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_13 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_7 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_6 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_6 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_5 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_5 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_5 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_5 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_5 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_5 = core_id_ctrl_decoder_decoded_invInputs [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_5 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_5 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_5 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_2 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_2 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_2 = core_id_ctrl_decoder_decoded_invInputs [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_31 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_lo ={ core_id_ctrl_decoder_decoded_andMatrixInput_30_2 , core_id_ctrl_decoder_decoded_andMatrixInput_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_2 , core_id_ctrl_decoder_decoded_andMatrixInput_29_2 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_lo_13 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_5 , core_id_ctrl_decoder_decoded_andMatrixInput_27_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_5 , core_id_ctrl_decoder_decoded_andMatrixInput_25_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_39 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_lo_71 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_39 , core_id_ctrl_decoder_decoded_lo_lo_lo_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_5 , core_id_ctrl_decoder_decoded_andMatrixInput_23_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_5 , core_id_ctrl_decoder_decoded_andMatrixInput_21_5 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_36 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_6 , core_id_ctrl_decoder_decoded_andMatrixInput_19_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_7 , core_id_ctrl_decoder_decoded_andMatrixInput_17_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_43 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_76 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_43 , core_id_ctrl_decoder_decoded_lo_hi_lo_36 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_lo_76 ={ core_id_ctrl_decoder_decoded_lo_hi_76 , core_id_ctrl_decoder_decoded_lo_lo_71 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_31 , core_id_ctrl_decoder_decoded_andMatrixInput_15_13 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_38 , core_id_ctrl_decoder_decoded_andMatrixInput_13_36 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_31 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_40 , core_id_ctrl_decoder_decoded_andMatrixInput_11_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_58 , core_id_ctrl_decoder_decoded_andMatrixInput_9_43 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_40 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_75 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_40 , core_id_ctrl_decoder_decoded_hi_lo_lo_31 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_2 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_75 , core_id_ctrl_decoder_decoded_andMatrixInput_7_71 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_76 , core_id_ctrl_decoder_decoded_andMatrixInput_5_76 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_38 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_76 , core_id_ctrl_decoder_decoded_andMatrixInput_3_76 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_76 , core_id_ctrl_decoder_decoded_andMatrixInput_1_76 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_58 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_5 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_76 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_58 , core_id_ctrl_decoder_decoded_hi_hi_lo_38 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_76 ={ core_id_ctrl_decoder_decoded_hi_hi_76 , core_id_ctrl_decoder_decoded_hi_lo_75 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_77 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_77 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_77 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_77 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_77 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_77 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_76 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_72 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_59 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_44 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_41 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_40 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_39 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_37 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_32 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_14 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_14 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_32 , core_id_ctrl_decoder_decoded_andMatrixInput_15_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_39 , core_id_ctrl_decoder_decoded_andMatrixInput_13_37 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_72 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_40 , core_id_ctrl_decoder_decoded_lo_lo_lo_14 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_37 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_41 , core_id_ctrl_decoder_decoded_andMatrixInput_11_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_59 , core_id_ctrl_decoder_decoded_andMatrixInput_9_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_77 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_44 , core_id_ctrl_decoder_decoded_lo_hi_lo_37 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_77 ={ core_id_ctrl_decoder_decoded_lo_hi_77 , core_id_ctrl_decoder_decoded_lo_lo_72 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_32 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_76 , core_id_ctrl_decoder_decoded_andMatrixInput_7_72 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_77 , core_id_ctrl_decoder_decoded_andMatrixInput_5_77 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_76 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_41 , core_id_ctrl_decoder_decoded_hi_lo_lo_32 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_39 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_77 , core_id_ctrl_decoder_decoded_andMatrixInput_3_77 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_59 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_77 , core_id_ctrl_decoder_decoded_andMatrixInput_1_77 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_77 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_59 , core_id_ctrl_decoder_decoded_hi_hi_lo_39 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_77 ={ core_id_ctrl_decoder_decoded_hi_hi_77 , core_id_ctrl_decoder_decoded_hi_lo_76 }; 
    wire core__GEN_53 =&{ core_id_ctrl_decoder_decoded_hi_77 , core_id_ctrl_decoder_decoded_lo_77 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_78 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_78 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_78 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_78 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_78 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_78 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_77 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_73 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_60 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_45 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_42 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_41 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_45 , core_id_ctrl_decoder_decoded_andMatrixInput_10_42 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_73 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_41 , core_id_ctrl_decoder_decoded_andMatrixInput_11_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_77 , core_id_ctrl_decoder_decoded_andMatrixInput_7_73 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_78 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_45 , core_id_ctrl_decoder_decoded_andMatrixInput_8_60 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_78 ={ core_id_ctrl_decoder_decoded_lo_hi_78 , core_id_ctrl_decoder_decoded_lo_lo_73 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_78 , core_id_ctrl_decoder_decoded_andMatrixInput_4_78 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_77 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_42 , core_id_ctrl_decoder_decoded_andMatrixInput_5_78 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_60 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_78 , core_id_ctrl_decoder_decoded_andMatrixInput_1_78 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_78 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_60 , core_id_ctrl_decoder_decoded_andMatrixInput_2_78 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_hi_78 ={ core_id_ctrl_decoder_decoded_hi_hi_78 , core_id_ctrl_decoder_decoded_hi_lo_77 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_79 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_79 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_79 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_79 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_79 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_79 = core_id_ctrl_decoder_decoded_invInputs [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_78 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_74 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_61 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_46 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_43 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_42 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_40 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_38 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_33 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_15 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_15 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_33 , core_id_ctrl_decoder_decoded_andMatrixInput_15_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_40 , core_id_ctrl_decoder_decoded_andMatrixInput_13_38 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_74 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_42 , core_id_ctrl_decoder_decoded_lo_lo_lo_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_38 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_43 , core_id_ctrl_decoder_decoded_andMatrixInput_11_42 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_46 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_61 , core_id_ctrl_decoder_decoded_andMatrixInput_9_46 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_79 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_46 , core_id_ctrl_decoder_decoded_lo_hi_lo_38 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_79 ={ core_id_ctrl_decoder_decoded_lo_hi_79 , core_id_ctrl_decoder_decoded_lo_lo_74 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_33 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_78 , core_id_ctrl_decoder_decoded_andMatrixInput_7_74 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_79 , core_id_ctrl_decoder_decoded_andMatrixInput_5_79 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_78 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_43 , core_id_ctrl_decoder_decoded_hi_lo_lo_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_79 , core_id_ctrl_decoder_decoded_andMatrixInput_3_79 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_61 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_79 , core_id_ctrl_decoder_decoded_andMatrixInput_1_79 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_79 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_61 , core_id_ctrl_decoder_decoded_hi_hi_lo_40 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_79 ={ core_id_ctrl_decoder_decoded_hi_hi_79 , core_id_ctrl_decoder_decoded_hi_lo_78 }; 
    wire core__GEN_54 =&{ core_id_ctrl_decoder_decoded_hi_79 , core_id_ctrl_decoder_decoded_lo_79 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_80 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_80 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_80 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_80 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_80 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_80 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_79 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_75 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_62 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_47 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_44 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_43 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_41 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_39 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_34 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_16 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_16 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_34 , core_id_ctrl_decoder_decoded_andMatrixInput_15_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_43 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_41 , core_id_ctrl_decoder_decoded_andMatrixInput_13_39 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_75 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_43 , core_id_ctrl_decoder_decoded_lo_lo_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_39 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_44 , core_id_ctrl_decoder_decoded_andMatrixInput_11_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_62 , core_id_ctrl_decoder_decoded_andMatrixInput_9_47 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_80 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_47 , core_id_ctrl_decoder_decoded_lo_hi_lo_39 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_80 ={ core_id_ctrl_decoder_decoded_lo_hi_80 , core_id_ctrl_decoder_decoded_lo_lo_75 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_34 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_79 , core_id_ctrl_decoder_decoded_andMatrixInput_7_75 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_80 , core_id_ctrl_decoder_decoded_andMatrixInput_5_80 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_79 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_44 , core_id_ctrl_decoder_decoded_hi_lo_lo_34 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_41 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_80 , core_id_ctrl_decoder_decoded_andMatrixInput_3_80 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_62 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_80 , core_id_ctrl_decoder_decoded_andMatrixInput_1_80 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_80 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_62 , core_id_ctrl_decoder_decoded_hi_hi_lo_41 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_80 ={ core_id_ctrl_decoder_decoded_hi_hi_80 , core_id_ctrl_decoder_decoded_hi_lo_79 }; 
    wire core__GEN_55 =&{ core_id_ctrl_decoder_decoded_hi_80 , core_id_ctrl_decoder_decoded_lo_80 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_81 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_81 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_81 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_81 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_81 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_81 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_80 = core_id_ctrl_decoder_decoded_plaInput [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_76 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_63 = core_id_ctrl_decoder_decoded_plaInput [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_48 = core_id_ctrl_decoder_decoded_invInputs [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_45 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_44 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_42 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_40 = core_id_ctrl_decoder_decoded_invInputs [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_35 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_17 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_17 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_35 , core_id_ctrl_decoder_decoded_andMatrixInput_15_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_44 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_42 , core_id_ctrl_decoder_decoded_andMatrixInput_13_40 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_76 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_44 , core_id_ctrl_decoder_decoded_lo_lo_lo_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_40 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_45 , core_id_ctrl_decoder_decoded_andMatrixInput_11_44 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_63 , core_id_ctrl_decoder_decoded_andMatrixInput_9_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_81 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_48 , core_id_ctrl_decoder_decoded_lo_hi_lo_40 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_81 ={ core_id_ctrl_decoder_decoded_lo_hi_81 , core_id_ctrl_decoder_decoded_lo_lo_76 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_35 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_80 , core_id_ctrl_decoder_decoded_andMatrixInput_7_76 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_45 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_81 , core_id_ctrl_decoder_decoded_andMatrixInput_5_81 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_80 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_45 , core_id_ctrl_decoder_decoded_hi_lo_lo_35 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_42 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_81 , core_id_ctrl_decoder_decoded_andMatrixInput_3_81 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_63 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_81 , core_id_ctrl_decoder_decoded_andMatrixInput_1_81 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_81 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_63 , core_id_ctrl_decoder_decoded_hi_hi_lo_42 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_81 ={ core_id_ctrl_decoder_decoded_hi_hi_81 , core_id_ctrl_decoder_decoded_hi_lo_80 }; 
    wire core__GEN_56 =&{ core_id_ctrl_decoder_decoded_hi_81 , core_id_ctrl_decoder_decoded_lo_81 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_82 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_82 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_82 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_82 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_82 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_82 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_81 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_77 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_64 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_49 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_46 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_45 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_43 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_41 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_36 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_18 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_8 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_7 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_7 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_6 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_6 = core_id_ctrl_decoder_decoded_plaInput [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_6 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_6 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_6 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_6 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_6 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_6 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_6 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_25_6 , core_id_ctrl_decoder_decoded_andMatrixInput_26_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_lo_18 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_27_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_23_6 , core_id_ctrl_decoder_decoded_andMatrixInput_24_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_21_6 , core_id_ctrl_decoder_decoded_andMatrixInput_22_6 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_45 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_lo_77 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_45 , core_id_ctrl_decoder_decoded_lo_lo_lo_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_7 , core_id_ctrl_decoder_decoded_andMatrixInput_19_6 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_lo_41 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_20_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_8 , core_id_ctrl_decoder_decoded_andMatrixInput_17_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_36 , core_id_ctrl_decoder_decoded_andMatrixInput_15_18 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_49 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_lo_hi_82 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_49 , core_id_ctrl_decoder_decoded_lo_hi_lo_41 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_lo_82 ={ core_id_ctrl_decoder_decoded_lo_hi_82 , core_id_ctrl_decoder_decoded_lo_lo_77 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_11_45 , core_id_ctrl_decoder_decoded_andMatrixInput_12_43 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_lo_36 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_13_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_49 , core_id_ctrl_decoder_decoded_andMatrixInput_10_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_7_77 , core_id_ctrl_decoder_decoded_andMatrixInput_8_64 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_46 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_lo_81 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_46 , core_id_ctrl_decoder_decoded_hi_lo_lo_36 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_82 , core_id_ctrl_decoder_decoded_andMatrixInput_5_82 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_lo_43 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_6 , core_id_ctrl_decoder_decoded_andMatrixInput_6_81 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_82 , core_id_ctrl_decoder_decoded_andMatrixInput_3_82 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_82 , core_id_ctrl_decoder_decoded_andMatrixInput_1_82 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_64 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_6 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_hi_hi_82 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_64 , core_id_ctrl_decoder_decoded_hi_hi_lo_43 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_hi_82 ={ core_id_ctrl_decoder_decoded_hi_hi_82 , core_id_ctrl_decoder_decoded_hi_lo_81 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_83 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_83 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_83 = core_id_ctrl_decoder_decoded_invInputs [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_83 = core_id_ctrl_decoder_decoded_invInputs [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_83 = core_id_ctrl_decoder_decoded_plaInput [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_83 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_82 = core_id_ctrl_decoder_decoded_plaInput [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_78 = core_id_ctrl_decoder_decoded_invInputs [7]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_65 = core_id_ctrl_decoder_decoded_invInputs [8]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_50 = core_id_ctrl_decoder_decoded_invInputs [9]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_47 = core_id_ctrl_decoder_decoded_invInputs [10]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_46 = core_id_ctrl_decoder_decoded_invInputs [11]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_12_44 = core_id_ctrl_decoder_decoded_invInputs [12]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_13_42 = core_id_ctrl_decoder_decoded_invInputs [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_14_37 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_15_19 = core_id_ctrl_decoder_decoded_invInputs [15]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_16_9 = core_id_ctrl_decoder_decoded_invInputs [16]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_17_8 = core_id_ctrl_decoder_decoded_invInputs [17]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_18_8 = core_id_ctrl_decoder_decoded_invInputs [18]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_19_7 = core_id_ctrl_decoder_decoded_invInputs [19]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_20_7 = core_id_ctrl_decoder_decoded_invInputs [20]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_21_7 = core_id_ctrl_decoder_decoded_plaInput [21]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_22_7 = core_id_ctrl_decoder_decoded_invInputs [22]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_23_7 = core_id_ctrl_decoder_decoded_invInputs [23]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_24_7 = core_id_ctrl_decoder_decoded_plaInput [24]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_25_7 = core_id_ctrl_decoder_decoded_plaInput [25]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_26_7 = core_id_ctrl_decoder_decoded_invInputs [26]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_27_7 = core_id_ctrl_decoder_decoded_plaInput [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_28_3 = core_id_ctrl_decoder_decoded_plaInput [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_29_3 = core_id_ctrl_decoder_decoded_plaInput [29]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_30_3 = core_id_ctrl_decoder_decoded_plaInput [30]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_31_1 = core_id_ctrl_decoder_decoded_invInputs [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_lo_1 ={ core_id_ctrl_decoder_decoded_andMatrixInput_30_3 , core_id_ctrl_decoder_decoded_andMatrixInput_31_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_28_3 , core_id_ctrl_decoder_decoded_andMatrixInput_29_3 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_lo_19 ={ core_id_ctrl_decoder_decoded_lo_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_lo_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_26_7 , core_id_ctrl_decoder_decoded_andMatrixInput_27_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_24_7 , core_id_ctrl_decoder_decoded_andMatrixInput_25_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_lo_hi_46 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_lo_lo_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_lo_78 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_46 , core_id_ctrl_decoder_decoded_lo_lo_lo_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_22_7 , core_id_ctrl_decoder_decoded_andMatrixInput_23_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_20_7 , core_id_ctrl_decoder_decoded_andMatrixInput_21_7 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_lo_42 ={ core_id_ctrl_decoder_decoded_lo_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_lo_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_18_8 , core_id_ctrl_decoder_decoded_andMatrixInput_19_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_16_9 , core_id_ctrl_decoder_decoded_andMatrixInput_17_8 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_lo_hi_hi_50 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_lo_hi_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_lo_hi_83 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_50 , core_id_ctrl_decoder_decoded_lo_hi_lo_42 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_lo_83 ={ core_id_ctrl_decoder_decoded_lo_hi_83 , core_id_ctrl_decoder_decoded_lo_lo_78 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_14_37 , core_id_ctrl_decoder_decoded_andMatrixInput_15_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_12_44 , core_id_ctrl_decoder_decoded_andMatrixInput_13_42 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_lo_37 ={ core_id_ctrl_decoder_decoded_hi_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_hi_lo_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_10_47 , core_id_ctrl_decoder_decoded_andMatrixInput_11_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_andMatrixInput_8_65 , core_id_ctrl_decoder_decoded_andMatrixInput_9_50 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_lo_hi_47 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_hi_lo_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_lo_82 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_47 , core_id_ctrl_decoder_decoded_hi_lo_lo_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_lo_3 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_82 , core_id_ctrl_decoder_decoded_andMatrixInput_7_78 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_4_83 , core_id_ctrl_decoder_decoded_andMatrixInput_5_83 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_lo_44 ={ core_id_ctrl_decoder_decoded_hi_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_hi_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_andMatrixInput_2_83 , core_id_ctrl_decoder_decoded_andMatrixInput_3_83 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_hi_9 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_83 , core_id_ctrl_decoder_decoded_andMatrixInput_1_83 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_hi_hi_hi_65 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_hi_9 , core_id_ctrl_decoder_decoded_hi_hi_hi_lo_7 }; 
    wire[7:0] core_id_ctrl_decoder_decoded_hi_hi_83 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_65 , core_id_ctrl_decoder_decoded_hi_hi_lo_44 }; 
    wire[15:0] core_id_ctrl_decoder_decoded_hi_83 ={ core_id_ctrl_decoder_decoded_hi_hi_83 , core_id_ctrl_decoder_decoded_hi_lo_82 }; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_0_84 = core_id_ctrl_decoder_decoded_plaInput [0]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_1_84 = core_id_ctrl_decoder_decoded_plaInput [1]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_2_84 = core_id_ctrl_decoder_decoded_plaInput [2]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_3_84 = core_id_ctrl_decoder_decoded_plaInput [3]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_4_84 = core_id_ctrl_decoder_decoded_invInputs [4]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_5_84 = core_id_ctrl_decoder_decoded_plaInput [5]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_6_83 = core_id_ctrl_decoder_decoded_invInputs [6]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_7_79 = core_id_ctrl_decoder_decoded_plaInput [13]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_8_66 = core_id_ctrl_decoder_decoded_invInputs [14]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_9_51 = core_id_ctrl_decoder_decoded_invInputs [27]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_10_48 = core_id_ctrl_decoder_decoded_invInputs [28]; 
    wire core_id_ctrl_decoder_decoded_andMatrixInput_11_47 = core_id_ctrl_decoder_decoded_plaInput [31]; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_lo_hi_47 ={ core_id_ctrl_decoder_decoded_andMatrixInput_9_51 , core_id_ctrl_decoder_decoded_andMatrixInput_10_48 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_lo_79 ={ core_id_ctrl_decoder_decoded_lo_lo_hi_47 , core_id_ctrl_decoder_decoded_andMatrixInput_11_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_lo_hi_hi_51 ={ core_id_ctrl_decoder_decoded_andMatrixInput_6_83 , core_id_ctrl_decoder_decoded_andMatrixInput_7_79 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_lo_hi_84 ={ core_id_ctrl_decoder_decoded_lo_hi_hi_51 , core_id_ctrl_decoder_decoded_andMatrixInput_8_66 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_lo_84 ={ core_id_ctrl_decoder_decoded_lo_hi_84 , core_id_ctrl_decoder_decoded_lo_lo_79 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_lo_hi_48 ={ core_id_ctrl_decoder_decoded_andMatrixInput_3_84 , core_id_ctrl_decoder_decoded_andMatrixInput_4_84 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_lo_83 ={ core_id_ctrl_decoder_decoded_hi_lo_hi_48 , core_id_ctrl_decoder_decoded_andMatrixInput_5_84 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_hi_hi_hi_66 ={ core_id_ctrl_decoder_decoded_andMatrixInput_0_84 , core_id_ctrl_decoder_decoded_andMatrixInput_1_84 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_hi_hi_84 ={ core_id_ctrl_decoder_decoded_hi_hi_hi_66 , core_id_ctrl_decoder_decoded_andMatrixInput_2_84 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_hi_84 ={ core_id_ctrl_decoder_decoded_hi_hi_84 , core_id_ctrl_decoder_decoded_hi_lo_83 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi ={ core__GEN_36 , core__GEN_49 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi ={&{ core_id_ctrl_decoder_decoded_hi_71 , core_id_ctrl_decoder_decoded_lo_71 },&{ core_id_ctrl_decoder_decoded_hi_75 , core_id_ctrl_decoder_decoded_lo_75 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi ,&{ core_id_ctrl_decoder_decoded_hi_82 , core_id_ctrl_decoder_decoded_lo_82 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi ={&{ core_id_ctrl_decoder_decoded_hi_21 , core_id_ctrl_decoder_decoded_lo_21 }, core__GEN_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi , core__GEN_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo ={ core__GEN_49 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi ={ core__GEN_41 , core__GEN_43 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi , core__GEN_48 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi ={ core__GEN_36 , core__GEN_37 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi , core__GEN_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi ={ core__GEN_30 , core__GEN_34 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi , core__GEN_35 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo }; 
    wire[10:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo ={ core__GEN_27 , core__GEN_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi ={ core__GEN_22 , core__GEN_23 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi , core__GEN_26 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi ={ core__GEN_18 , core__GEN_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi , core__GEN_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi , core__GEN_16 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo }; 
    wire[10:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_3 ={&{ core_id_ctrl_decoder_decoded_hi_61 , core_id_ctrl_decoder_decoded_lo_61 },&{ core_id_ctrl_decoder_decoded_hi_62 , core_id_ctrl_decoder_decoded_lo_62 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_4 ={ core__GEN_20 , core__GEN_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_5 ={ core__GEN_50 , core__GEN_52 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_6 ={ core__GEN_49 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_2 ={ core__GEN_36 , core__GEN_49 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_2 , core__GEN_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_2 ={&{ core_id_ctrl_decoder_decoded_hi_1 , core_id_ctrl_decoder_decoded_lo_1 }, core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_2 , core__GEN_15 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_1 ={&{ core_id_ctrl_decoder_decoded_hi_63 , core_id_ctrl_decoder_decoded_lo_63 },&{ core_id_ctrl_decoder_decoded_hi_66 , core_id_ctrl_decoder_decoded_lo_66 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_1 ={&{ core_id_ctrl_decoder_decoded_hi_51 , core_id_ctrl_decoder_decoded_lo_51 },&{ core_id_ctrl_decoder_decoded_hi_53 , core_id_ctrl_decoder_decoded_lo_53 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_1 ,&{ core_id_ctrl_decoder_decoded_hi_60 , core_id_ctrl_decoder_decoded_lo_60 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_1 ={ core__GEN_40 , core__GEN_41 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_1 , core__GEN_43 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_1 ={ core__GEN_28 , core__GEN_30 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_1 ,&{ core_id_ctrl_decoder_decoded_hi_29 , core_id_ctrl_decoder_decoded_lo_29 }}; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_1 ={ core__GEN_54 , core__GEN_55 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_1 , core__GEN_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_2 ={&{ core_id_ctrl_decoder_decoded_hi_64 , core_id_ctrl_decoder_decoded_lo_64 },&{ core_id_ctrl_decoder_decoded_hi_67 , core_id_ctrl_decoder_decoded_lo_67 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_2 , core__GEN_53 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_2 ={&{ core_id_ctrl_decoder_decoded_hi_55 , core_id_ctrl_decoder_decoded_lo_55 },&{ core_id_ctrl_decoder_decoded_hi_56 , core_id_ctrl_decoder_decoded_lo_56 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_2 ,&{ core_id_ctrl_decoder_decoded_hi_58 , core_id_ctrl_decoder_decoded_lo_58 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_2 ={&{ core_id_ctrl_decoder_decoded_hi_17 , core_id_ctrl_decoder_decoded_lo_17 },&{ core_id_ctrl_decoder_decoded_hi_39 , core_id_ctrl_decoder_decoded_lo_39 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_2 ,&{ core_id_ctrl_decoder_decoded_hi_40 , core_id_ctrl_decoder_decoded_lo_40 }}; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_3 ={&{ core_id_ctrl_decoder_decoded_hi_48 , core_id_ctrl_decoder_decoded_lo_48 }, core__GEN_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_5 ={ core__GEN_39 ,&{ core_id_ctrl_decoder_decoded_hi_45 , core_id_ctrl_decoder_decoded_lo_45 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_3 ={&{ core_id_ctrl_decoder_decoded_hi_41 , core_id_ctrl_decoder_decoded_lo_41 },&{ core_id_ctrl_decoder_decoded_hi_42 , core_id_ctrl_decoder_decoded_lo_42 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_5 ={ core__GEN_35 ,&{ core_id_ctrl_decoder_decoded_hi_35 , core_id_ctrl_decoder_decoded_lo_35 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_6 ={ core__GEN_54 , core__GEN_55 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_6 , core__GEN_56 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_4 ={ core__GEN_39 , core__GEN_53 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_6 ={&{ core_id_ctrl_decoder_decoded_hi_33 , core_id_ctrl_decoder_decoded_lo_33 },&{ core_id_ctrl_decoder_decoded_hi_36 , core_id_ctrl_decoder_decoded_lo_36 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_1 ={ core__GEN_49 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_2 ={ core__GEN_40 ,&{ core_id_ctrl_decoder_decoded_hi_50 , core_id_ctrl_decoder_decoded_lo_50 }}; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_1 ={ core__GEN_37 , core__GEN_39 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_1 ={ core__GEN_32 , core__GEN_35 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_1 , core__GEN_36 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_1 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_1 ={ core__GEN_27 , core__GEN_28 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_3 ={ core__GEN_22 , core__GEN_25 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_1 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_1 ={ core__GEN_19 ,&{ core_id_ctrl_decoder_decoded_hi_12 , core_id_ctrl_decoder_decoded_lo_12 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_1 ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_3 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_1 , core__GEN_15 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_1 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_8 ={ core__GEN_44 , core__GEN_46 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_13 ={ core__GEN_24 , core__GEN_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_3 ={ core__GEN_42 , core__GEN_45 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_3 , core__GEN_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_4 ={ core__GEN_31 , core__GEN_35 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_4 , core__GEN_40 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_4 ={ core__GEN_18 , core__GEN_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_4 , core__GEN_29 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_4 ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_4 , core__GEN_16 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_2 ={ core__GEN_49 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_1 ={ core__GEN_41 , core__GEN_43 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_1 , core__GEN_48 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_2 ={ core__GEN_39 , core__GEN_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_2 ={ core__GEN_35 , core__GEN_36 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_2 , core__GEN_38 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_2 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_2 ={ core__GEN_30 , core__GEN_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_1 ={ core__GEN_23 , core__GEN_25 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_1 , core__GEN_28 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_2 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_1 ={ core__GEN_18 , core__GEN_21 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_1 , core__GEN_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_2 ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_2 , core__GEN_15 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_2 }; 
    wire[10:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_5 ={ core__GEN_42 , core__GEN_45 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_5 , core__GEN_47 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_3 ={ core__GEN_35 , core__GEN_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_6 ={ core__GEN_29 , core__GEN_31 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_7 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_6 ={ core__GEN_19 , core__GEN_26 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_6 , core__GEN_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_3 ={ core__GEN_15 , core__GEN_18 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_6 ={ core__GEN_13 , core__GEN_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_3 }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_16 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_3 ={ core__GEN_46 , core__GEN_48 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_6 ={ core__GEN_43 , core__GEN_44 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_4 ={ core__GEN_40 , core__GEN_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_3 ={ core__GEN_28 , core__GEN_30 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_3 , core__GEN_35 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_4 }; 
    wire[8:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_8 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_3 ={ core__GEN_24 , core__GEN_25 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_2 ={ core__GEN_21 , core__GEN_22 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_2 , core__GEN_23 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_3 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_4 ={ core__GEN_18 , core__GEN_19 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_3 ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_3 , core__GEN_15 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_4 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_4 ={ core__GEN_49 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_2 ={ core__GEN_41 , core__GEN_43 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_2 , core__GEN_48 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_5 ={ core__GEN_39 , core__GEN_40 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_4 ={ core__GEN_35 , core__GEN_36 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_4 , core__GEN_38 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_5 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_9 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_4 ={ core__GEN_30 , core__GEN_33 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_3 ={ core__GEN_23 , core__GEN_25 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_3 , core__GEN_28 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_4 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_2 ={ core__GEN_18 , core__GEN_21 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_2 , core__GEN_22 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_4 ={ core__GEN_13 , core__GEN_14 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_8 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_4 , core__GEN_15 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_5 }; 
    wire[10:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_18 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_8 ={ core__GEN_48 , core__GEN_49 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_8 , core__GEN_50 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_9 ={ core__GEN_36 , core__GEN_39 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_9 , core__GEN_43 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_10 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_9 ={ core__GEN_22 , core__GEN_23 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_9 ,&{ core_id_ctrl_decoder_decoded_hi_15 , core_id_ctrl_decoder_decoded_lo_15 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_9 ={ core__GEN_20 ,&{ core_id_ctrl_decoder_decoded_hi_10 , core_id_ctrl_decoder_decoded_lo_10 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_9 , core__GEN_21 }; 
    wire[5:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_19 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi ={&{ core_id_ctrl_decoder_decoded_hi_72 , core_id_ctrl_decoder_decoded_lo_72 },&{ core_id_ctrl_decoder_decoded_hi_76 , core_id_ctrl_decoder_decoded_lo_76 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi ,&{ core_id_ctrl_decoder_decoded_hi_83 , core_id_ctrl_decoder_decoded_lo_83 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo ={ core__GEN_49 , core__GEN_51 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_3 ={ core__GEN_43 , core__GEN_48 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_9 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_3 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_1 ={ core__GEN_39 , core__GEN_40 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_1 , core__GEN_41 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo ={ core__GEN_36 , core__GEN_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_5 ={ core__GEN_32 , core__GEN_35 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_6 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_11 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi ={&{ core_id_ctrl_decoder_decoded_hi_22 , core_id_ctrl_decoder_decoded_lo_22 }, core__GEN_28 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi , core__GEN_30 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo ={ core__GEN_25 , core__GEN_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_4 ={ core__GEN_22 , core__GEN_23 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_5 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_3 ={ core__GEN_18 , core__GEN_19 }; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_3 , core__GEN_21 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo ={ core__GEN_15 , core__GEN_17 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_5 ={ core__GEN_13 , core__GEN_14 }; 
    wire[3:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo }; 
    wire[6:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_14 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_6 }; 
    wire[13:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_20 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi , core__GEN_50 },1'h0}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ={| core__GEN_34 ,|(&{ core_id_ctrl_decoder_decoded_hi_23 , core_id_ctrl_decoder_decoded_lo_23 })}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ,| core__GEN_17 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo_1 ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo },| core__GEN_37 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ={1'h0,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_3 , core__GEN_48 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_1 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_10 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_lo_1 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_12 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_4 ,&{ core_id_ctrl_decoder_decoded_hi_74 , core_id_ctrl_decoder_decoded_lo_74 }},1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_2 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ,1'h0}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_hi_2 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo_1 ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_6 ,&{ core_id_ctrl_decoder_decoded_hi_84 , core_id_ctrl_decoder_decoded_lo_84 }},|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_5 ,&{ core_id_ctrl_decoder_decoded_hi_78 , core_id_ctrl_decoder_decoded_lo_78 }}}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_7 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_2 },1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ,| core__GEN_36 }; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_lo_1 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_lo_7 }; 
    wire[19:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_hi_15 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_lo_12 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_9 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_4 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_8 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_3 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_12 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_7 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_6 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_1 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_10 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_5 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_hi_1 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo_1 ={|{ core__GEN_19 , core__GEN_27 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_13 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_8 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ={|{&{ core_id_ctrl_decoder_decoded_hi_8 , core_id_ctrl_decoder_decoded_lo_8 }, core__GEN_27 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_15 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_10 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_5 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_14 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_9 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_hi_5 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_lo_1 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_13 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_lo_6 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_lo ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_17 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_12 },|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_16 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_11 }}; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ={| core__GEN_26 ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_19 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_14 }}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_4 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ,|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_18 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_13 }}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_7 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_hi_4 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo_1 ={|{ core__GEN_24 , core__GEN_39 },| core__GEN_27 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ={|{ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_20 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_15 },1'h0}; 
    wire[2:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_6 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ,1'h0}; 
    wire[4:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_11 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_hi_6 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_lo_1 }; 
    wire[9:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_hi_11 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_lo_7 }; 
    wire[19:0] core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_21 ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_hi_15 , core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_lo_13 }; 
    wire[39:0] core_id_ctrl_decoder_decoded_orMatrixOutputs ={ core_id_ctrl_decoder_decoded_orMatrixOutputs_hi_21 , core_id_ctrl_decoder_decoded_orMatrixOutputs_lo_16 }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [1], core_id_ctrl_decoder_decoded_orMatrixOutputs [0]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [4], core_id_ctrl_decoder_decoded_orMatrixOutputs [3]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [2]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [6], core_id_ctrl_decoder_decoded_orMatrixOutputs [5]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [9], core_id_ctrl_decoder_decoded_orMatrixOutputs [8]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [7]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [11], core_id_ctrl_decoder_decoded_orMatrixOutputs [10]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [14], core_id_ctrl_decoder_decoded_orMatrixOutputs [13]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [12]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [16], core_id_ctrl_decoder_decoded_orMatrixOutputs [15]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [19], core_id_ctrl_decoder_decoded_orMatrixOutputs [18]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [17]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi_lo }; 
    wire[19:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [21], core_id_ctrl_decoder_decoded_orMatrixOutputs [20]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [24], core_id_ctrl_decoder_decoded_orMatrixOutputs [23]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [22]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [26], core_id_ctrl_decoder_decoded_orMatrixOutputs [25]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [29], core_id_ctrl_decoder_decoded_orMatrixOutputs [28]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [27]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [31], core_id_ctrl_decoder_decoded_orMatrixOutputs [30]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [34], core_id_ctrl_decoder_decoded_orMatrixOutputs [33]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [32]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_lo ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [36], core_id_ctrl_decoder_decoded_orMatrixOutputs [35]}; 
    wire[1:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_orMatrixOutputs [39], core_id_ctrl_decoder_decoded_orMatrixOutputs [38]}; 
    wire[2:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_orMatrixOutputs [37]}; 
    wire[4:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi_lo }; 
    wire[9:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi_lo }; 
    wire[19:0] core_id_ctrl_decoder_decoded_invMatrixOutputs_hi ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_id_ctrl_decoder_decoded_invMatrixOutputs ={ core_id_ctrl_decoder_decoded_invMatrixOutputs_hi , core_id_ctrl_decoder_decoded_invMatrixOutputs_lo }; 
    wire[39:0] core_id_ctrl_decoder_decoded = core_id_ctrl_decoder_decoded_invMatrixOutputs ; 
  assign  core_id_ctrl_decoder_0 = core_id_ctrl_decoder_decoded [39]; 
    wire core_id_ctrl_legal = core_id_ctrl_decoder_0 ; 
  assign  core_id_ctrl_decoder_1 = core_id_ctrl_decoder_decoded [38]; 
    wire core_id_ctrl_fp = core_id_ctrl_decoder_1 ; 
  assign  core_id_ctrl_decoder_2 = core_id_ctrl_decoder_decoded [37]; 
    wire core_id_ctrl_rocc = core_id_ctrl_decoder_2 ; 
  assign  core_id_ctrl_decoder_3 = core_id_ctrl_decoder_decoded [36]; 
    wire core_id_ctrl_branch = core_id_ctrl_decoder_3 ; 
  assign  core_id_ctrl_decoder_4 = core_id_ctrl_decoder_decoded [35]; 
    wire core_id_ctrl_jal = core_id_ctrl_decoder_4 ; 
  assign  core_id_ctrl_decoder_5 = core_id_ctrl_decoder_decoded [34]; 
    wire core_id_ctrl_jalr = core_id_ctrl_decoder_5 ; 
  assign  core_id_ctrl_decoder_6 = core_id_ctrl_decoder_decoded [33]; 
    wire core_id_ctrl_rxs2 = core_id_ctrl_decoder_6 ; 
  assign  core_id_ctrl_decoder_7 = core_id_ctrl_decoder_decoded [32]; 
    wire core_id_ctrl_rxs1 = core_id_ctrl_decoder_7 ; 
  assign  core_id_ctrl_decoder_8 = core_id_ctrl_decoder_decoded [31:30]; 
    wire[1:0] core_id_ctrl_sel_alu2 = core_id_ctrl_decoder_8 ; 
  assign  core_id_ctrl_decoder_9 = core_id_ctrl_decoder_decoded [29:28]; 
    wire[1:0] core_id_ctrl_sel_alu1 = core_id_ctrl_decoder_9 ; 
  assign  core_id_ctrl_decoder_10 = core_id_ctrl_decoder_decoded [27:25]; 
    wire[2:0] core_id_ctrl_sel_imm = core_id_ctrl_decoder_10 ; 
  assign  core_id_ctrl_decoder_11 = core_id_ctrl_decoder_decoded [24]; 
    wire core_id_ctrl_alu_dw = core_id_ctrl_decoder_11 ; 
  assign  core_id_ctrl_decoder_12 = core_id_ctrl_decoder_decoded [23:20]; 
    wire[3:0] core_id_ctrl_alu_fn = core_id_ctrl_decoder_12 ; 
  assign  core_id_ctrl_decoder_13 = core_id_ctrl_decoder_decoded [19]; 
    wire core_id_ctrl_mem = core_id_ctrl_decoder_13 ; 
  assign  core_id_ctrl_decoder_14 = core_id_ctrl_decoder_decoded [18:14]; 
    wire[4:0] core_id_ctrl_mem_cmd = core_id_ctrl_decoder_14 ; 
  assign  core_id_ctrl_decoder_15 = core_id_ctrl_decoder_decoded [13]; 
    wire core_id_ctrl_rfs1 = core_id_ctrl_decoder_15 ; 
  assign  core_id_ctrl_decoder_16 = core_id_ctrl_decoder_decoded [12]; 
    wire core_id_ctrl_rfs2 = core_id_ctrl_decoder_16 ; 
  assign  core_id_ctrl_decoder_17 = core_id_ctrl_decoder_decoded [11]; 
    wire core_id_ctrl_rfs3 = core_id_ctrl_decoder_17 ; 
  assign  core_id_ctrl_decoder_18 = core_id_ctrl_decoder_decoded [10]; 
    wire core_id_ctrl_wfd = core_id_ctrl_decoder_18 ; 
  assign  core_id_ctrl_decoder_19 = core_id_ctrl_decoder_decoded [9]; 
    wire core_id_ctrl_mul = core_id_ctrl_decoder_19 ; 
  assign  core_id_ctrl_decoder_20 = core_id_ctrl_decoder_decoded [8]; 
    wire core_id_ctrl_div = core_id_ctrl_decoder_20 ; 
  assign  core_id_ctrl_decoder_21 = core_id_ctrl_decoder_decoded [7]; 
    wire core_id_ctrl_wxd = core_id_ctrl_decoder_21 ; 
  assign  core_id_ctrl_decoder_22 = core_id_ctrl_decoder_decoded [6:4]; 
    wire[2:0] core_id_ctrl_csr = core_id_ctrl_decoder_22 ; 
  assign  core_id_ctrl_decoder_23 = core_id_ctrl_decoder_decoded [3]; 
    wire core_id_ctrl_fence_i = core_id_ctrl_decoder_23 ; 
  assign  core_id_ctrl_decoder_24 = core_id_ctrl_decoder_decoded [2]; 
    wire core_id_ctrl_fence = core_id_ctrl_decoder_24 ; 
  assign  core_id_ctrl_decoder_25 = core_id_ctrl_decoder_decoded [1]; 
    wire core_id_ctrl_amo = core_id_ctrl_decoder_25 ; 
  assign  core_id_ctrl_decoder_26 = core_id_ctrl_decoder_decoded [0]; 
    wire core_id_ctrl_dp = core_id_ctrl_decoder_26 ; 
    reg core_id_reg_fence ; 
    wire[63:0] core_rf_wdata ;  
    wire[4:0] core_rf_ext_R0_addr;
    wire core_rf_ext_R0_en;
    wire core_rf_ext_R0_clk;
    wire[63:0] core_rf_ext_R0_data;
    wire[4:0] core_rf_ext_R1_addr;
    wire core_rf_ext_R1_en;
    wire core_rf_ext_R1_clk;
    wire[63:0] core_rf_ext_R1_data;
    wire[4:0] core_rf_ext_W0_addr;
    wire core_rf_ext_W0_en;
    wire core_rf_ext_W0_clk;
    wire[63:0] core_rf_ext_W0_data;

    reg[63:0] core_rf_ext_Memory [0:30]; 
  always @( posedge  core_rf_ext_W0_clk )
         begin 
             if ( core_rf_ext_W0_en &1'h1) 
                 core_rf_ext_Memory  [ core_rf_ext_W0_addr ]<= core_rf_ext_W0_data ;
         end
  assign  core_rf_ext_R0_data = core_rf_ext_R0_en  ?  core_rf_ext_Memory [ core_rf_ext_R0_addr ]:64'bx; 
  assign  core_rf_ext_R1_data = core_rf_ext_R1_en  ?  core_rf_ext_Memory [ core_rf_ext_R1_addr ]:64'bx;
    assign core_rf_ext_R0_addr = core__GEN_10;
    assign core_rf_ext_R0_en = 1'h1;
    assign core_rf_ext_R0_clk = core_clock;
    assign core__rf_ext_R0_data = core_rf_ext_R0_data;
    assign core_rf_ext_R1_addr = core__GEN_11;
    assign core_rf_ext_R1_en = 1'h1;
    assign core_rf_ext_R1_clk = core_clock;
    assign core__rf_ext_R1_data = core_rf_ext_R1_data;
    assign core_rf_ext_W0_addr = core__GEN_6;
    assign core_rf_ext_W0_en = core__GEN_12;
    assign core_rf_ext_W0_clk = core_clock;
    assign core_rf_ext_W0_data = core_rf_wdata;
     
  assign  core__GEN_12 = core__GEN_5 &1'h1; 
  assign  core__GEN_11 =~ core_id_raddr1 ; 
  assign  core__GEN_10 =~ core_id_raddr2 ; 
    wire core_id_npc_sign = core__ibuf_io_inst_0_bits_inst_bits [31]; 
    wire core_id_npc_hi_hi_hi = core_id_npc_sign ; 
    wire[10:0] core_id_npc_b30_20 ={{10{ core_id_npc_sign }}, core_id_npc_sign }; 
    wire[10:0] core_id_npc_hi_hi_lo = core_id_npc_b30_20 ; 
    wire[7:0] core_id_npc_b19_12 = core__ibuf_io_inst_0_bits_inst_bits [19:12]; 
    wire[7:0] core_id_npc_hi_lo_hi = core_id_npc_b19_12 ; 
    wire core_id_npc_b11 = core__ibuf_io_inst_0_bits_inst_bits [20]; 
    wire core_id_npc_hi_lo_lo = core_id_npc_b11 ; 
    wire[5:0] core_id_npc_b10_5 = core__ibuf_io_inst_0_bits_inst_bits [30:25]; 
    wire[3:0] core_id_npc_b4_1 = core__ibuf_io_inst_0_bits_inst_bits [24:21]; 
    wire[9:0] core_id_npc_lo_hi ={ core_id_npc_b10_5 , core_id_npc_b4_1 }; 
    wire[10:0] core_id_npc_lo ={ core_id_npc_lo_hi , core_id_npc_b0 }; 
    wire[8:0] core_id_npc_hi_lo ={ core_id_npc_hi_lo_hi , core_id_npc_hi_lo_lo }; 
    wire[11:0] core_id_npc_hi_hi ={ core_id_npc_hi_hi_hi , core_id_npc_hi_hi_lo }; 
    wire[20:0] core_id_npc_hi ={ core_id_npc_hi_hi , core_id_npc_hi_lo }; 
    wire[31:0] core__GEN_57 ={ core_id_npc_hi , core_id_npc_lo }; 
    wire[34:0] core__GEN_58 ={ core__ibuf_io_pc [33], core__ibuf_io_pc }+{{3{ core__GEN_57 [31]}}, core__GEN_57 }; 
    wire[33:0] core_id_npc = core__GEN_58 [33:0]; 
    wire core_wb_xcpt ; 
    wire[63:0] core_wb_cause ; 
    wire core_wb_valid ;  
    wire core_csr_clock;
    wire core_csr_reset;
    wire core_csr_io_ungated_clock;
    wire core_csr_io_interrupts_debug;
    wire core_csr_io_interrupts_mtip;
    wire core_csr_io_interrupts_msip;
    wire core_csr_io_interrupts_meip;
    wire core_csr_io_hartid;
    wire[11:0] core_csr_io_rw_addr;
    wire[2:0] core_csr_io_rw_cmd;
    wire[63:0] core_csr_io_rw_rdata;
    wire[63:0] core_csr_io_rw_wdata;
    wire[31:0] core_csr_io_decode_0_inst;
    wire core_csr_io_decode_0_fp_illegal;
    wire core_csr_io_decode_0_vector_illegal;
    wire core_csr_io_decode_0_fp_csr;
    wire core_csr_io_decode_0_rocc_illegal;
    wire core_csr_io_decode_0_read_illegal;
    wire core_csr_io_decode_0_write_illegal;
    wire core_csr_io_decode_0_write_flush;
    wire core_csr_io_decode_0_system_illegal;
    wire core_csr_io_decode_0_virtual_access_illegal;
    wire core_csr_io_decode_0_virtual_system_illegal;
    wire core_csr_io_csr_stall;
    wire core_csr_io_rw_stall;
    wire core_csr_io_eret;
    wire core_csr_io_singleStep;
    wire core_csr_io_status_debug;
    wire core_csr_io_status_cease;
    wire core_csr_io_status_wfi;
    wire[31:0] core_csr_io_status_isa;
    wire[1:0] core_csr_io_status_dprv;
    wire core_csr_io_status_dv;
    wire[1:0] core_csr_io_status_prv;
    wire core_csr_io_status_v;
    wire core_csr_io_status_sd;
    wire[22:0] core_csr_io_status_zero2;
    wire core_csr_io_status_mpv;
    wire core_csr_io_status_gva;
    wire core_csr_io_status_mbe;
    wire core_csr_io_status_sbe;
    wire[1:0] core_csr_io_status_sxl;
    wire[1:0] core_csr_io_status_uxl;
    wire core_csr_io_status_sd_rv32;
    wire[7:0] core_csr_io_status_zero1;
    wire core_csr_io_status_tsr;
    wire core_csr_io_status_tw;
    wire core_csr_io_status_tvm;
    wire core_csr_io_status_mxr;
    wire core_csr_io_status_sum;
    wire core_csr_io_status_mprv;
    wire[1:0] core_csr_io_status_xs;
    wire[1:0] core_csr_io_status_fs;
    wire[1:0] core_csr_io_status_mpp;
    wire[1:0] core_csr_io_status_vs;
    wire core_csr_io_status_spp;
    wire core_csr_io_status_mpie;
    wire core_csr_io_status_ube;
    wire core_csr_io_status_spie;
    wire core_csr_io_status_upie;
    wire core_csr_io_status_mie;
    wire core_csr_io_status_hie;
    wire core_csr_io_status_sie;
    wire core_csr_io_status_uie;
    wire[29:0] core_csr_io_hstatus_zero6;
    wire[1:0] core_csr_io_hstatus_vsxl;
    wire[8:0] core_csr_io_hstatus_zero5;
    wire core_csr_io_hstatus_vtsr;
    wire core_csr_io_hstatus_vtw;
    wire core_csr_io_hstatus_vtvm;
    wire[1:0] core_csr_io_hstatus_zero3;
    wire[5:0] core_csr_io_hstatus_vgein;
    wire[1:0] core_csr_io_hstatus_zero2;
    wire core_csr_io_hstatus_hu;
    wire core_csr_io_hstatus_spvp;
    wire core_csr_io_hstatus_spv;
    wire core_csr_io_hstatus_gva;
    wire core_csr_io_hstatus_vsbe;
    wire[4:0] core_csr_io_hstatus_zero1;
    wire core_csr_io_gstatus_debug;
    wire core_csr_io_gstatus_cease;
    wire core_csr_io_gstatus_wfi;
    wire[31:0] core_csr_io_gstatus_isa;
    wire[1:0] core_csr_io_gstatus_dprv;
    wire core_csr_io_gstatus_dv;
    wire[1:0] core_csr_io_gstatus_prv;
    wire core_csr_io_gstatus_v;
    wire core_csr_io_gstatus_sd;
    wire[22:0] core_csr_io_gstatus_zero2;
    wire core_csr_io_gstatus_mpv;
    wire core_csr_io_gstatus_gva;
    wire core_csr_io_gstatus_mbe;
    wire core_csr_io_gstatus_sbe;
    wire[1:0] core_csr_io_gstatus_sxl;
    wire[1:0] core_csr_io_gstatus_uxl;
    wire core_csr_io_gstatus_sd_rv32;
    wire[7:0] core_csr_io_gstatus_zero1;
    wire core_csr_io_gstatus_tsr;
    wire core_csr_io_gstatus_tw;
    wire core_csr_io_gstatus_tvm;
    wire core_csr_io_gstatus_mxr;
    wire core_csr_io_gstatus_sum;
    wire core_csr_io_gstatus_mprv;
    wire[1:0] core_csr_io_gstatus_xs;
    wire[1:0] core_csr_io_gstatus_fs;
    wire[1:0] core_csr_io_gstatus_mpp;
    wire[1:0] core_csr_io_gstatus_vs;
    wire core_csr_io_gstatus_spp;
    wire core_csr_io_gstatus_mpie;
    wire core_csr_io_gstatus_ube;
    wire core_csr_io_gstatus_spie;
    wire core_csr_io_gstatus_upie;
    wire core_csr_io_gstatus_mie;
    wire core_csr_io_gstatus_hie;
    wire core_csr_io_gstatus_sie;
    wire core_csr_io_gstatus_uie;
    wire[3:0] core_csr_io_ptbr_mode;
    wire[15:0] core_csr_io_ptbr_asid;
    wire[43:0] core_csr_io_ptbr_ppn;
    wire[3:0] core_csr_io_hgatp_mode;
    wire[15:0] core_csr_io_hgatp_asid;
    wire[43:0] core_csr_io_hgatp_ppn;
    wire[3:0] core_csr_io_vsatp_mode;
    wire[15:0] core_csr_io_vsatp_asid;
    wire[43:0] core_csr_io_vsatp_ppn;
    wire[33:0] core_csr_io_evec;
    wire core_csr_io_exception;
    wire core_csr_io_retire;
    wire[63:0] core_csr_io_cause;
    wire[33:0] core_csr_io_pc;
    wire[33:0] core_csr_io_tval;
    wire[39:0] core_csr_io_htval;
    wire core_csr_io_gva;
    wire[63:0] core_csr_io_time;
    wire[2:0] core_csr_io_fcsr_rm;
    wire core_csr_io_fcsr_flags_valid;
    wire[4:0] core_csr_io_fcsr_flags_bits;
    wire core_csr_io_rocc_interrupt;
    wire core_csr_io_interrupt;
    wire[63:0] core_csr_io_interrupt_cause;
    wire[3:0] core_csr_io_bp_0_control_ttype;
    wire core_csr_io_bp_0_control_dmode;
    wire[5:0] core_csr_io_bp_0_control_maskmax;
    wire[39:0] core_csr_io_bp_0_control_reserved;
    wire core_csr_io_bp_0_control_action;
    wire core_csr_io_bp_0_control_chain;
    wire[1:0] core_csr_io_bp_0_control_zero;
    wire[1:0] core_csr_io_bp_0_control_tmatch;
    wire core_csr_io_bp_0_control_m;
    wire core_csr_io_bp_0_control_h;
    wire core_csr_io_bp_0_control_s;
    wire core_csr_io_bp_0_control_u;
    wire core_csr_io_bp_0_control_x;
    wire core_csr_io_bp_0_control_w;
    wire core_csr_io_bp_0_control_r;
    wire[32:0] core_csr_io_bp_0_address;
    wire core_csr_io_bp_0_textra_mselect;
    wire[47:0] core_csr_io_bp_0_textra_pad2;
    wire core_csr_io_bp_0_textra_pad1;
    wire core_csr_io_bp_0_textra_sselect;
    wire core_csr_io_pmp_0_cfg_l;
    wire[1:0] core_csr_io_pmp_0_cfg_res;
    wire[1:0] core_csr_io_pmp_0_cfg_a;
    wire core_csr_io_pmp_0_cfg_x;
    wire core_csr_io_pmp_0_cfg_w;
    wire core_csr_io_pmp_0_cfg_r;
    wire[29:0] core_csr_io_pmp_0_addr;
    wire[31:0] core_csr_io_pmp_0_mask;
    wire core_csr_io_pmp_1_cfg_l;
    wire[1:0] core_csr_io_pmp_1_cfg_res;
    wire[1:0] core_csr_io_pmp_1_cfg_a;
    wire core_csr_io_pmp_1_cfg_x;
    wire core_csr_io_pmp_1_cfg_w;
    wire core_csr_io_pmp_1_cfg_r;
    wire[29:0] core_csr_io_pmp_1_addr;
    wire[31:0] core_csr_io_pmp_1_mask;
    wire core_csr_io_pmp_2_cfg_l;
    wire[1:0] core_csr_io_pmp_2_cfg_res;
    wire[1:0] core_csr_io_pmp_2_cfg_a;
    wire core_csr_io_pmp_2_cfg_x;
    wire core_csr_io_pmp_2_cfg_w;
    wire core_csr_io_pmp_2_cfg_r;
    wire[29:0] core_csr_io_pmp_2_addr;
    wire[31:0] core_csr_io_pmp_2_mask;
    wire core_csr_io_pmp_3_cfg_l;
    wire[1:0] core_csr_io_pmp_3_cfg_res;
    wire[1:0] core_csr_io_pmp_3_cfg_a;
    wire core_csr_io_pmp_3_cfg_x;
    wire core_csr_io_pmp_3_cfg_w;
    wire core_csr_io_pmp_3_cfg_r;
    wire[29:0] core_csr_io_pmp_3_addr;
    wire[31:0] core_csr_io_pmp_3_mask;
    wire core_csr_io_pmp_4_cfg_l;
    wire[1:0] core_csr_io_pmp_4_cfg_res;
    wire[1:0] core_csr_io_pmp_4_cfg_a;
    wire core_csr_io_pmp_4_cfg_x;
    wire core_csr_io_pmp_4_cfg_w;
    wire core_csr_io_pmp_4_cfg_r;
    wire[29:0] core_csr_io_pmp_4_addr;
    wire[31:0] core_csr_io_pmp_4_mask;
    wire core_csr_io_pmp_5_cfg_l;
    wire[1:0] core_csr_io_pmp_5_cfg_res;
    wire[1:0] core_csr_io_pmp_5_cfg_a;
    wire core_csr_io_pmp_5_cfg_x;
    wire core_csr_io_pmp_5_cfg_w;
    wire core_csr_io_pmp_5_cfg_r;
    wire[29:0] core_csr_io_pmp_5_addr;
    wire[31:0] core_csr_io_pmp_5_mask;
    wire core_csr_io_pmp_6_cfg_l;
    wire[1:0] core_csr_io_pmp_6_cfg_res;
    wire[1:0] core_csr_io_pmp_6_cfg_a;
    wire core_csr_io_pmp_6_cfg_x;
    wire core_csr_io_pmp_6_cfg_w;
    wire core_csr_io_pmp_6_cfg_r;
    wire[29:0] core_csr_io_pmp_6_addr;
    wire[31:0] core_csr_io_pmp_6_mask;
    wire core_csr_io_pmp_7_cfg_l;
    wire[1:0] core_csr_io_pmp_7_cfg_res;
    wire[1:0] core_csr_io_pmp_7_cfg_a;
    wire core_csr_io_pmp_7_cfg_x;
    wire core_csr_io_pmp_7_cfg_w;
    wire core_csr_io_pmp_7_cfg_r;
    wire[29:0] core_csr_io_pmp_7_addr;
    wire[31:0] core_csr_io_pmp_7_mask;
    wire[31:0] core_csr_io_csrw_counter;
    wire core_csr_io_inhibit_cycle;
    wire[31:0] core_csr_io_inst_0;
    wire core_csr_io_trace_0_valid;
    wire[33:0] core_csr_io_trace_0_iaddr;
    wire[31:0] core_csr_io_trace_0_insn;
    wire[2:0] core_csr_io_trace_0_priv;
    wire core_csr_io_trace_0_exception;
    wire core_csr_io_trace_0_interrupt;
    wire[63:0] core_csr_io_trace_0_cause;
    wire[33:0] core_csr_io_trace_0_tval;
    wire core_csr_io_fiom;
    wire core_csr_io_customCSRs_0_ren;
    wire core_csr_io_customCSRs_0_wen;
    wire[63:0] core_csr_io_customCSRs_0_wdata;
    wire[63:0] core_csr_io_customCSRs_0_value;
    wire core_csr_io_customCSRs_0_stall;
    wire core_csr_io_customCSRs_0_set;
    wire[63:0] core_csr_io_customCSRs_0_sdata;
    wire core_csr_io_customCSRs_1_ren;
    wire core_csr_io_customCSRs_1_wen;
    wire[63:0] core_csr_io_customCSRs_1_wdata;
    wire[63:0] core_csr_io_customCSRs_1_value;
    wire core_csr_io_customCSRs_1_stall;
    wire core_csr_io_customCSRs_1_set;
    wire[63:0] core_csr_io_customCSRs_1_sdata;
    wire core_csr_io_customCSRs_2_ren;
    wire core_csr_io_customCSRs_2_wen;
    wire[63:0] core_csr_io_customCSRs_2_wdata;
    wire[63:0] core_csr_io_customCSRs_2_value;
    wire core_csr_io_customCSRs_2_stall;
    wire core_csr_io_customCSRs_2_set;
    wire[63:0] core_csr_io_customCSRs_2_sdata;
    wire core_csr_io_customCSRs_3_ren;
    wire core_csr_io_customCSRs_3_wen;
    wire[63:0] core_csr_io_customCSRs_3_wdata;
    wire[63:0] core_csr_io_customCSRs_3_value;
    wire core_csr_io_customCSRs_3_stall;
    wire core_csr_io_customCSRs_3_set;
    wire[63:0] core_csr_io_customCSRs_3_sdata;

    wire core_csr_mip_rocc = core_csr_io_rocc_interrupt ; 
    wire core_csr_mip_meip = core_csr_io_interrupts_meip ; 
    wire core_csr_mip_mtip = core_csr_io_interrupts_mtip ; 
    wire core_csr_mip_msip = core_csr_io_interrupts_msip ; 
    wire[31:0] core_csr_decoded_plaInput_1 = core_csr_io_decode_0_inst ; 
    wire core_csr_set_fs_dirty = core_csr_io_fcsr_flags_valid ; 
    wire[39:0] core_csr__reg_bp_1_WIRE_control_reserved =40'h0; 
    wire[3:0] core_csr__reg_bp_1_WIRE_control_ttype =4'h0; 
    wire[32:0] core_csr__reg_bp_1_WIRE_address =33'h0; 
    wire[29:0] core_csr__reg_hstatus_WIRE_zero6 =30'h0; 
    wire[29:0] core_csr_read_pmp_15_addr =30'h0; 
    wire[8:0] core_csr__reg_hstatus_WIRE_zero5 =9'h0; 
    wire[5:0] core_csr__reg_hstatus_WIRE_vgein =6'h0; 
    wire[5:0] core_csr__reg_bp_1_WIRE_control_maskmax =6'h0; 
    wire[4:0] core_csr__reg_hstatus_WIRE_zero1 =5'h0; 
    wire[53:0] core_csr__reg_menvcfg_WIRE_zero54 =54'h0; 
    wire[53:0] core_csr__reg_senvcfg_WIRE_zero54 =54'h0; 
    wire[53:0] core_csr__reg_henvcfg_WIRE_zero54 =54'h0; 
    wire[63:0] core_csr_read_mideleg =64'h0; 
    wire[63:0] core_csr_read_medeleg =64'h0; 
    wire[63:0] core_csr_read_hideleg =64'h0; 
    wire[63:0] core_csr_read_hedeleg =64'h0; 
    wire[47:0] core_csr__reg_bp_1_WIRE_textra_pad2 =48'h0; 
    wire core_csr_sup_meip =1'h1; 
    wire core_csr_sup_mtip =1'h1; 
    wire core_csr_sup_msip =1'h1; 
    wire core_csr_sie_mask_sgeip_mask_sgeip =1'h1; 
    wire core_csr_allow_wfi =1'h1; 
    wire core_csr_allow_sfence_vma =1'h1; 
    wire core_csr_allow_hfence_vvma =1'h1; 
    wire core_csr_allow_hlsv =1'h1; 
    wire core_csr_allow_sret =1'h1; 
    wire core_csr_delegable_16 =1'h1; 
    wire core_csr_delegable_18 =1'h1; 
    wire core_csr_delegable_19 =1'h1; 
    wire core_csr_delegable_20 =1'h1; 
    wire core_csr_delegable_22 =1'h1; 
    wire[11:0] core_csr__reset_dcsr_WIRE_zero3 =12'h0; 
    wire[2:0] core_csr__reset_dcsr_WIRE_cause =3'h0; 
    wire[2:0] core_csr__reset_mnstatus_WIRE_zero3 =3'h0; 
    wire[2:0] core_csr__reset_mnstatus_WIRE_zero2 =3'h0; 
    wire[2:0] core_csr__reset_mnstatus_WIRE_zero1 =3'h0; 
    wire[2:0] core_csr__reg_menvcfg_WIRE_zero3 =3'h0; 
    wire[2:0] core_csr__reg_senvcfg_WIRE_zero3 =3'h0; 
    wire[2:0] core_csr__reg_henvcfg_WIRE_zero3 =3'h0; 
    wire[2:0] core_csr__read_mnstatus_WIRE_zero3 =3'h0; 
    wire[2:0] core_csr__read_mnstatus_WIRE_zero2 =3'h0; 
    wire[2:0] core_csr__read_mnstatus_WIRE_zero1 =3'h0; 
    wire[1:0] core_csr_reset_mstatus_prv =2'h3; 
    wire[1:0] core_csr_reset_mstatus_mpp =2'h3; 
    wire[1:0] core_csr_reset_dcsr_prv =2'h3; 
    wire[1:0] core_csr_reset_mnstatus_mpp =2'h3; 
    wire[31:0] core_csr__reset_mstatus_WIRE_isa =32'h0; 
    wire[31:0] core_csr_read_mcounteren =32'h0; 
    wire[31:0] core_csr_read_scounteren =32'h0; 
    wire[31:0] core_csr_read_hcounteren =32'h0; 
    wire[31:0] core_csr_read_pmp_15_mask =32'h0; 
    wire[22:0] core_csr__reset_mstatus_WIRE_zero2 =23'h0; 
    wire[7:0] core_csr__reset_mstatus_WIRE_zero1 =8'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_dprv =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_prv =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_sxl =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_uxl =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_xs =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_fs =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_mpp =2'h0; 
    wire[1:0] core_csr__reset_mstatus_WIRE_vs =2'h0; 
    wire[1:0] core_csr__reset_dcsr_WIRE_xdebugver =2'h0; 
    wire[1:0] core_csr__reset_dcsr_WIRE_zero4 =2'h0; 
    wire[1:0] core_csr__reset_dcsr_WIRE_zero1 =2'h0; 
    wire[1:0] core_csr__reset_dcsr_WIRE_prv =2'h0; 
    wire[1:0] core_csr__reset_mnstatus_WIRE_mpp =2'h0; 
    wire[1:0] core_csr__reg_menvcfg_WIRE_cbie =2'h0; 
    wire[1:0] core_csr__reg_senvcfg_WIRE_cbie =2'h0; 
    wire[1:0] core_csr__reg_henvcfg_WIRE_cbie =2'h0; 
    wire[1:0] core_csr__reg_hstatus_WIRE_vsxl =2'h0; 
    wire[1:0] core_csr__reg_hstatus_WIRE_zero3 =2'h0; 
    wire[1:0] core_csr__reg_hstatus_WIRE_zero2 =2'h0; 
    wire[1:0] core_csr__read_mnstatus_WIRE_mpp =2'h0; 
    wire[1:0] core_csr_read_vcsr =2'h0; 
    wire[1:0] core_csr_read_pmp_15_cfg_res =2'h0; 
    wire[1:0] core_csr_read_pmp_15_cfg_a =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_lo =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_hi =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_lo_1 =2'h0; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_lo_hi_1 =2'h0; 
    wire[1:0] core_csr_nmiTVec =2'h0; 
    wire[1:0] core_csr__reg_bp_1_WIRE_control_zero =2'h0; 
    wire[1:0] core_csr__reg_bp_1_WIRE_control_tmatch =2'h0; 
    wire core_csr__io_status_sd_rv32_output =1'h0; 
    wire core_csr__reset_mstatus_WIRE_debug =1'h0; 
    wire core_csr__reset_mstatus_WIRE_cease =1'h0; 
    wire core_csr__reset_mstatus_WIRE_wfi =1'h0; 
    wire core_csr__reset_mstatus_WIRE_dv =1'h0; 
    wire core_csr__reset_mstatus_WIRE_v =1'h0; 
    wire core_csr__reset_mstatus_WIRE_sd =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mpv =1'h0; 
    wire core_csr__reset_mstatus_WIRE_gva =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mbe =1'h0; 
    wire core_csr__reset_mstatus_WIRE_sbe =1'h0; 
    wire core_csr__reset_mstatus_WIRE_sd_rv32 =1'h0; 
    wire core_csr__reset_mstatus_WIRE_tsr =1'h0; 
    wire core_csr__reset_mstatus_WIRE_tw =1'h0; 
    wire core_csr__reset_mstatus_WIRE_tvm =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mxr =1'h0; 
    wire core_csr__reset_mstatus_WIRE_sum =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mprv =1'h0; 
    wire core_csr__reset_mstatus_WIRE_spp =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mpie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_ube =1'h0; 
    wire core_csr__reset_mstatus_WIRE_spie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_upie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_mie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_hie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_sie =1'h0; 
    wire core_csr__reset_mstatus_WIRE_uie =1'h0; 
    wire core_csr__reset_dcsr_WIRE_ebreakm =1'h0; 
    wire core_csr__reset_dcsr_WIRE_ebreakh =1'h0; 
    wire core_csr__reset_dcsr_WIRE_ebreaks =1'h0; 
    wire core_csr__reset_dcsr_WIRE_ebreaku =1'h0; 
    wire core_csr__reset_dcsr_WIRE_zero2 =1'h0; 
    wire core_csr__reset_dcsr_WIRE_stopcycle =1'h0; 
    wire core_csr__reset_dcsr_WIRE_stoptime =1'h0; 
    wire core_csr__reset_dcsr_WIRE_v =1'h0; 
    wire core_csr__reset_dcsr_WIRE_step =1'h0; 
    wire core_csr_sup_zero1 =1'h0; 
    wire core_csr_sup_debug =1'h0; 
    wire core_csr_sup_rocc =1'h0; 
    wire core_csr_sup_sgeip =1'h0; 
    wire core_csr_sup_vseip =1'h0; 
    wire core_csr_sup_seip =1'h0; 
    wire core_csr_sup_ueip =1'h0; 
    wire core_csr_sup_vstip =1'h0; 
    wire core_csr_sup_stip =1'h0; 
    wire core_csr_sup_utip =1'h0; 
    wire core_csr_sup_vssip =1'h0; 
    wire core_csr_sup_ssip =1'h0; 
    wire core_csr_sup_usip =1'h0; 
    wire core_csr_del_meip =1'h0; 
    wire core_csr_del_mtip =1'h0; 
    wire core_csr_del_msip =1'h0; 
    wire core_csr__always_WIRE_zero1 =1'h0; 
    wire core_csr__always_WIRE_debug =1'h0; 
    wire core_csr__always_WIRE_rocc =1'h0; 
    wire core_csr__always_WIRE_sgeip =1'h0; 
    wire core_csr__always_WIRE_meip =1'h0; 
    wire core_csr__always_WIRE_vseip =1'h0; 
    wire core_csr__always_WIRE_seip =1'h0; 
    wire core_csr__always_WIRE_ueip =1'h0; 
    wire core_csr__always_WIRE_mtip =1'h0; 
    wire core_csr__always_WIRE_vstip =1'h0; 
    wire core_csr__always_WIRE_stip =1'h0; 
    wire core_csr__always_WIRE_utip =1'h0; 
    wire core_csr__always_WIRE_msip =1'h0; 
    wire core_csr__always_WIRE_vssip =1'h0; 
    wire core_csr__always_WIRE_ssip =1'h0; 
    wire core_csr__always_WIRE_usip =1'h0; 
    wire core_csr_always_vseip =1'h0; 
    wire core_csr_always_vstip =1'h0; 
    wire core_csr_always_vssip =1'h0; 
    wire core_csr__reset_mnstatus_WIRE_mpv =1'h0; 
    wire core_csr__reset_mnstatus_WIRE_mie =1'h0; 
    wire core_csr__reg_menvcfg_WIRE_stce =1'h0; 
    wire core_csr__reg_menvcfg_WIRE_pbmte =1'h0; 
    wire core_csr__reg_menvcfg_WIRE_cbze =1'h0; 
    wire core_csr__reg_menvcfg_WIRE_cbcfe =1'h0; 
    wire core_csr__reg_menvcfg_WIRE_fiom =1'h0; 
    wire core_csr__reg_senvcfg_WIRE_stce =1'h0; 
    wire core_csr__reg_senvcfg_WIRE_pbmte =1'h0; 
    wire core_csr__reg_senvcfg_WIRE_cbze =1'h0; 
    wire core_csr__reg_senvcfg_WIRE_cbcfe =1'h0; 
    wire core_csr__reg_senvcfg_WIRE_fiom =1'h0; 
    wire core_csr__reg_henvcfg_WIRE_stce =1'h0; 
    wire core_csr__reg_henvcfg_WIRE_pbmte =1'h0; 
    wire core_csr__reg_henvcfg_WIRE_cbze =1'h0; 
    wire core_csr__reg_henvcfg_WIRE_cbcfe =1'h0; 
    wire core_csr__reg_henvcfg_WIRE_fiom =1'h0; 
    wire core_csr__reg_hstatus_WIRE_vtsr =1'h0; 
    wire core_csr__reg_hstatus_WIRE_vtw =1'h0; 
    wire core_csr__reg_hstatus_WIRE_vtvm =1'h0; 
    wire core_csr__reg_hstatus_WIRE_hu =1'h0; 
    wire core_csr__reg_hstatus_WIRE_spvp =1'h0; 
    wire core_csr__reg_hstatus_WIRE_spv =1'h0; 
    wire core_csr__reg_hstatus_WIRE_gva =1'h0; 
    wire core_csr__reg_hstatus_WIRE_vsbe =1'h0; 
    wire core_csr__read_mnstatus_WIRE_mpv =1'h0; 
    wire core_csr__read_mnstatus_WIRE_mie =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_zero1 =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_debug =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_rocc =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_sgeip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_meip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_vseip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_seip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_ueip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_mtip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_vstip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_stip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_utip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_msip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_vssip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_ssip =1'h0; 
    wire core_csr__sie_mask_sgeip_mask_WIRE_usip =1'h0; 
    wire core_csr_read_pmp_15_cfg_l =1'h0; 
    wire core_csr_read_pmp_15_cfg_x =1'h0; 
    wire core_csr_read_pmp_15_cfg_w =1'h0; 
    wire core_csr_read_pmp_15_cfg_r =1'h0; 
    wire core_csr_io_decode_0_fp_csr_plaOutput =1'h0; 
    wire core_csr_io_decode_0_read_illegal_plaOutput_1 =1'h0; 
    wire core_csr_delegate =1'h0; 
    wire core_csr_trapToNmiInt =1'h0; 
    wire core_csr_trapToNmiXcpt =1'h0; 
    wire core_csr_delegable_17 =1'h0; 
    wire core_csr_delegable_21 =1'h0; 
    wire core_csr_delegable_23 =1'h0; 
    wire core_csr_delegable_24 =1'h0; 
    wire[63:0] core_csr__io_rw_rdata_WIRE ; 
    wire core_csr_set_vs_dirty =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_dmode =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_action =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_chain =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_m =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_h =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_s =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_u =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_x =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_w =1'h0; 
    wire core_csr__reg_bp_1_WIRE_control_r =1'h0; 
    wire core_csr__reg_bp_1_WIRE_textra_mselect =1'h0; 
    wire core_csr__reg_bp_1_WIRE_textra_pad1 =1'h0; 
    wire core_csr__reg_bp_1_WIRE_textra_sselect =1'h0; 
    wire core_csr_reset_mstatus_debug = core_csr__reset_mstatus_WIRE_debug ; 
    wire core_csr_reset_mstatus_cease = core_csr__reset_mstatus_WIRE_cease ; 
    wire core_csr_reset_mstatus_wfi = core_csr__reset_mstatus_WIRE_wfi ; 
    wire[31:0] core_csr_reset_mstatus_isa = core_csr__reset_mstatus_WIRE_isa ; 
    wire[1:0] core_csr_reset_mstatus_dprv = core_csr__reset_mstatus_WIRE_dprv ; 
    wire core_csr_reset_mstatus_dv = core_csr__reset_mstatus_WIRE_dv ; 
    wire core_csr_reset_mstatus_v = core_csr__reset_mstatus_WIRE_v ; 
    wire core_csr_reset_mstatus_sd = core_csr__reset_mstatus_WIRE_sd ; 
    wire[22:0] core_csr_reset_mstatus_zero2 = core_csr__reset_mstatus_WIRE_zero2 ; 
    wire core_csr_reset_mstatus_mpv = core_csr__reset_mstatus_WIRE_mpv ; 
    wire core_csr_reset_mstatus_gva = core_csr__reset_mstatus_WIRE_gva ; 
    wire core_csr_reset_mstatus_mbe = core_csr__reset_mstatus_WIRE_mbe ; 
    wire core_csr_reset_mstatus_sbe = core_csr__reset_mstatus_WIRE_sbe ; 
    wire[1:0] core_csr_reset_mstatus_sxl = core_csr__reset_mstatus_WIRE_sxl ; 
    wire[1:0] core_csr_reset_mstatus_uxl = core_csr__reset_mstatus_WIRE_uxl ; 
    wire core_csr_reset_mstatus_sd_rv32 = core_csr__reset_mstatus_WIRE_sd_rv32 ; 
    wire[7:0] core_csr_reset_mstatus_zero1 = core_csr__reset_mstatus_WIRE_zero1 ; 
    wire core_csr_reset_mstatus_tsr = core_csr__reset_mstatus_WIRE_tsr ; 
    wire core_csr_reset_mstatus_tw = core_csr__reset_mstatus_WIRE_tw ; 
    wire core_csr_reset_mstatus_tvm = core_csr__reset_mstatus_WIRE_tvm ; 
    wire core_csr_reset_mstatus_mxr = core_csr__reset_mstatus_WIRE_mxr ; 
    wire core_csr_reset_mstatus_sum = core_csr__reset_mstatus_WIRE_sum ; 
    wire core_csr_reset_mstatus_mprv = core_csr__reset_mstatus_WIRE_mprv ; 
    wire[1:0] core_csr_reset_mstatus_fs = core_csr__reset_mstatus_WIRE_fs ; 
    wire[1:0] core_csr_reset_mstatus_vs = core_csr__reset_mstatus_WIRE_vs ; 
    wire core_csr_reset_mstatus_spp = core_csr__reset_mstatus_WIRE_spp ; 
    wire core_csr_reset_mstatus_mpie = core_csr__reset_mstatus_WIRE_mpie ; 
    wire core_csr_reset_mstatus_ube = core_csr__reset_mstatus_WIRE_ube ; 
    wire core_csr_reset_mstatus_spie = core_csr__reset_mstatus_WIRE_spie ; 
    wire core_csr_reset_mstatus_upie = core_csr__reset_mstatus_WIRE_upie ; 
    wire core_csr_reset_mstatus_mie = core_csr__reset_mstatus_WIRE_mie ; 
    wire core_csr_reset_mstatus_hie = core_csr__reset_mstatus_WIRE_hie ; 
    wire core_csr_reset_mstatus_sie = core_csr__reset_mstatus_WIRE_sie ; 
    wire core_csr_reset_mstatus_uie = core_csr__reset_mstatus_WIRE_uie ; 
    wire[1:0] core_csr_reset_mstatus_xs =2'h0; 
    reg core_csr_reg_mstatus_debug ; 
    reg core_csr_reg_mstatus_cease ; 
    reg core_csr_reg_mstatus_wfi ; reg[31:0] core_csr_reg_mstatus_isa ; reg[1:0] core_csr_reg_mstatus_dprv ; 
    reg core_csr_reg_mstatus_dv ; reg[1:0] core_csr_reg_mstatus_prv ; 
    wire[1:0] core_csr__io_status_prv_output = core_csr_reg_mstatus_prv ; 
    reg core_csr_reg_mstatus_v ; 
    wire core_csr__io_status_v_output = core_csr_reg_mstatus_v ; 
    reg core_csr_reg_mstatus_sd ; reg[22:0] core_csr_reg_mstatus_zero2 ; 
    wire[22:0] core_csr__io_status_zero2_output = core_csr_reg_mstatus_zero2 ; 
    reg core_csr_reg_mstatus_mpv ; 
    wire core_csr__io_status_mpv_output = core_csr_reg_mstatus_mpv ; 
    reg core_csr_reg_mstatus_gva ; 
    wire core_csr__io_status_gva_output = core_csr_reg_mstatus_gva ; 
    reg core_csr_reg_mstatus_mbe ; 
    wire core_csr__io_status_mbe_output = core_csr_reg_mstatus_mbe ; 
    reg core_csr_reg_mstatus_sbe ; 
    wire core_csr__io_status_sbe_output = core_csr_reg_mstatus_sbe ; reg[1:0] core_csr_reg_mstatus_sxl ; reg[1:0] core_csr_reg_mstatus_uxl ; 
    reg core_csr_reg_mstatus_sd_rv32 ; reg[7:0] core_csr_reg_mstatus_zero1 ; 
    wire[7:0] core_csr__io_status_zero1_output = core_csr_reg_mstatus_zero1 ; 
    reg core_csr_reg_mstatus_tsr ; 
    wire core_csr__io_status_tsr_output = core_csr_reg_mstatus_tsr ; 
    reg core_csr_reg_mstatus_tw ; 
    wire core_csr__io_status_tw_output = core_csr_reg_mstatus_tw ; 
    reg core_csr_reg_mstatus_tvm ; 
    wire core_csr__io_status_tvm_output = core_csr_reg_mstatus_tvm ; 
    reg core_csr_reg_mstatus_mxr ; 
    wire core_csr__io_status_mxr_output = core_csr_reg_mstatus_mxr ; 
    reg core_csr_reg_mstatus_sum ; 
    wire core_csr__io_status_sum_output = core_csr_reg_mstatus_sum ; 
    reg core_csr_reg_mstatus_mprv ; 
    wire core_csr__io_status_mprv_output = core_csr_reg_mstatus_mprv ; reg[1:0] core_csr_reg_mstatus_xs ; 
    wire[1:0] core_csr__io_status_xs_output = core_csr_reg_mstatus_xs ; reg[1:0] core_csr_reg_mstatus_fs ; 
    wire[1:0] core_csr__io_status_fs_output = core_csr_reg_mstatus_fs ; reg[1:0] core_csr_reg_mstatus_mpp ; 
    wire[1:0] core_csr__io_status_mpp_output = core_csr_reg_mstatus_mpp ; reg[1:0] core_csr_reg_mstatus_vs ; 
    wire[1:0] core_csr__io_status_vs_output = core_csr_reg_mstatus_vs ; 
    reg core_csr_reg_mstatus_spp ; 
    wire core_csr__io_status_spp_output = core_csr_reg_mstatus_spp ; 
    reg core_csr_reg_mstatus_mpie ; 
    wire core_csr__io_status_mpie_output = core_csr_reg_mstatus_mpie ; 
    reg core_csr_reg_mstatus_ube ; 
    wire core_csr__io_status_ube_output = core_csr_reg_mstatus_ube ; 
    reg core_csr_reg_mstatus_spie ; 
    wire core_csr__io_status_spie_output = core_csr_reg_mstatus_spie ; 
    reg core_csr_reg_mstatus_upie ; 
    wire core_csr__io_status_upie_output = core_csr_reg_mstatus_upie ; 
    reg core_csr_reg_mstatus_mie ; 
    wire core_csr__io_status_mie_output = core_csr_reg_mstatus_mie ; 
    reg core_csr_reg_mstatus_hie ; 
    wire core_csr__io_status_hie_output = core_csr_reg_mstatus_hie ; 
    reg core_csr_reg_mstatus_sie ; 
    wire core_csr__io_status_sie_output = core_csr_reg_mstatus_sie ; 
    reg core_csr_reg_mstatus_uie ; 
    wire core_csr__io_status_uie_output = core_csr_reg_mstatus_uie ; 
    wire[1:0] core_csr_reset_dcsr_zero4 = core_csr__reset_dcsr_WIRE_zero4 ; 
    wire[11:0] core_csr_reset_dcsr_zero3 = core_csr__reset_dcsr_WIRE_zero3 ; 
    wire core_csr_reset_dcsr_ebreakm = core_csr__reset_dcsr_WIRE_ebreakm ; 
    wire core_csr_reset_dcsr_ebreakh = core_csr__reset_dcsr_WIRE_ebreakh ; 
    wire core_csr_reset_dcsr_ebreaks = core_csr__reset_dcsr_WIRE_ebreaks ; 
    wire core_csr_reset_dcsr_ebreaku = core_csr__reset_dcsr_WIRE_ebreaku ; 
    wire core_csr_reset_dcsr_zero2 = core_csr__reset_dcsr_WIRE_zero2 ; 
    wire core_csr_reset_dcsr_stopcycle = core_csr__reset_dcsr_WIRE_stopcycle ; 
    wire core_csr_reset_dcsr_stoptime = core_csr__reset_dcsr_WIRE_stoptime ; 
    wire[2:0] core_csr_reset_dcsr_cause = core_csr__reset_dcsr_WIRE_cause ; 
    wire core_csr_reset_dcsr_v = core_csr__reset_dcsr_WIRE_v ; 
    wire[1:0] core_csr_reset_dcsr_zero1 = core_csr__reset_dcsr_WIRE_zero1 ; 
    wire core_csr_reset_dcsr_step = core_csr__reset_dcsr_WIRE_step ; 
    wire[1:0] core_csr_reset_dcsr_xdebugver =2'h1; reg[1:0] core_csr_reg_dcsr_xdebugver ; reg[1:0] core_csr_reg_dcsr_zero4 ; reg[11:0] core_csr_reg_dcsr_zero3 ; 
    reg core_csr_reg_dcsr_ebreakm ; 
    reg core_csr_reg_dcsr_ebreakh ; 
    reg core_csr_reg_dcsr_ebreaks ; 
    reg core_csr_reg_dcsr_ebreaku ; 
    reg core_csr_reg_dcsr_zero2 ; 
    reg core_csr_reg_dcsr_stopcycle ; 
    reg core_csr_reg_dcsr_stoptime ; reg[2:0] core_csr_reg_dcsr_cause ; 
    reg core_csr_reg_dcsr_v ; reg[1:0] core_csr_reg_dcsr_zero1 ; 
    reg core_csr_reg_dcsr_step ; reg[1:0] core_csr_reg_dcsr_prv ; 
    wire core_csr_del_zero1 = core_csr_sup_zero1 ; 
    wire core_csr_del_debug = core_csr_sup_debug ; 
    wire core_csr_del_rocc = core_csr_sup_rocc ; 
    wire core_csr_del_sgeip = core_csr_sup_sgeip ; 
    wire core_csr_del_vseip = core_csr_sup_vseip ; 
    wire core_csr_del_seip = core_csr_sup_seip ; 
    wire core_csr_del_ueip = core_csr_sup_ueip ; 
    wire core_csr_del_vstip = core_csr_sup_vstip ; 
    wire core_csr_del_stip = core_csr_sup_stip ; 
    wire core_csr_del_utip = core_csr_sup_utip ; 
    wire core_csr_del_vssip = core_csr_sup_vssip ; 
    wire core_csr_del_ssip = core_csr_sup_ssip ; 
    wire core_csr_del_usip = core_csr_sup_usip ; 
    wire[1:0] core_csr_lo_lo_lo ={ core_csr_sup_ssip , core_csr_sup_usip }; 
    wire[1:0] core_csr_lo_lo_hi ={ core_csr_sup_msip , core_csr_sup_vssip }; 
    wire[3:0] core_csr_lo_lo ={ core_csr_lo_lo_hi , core_csr_lo_lo_lo }; 
    wire[1:0] core_csr_lo_hi_lo ={ core_csr_sup_stip , core_csr_sup_utip }; 
    wire[1:0] core_csr_lo_hi_hi ={ core_csr_sup_mtip , core_csr_sup_vstip }; 
    wire[3:0] core_csr_lo_hi ={ core_csr_lo_hi_hi , core_csr_lo_hi_lo }; 
    wire[7:0] core_csr_lo ={ core_csr_lo_hi , core_csr_lo_lo }; 
    wire[1:0] core_csr_hi_lo_lo ={ core_csr_sup_seip , core_csr_sup_ueip }; 
    wire[1:0] core_csr_hi_lo_hi ={ core_csr_sup_meip , core_csr_sup_vseip }; 
    wire[3:0] core_csr_hi_lo ={ core_csr_hi_lo_hi , core_csr_hi_lo_lo }; 
    wire[1:0] core_csr_hi_hi_lo ={ core_csr_sup_rocc , core_csr_sup_sgeip }; 
    wire[1:0] core_csr_hi_hi_hi ={ core_csr_sup_zero1 , core_csr_sup_debug }; 
    wire[3:0] core_csr_hi_hi ={ core_csr_hi_hi_hi , core_csr_hi_hi_lo }; 
    wire[7:0] core_csr_hi ={ core_csr_hi_hi , core_csr_hi_lo }; 
    wire[15:0] core_csr_supported_interrupts ={ core_csr_hi , core_csr_lo }; 
    wire[1:0] core_csr_lo_lo_lo_1 ={ core_csr_del_ssip , core_csr_del_usip }; 
    wire[1:0] core_csr_lo_lo_hi_1 ={ core_csr_del_msip , core_csr_del_vssip }; 
    wire[3:0] core_csr_lo_lo_1 ={ core_csr_lo_lo_hi_1 , core_csr_lo_lo_lo_1 }; 
    wire[1:0] core_csr_lo_hi_lo_1 ={ core_csr_del_stip , core_csr_del_utip }; 
    wire[1:0] core_csr_lo_hi_hi_1 ={ core_csr_del_mtip , core_csr_del_vstip }; 
    wire[3:0] core_csr_lo_hi_1 ={ core_csr_lo_hi_hi_1 , core_csr_lo_hi_lo_1 }; 
    wire[7:0] core_csr_lo_1 ={ core_csr_lo_hi_1 , core_csr_lo_lo_1 }; 
    wire[1:0] core_csr_hi_lo_lo_1 ={ core_csr_del_seip , core_csr_del_ueip }; 
    wire[1:0] core_csr_hi_lo_hi_1 ={ core_csr_del_meip , core_csr_del_vseip }; 
    wire[3:0] core_csr_hi_lo_1 ={ core_csr_hi_lo_hi_1 , core_csr_hi_lo_lo_1 }; 
    wire[1:0] core_csr_hi_hi_lo_1 ={ core_csr_del_rocc , core_csr_del_sgeip }; 
    wire[1:0] core_csr_hi_hi_hi_1 ={ core_csr_del_zero1 , core_csr_del_debug }; 
    wire[3:0] core_csr_hi_hi_1 ={ core_csr_hi_hi_hi_1 , core_csr_hi_hi_lo_1 }; 
    wire[7:0] core_csr_hi_1 ={ core_csr_hi_hi_1 , core_csr_hi_lo_1 }; 
    wire[15:0] core_csr_delegable_interrupts ={ core_csr_hi_1 , core_csr_lo_1 }; 
    wire core_csr_always_zero1 = core_csr__always_WIRE_zero1 ; 
    wire core_csr_always_debug = core_csr__always_WIRE_debug ; 
    wire core_csr_always_rocc = core_csr__always_WIRE_rocc ; 
    wire core_csr_always_sgeip = core_csr__always_WIRE_sgeip ; 
    wire core_csr_always_meip = core_csr__always_WIRE_meip ; 
    wire core_csr_always_seip = core_csr__always_WIRE_seip ; 
    wire core_csr_always_ueip = core_csr__always_WIRE_ueip ; 
    wire core_csr_always_mtip = core_csr__always_WIRE_mtip ; 
    wire core_csr_always_stip = core_csr__always_WIRE_stip ; 
    wire core_csr_always_utip = core_csr__always_WIRE_utip ; 
    wire core_csr_always_msip = core_csr__always_WIRE_msip ; 
    wire core_csr_always_ssip = core_csr__always_WIRE_ssip ; 
    wire core_csr_always_usip = core_csr__always_WIRE_usip ; 
    wire core_csr_deleg_zero1 = core_csr_always_zero1 ; 
    wire core_csr_deleg_debug = core_csr_always_debug ; 
    wire core_csr_deleg_rocc = core_csr_always_rocc ; 
    wire core_csr_deleg_sgeip = core_csr_always_sgeip ; 
    wire core_csr_deleg_meip = core_csr_always_meip ; 
    wire core_csr_deleg_vseip = core_csr_always_vseip ; 
    wire core_csr_deleg_seip = core_csr_always_seip ; 
    wire core_csr_deleg_ueip = core_csr_always_ueip ; 
    wire core_csr_deleg_mtip = core_csr_always_mtip ; 
    wire core_csr_deleg_vstip = core_csr_always_vstip ; 
    wire core_csr_deleg_stip = core_csr_always_stip ; 
    wire core_csr_deleg_utip = core_csr_always_utip ; 
    wire core_csr_deleg_msip = core_csr_always_msip ; 
    wire core_csr_deleg_vssip = core_csr_always_vssip ; 
    wire core_csr_deleg_ssip = core_csr_always_ssip ; 
    wire core_csr_deleg_usip = core_csr_always_usip ; 
    wire[1:0] core_csr_lo_lo_lo_2 ={ core_csr_deleg_ssip , core_csr_deleg_usip }; 
    wire[1:0] core_csr_lo_lo_hi_2 ={ core_csr_deleg_msip , core_csr_deleg_vssip }; 
    wire[3:0] core_csr_lo_lo_2 ={ core_csr_lo_lo_hi_2 , core_csr_lo_lo_lo_2 }; 
    wire[1:0] core_csr_lo_hi_lo_2 ={ core_csr_deleg_stip , core_csr_deleg_utip }; 
    wire[1:0] core_csr_lo_hi_hi_2 ={ core_csr_deleg_mtip , core_csr_deleg_vstip }; 
    wire[3:0] core_csr_lo_hi_2 ={ core_csr_lo_hi_hi_2 , core_csr_lo_hi_lo_2 }; 
    wire[7:0] core_csr_lo_2 ={ core_csr_lo_hi_2 , core_csr_lo_lo_2 }; 
    wire[1:0] core_csr_hi_lo_lo_2 ={ core_csr_deleg_seip , core_csr_deleg_ueip }; 
    wire[1:0] core_csr_hi_lo_hi_2 ={ core_csr_deleg_meip , core_csr_deleg_vseip }; 
    wire[3:0] core_csr_hi_lo_2 ={ core_csr_hi_lo_hi_2 , core_csr_hi_lo_lo_2 }; 
    wire[1:0] core_csr_hi_hi_lo_2 ={ core_csr_deleg_rocc , core_csr_deleg_sgeip }; 
    wire[1:0] core_csr_hi_hi_hi_2 ={ core_csr_deleg_zero1 , core_csr_deleg_debug }; 
    wire[3:0] core_csr_hi_hi_2 ={ core_csr_hi_hi_hi_2 , core_csr_hi_hi_lo_2 }; 
    wire[7:0] core_csr_hi_2 ={ core_csr_hi_hi_2 , core_csr_hi_lo_2 }; 
    wire[15:0] core_csr_hs_delegable_interrupts ={ core_csr_hi_2 , core_csr_lo_2 }; 
    wire[1:0] core_csr_lo_lo_lo_3 ={ core_csr_always_ssip , core_csr_always_usip }; 
    wire[1:0] core_csr_lo_lo_hi_3 ={ core_csr_always_msip , core_csr_always_vssip }; 
    wire[3:0] core_csr_lo_lo_3 ={ core_csr_lo_lo_hi_3 , core_csr_lo_lo_lo_3 }; 
    wire[1:0] core_csr_lo_hi_lo_3 ={ core_csr_always_stip , core_csr_always_utip }; 
    wire[1:0] core_csr_lo_hi_hi_3 ={ core_csr_always_mtip , core_csr_always_vstip }; 
    wire[3:0] core_csr_lo_hi_3 ={ core_csr_lo_hi_hi_3 , core_csr_lo_hi_lo_3 }; 
    wire[7:0] core_csr_lo_3 ={ core_csr_lo_hi_3 , core_csr_lo_lo_3 }; 
    wire[1:0] core_csr_hi_lo_lo_3 ={ core_csr_always_seip , core_csr_always_ueip }; 
    wire[1:0] core_csr_hi_lo_hi_3 ={ core_csr_always_meip , core_csr_always_vseip }; 
    wire[3:0] core_csr_hi_lo_3 ={ core_csr_hi_lo_hi_3 , core_csr_hi_lo_lo_3 }; 
    wire[1:0] core_csr_hi_hi_lo_3 ={ core_csr_always_rocc , core_csr_always_sgeip }; 
    wire[1:0] core_csr_hi_hi_hi_3 ={ core_csr_always_zero1 , core_csr_always_debug }; 
    wire[3:0] core_csr_hi_hi_3 ={ core_csr_hi_hi_hi_3 , core_csr_hi_hi_lo_3 }; 
    wire[7:0] core_csr_hi_3 ={ core_csr_hi_hi_3 , core_csr_hi_lo_3 }; 
    wire[15:0] core_csr_mideleg_always_hs ={ core_csr_hi_3 , core_csr_lo_3 }; 
    reg core_csr_reg_debug ; 
    wire core_csr__io_status_debug_output = core_csr_reg_debug ; reg[33:0] core_csr_reg_dpc ; reg[63:0] core_csr_reg_dscratch0 ; 
    reg core_csr_reg_singleStepped ; 
    reg core_csr_reg_tselect ; reg[3:0] core_csr_reg_bp_0_control_ttype ; 
    reg core_csr_reg_bp_0_control_dmode ; reg[5:0] core_csr_reg_bp_0_control_maskmax ; reg[39:0] core_csr_reg_bp_0_control_reserved ; 
    reg core_csr_reg_bp_0_control_action ; 
    reg core_csr_reg_bp_0_control_chain ; reg[1:0] core_csr_reg_bp_0_control_zero ; reg[1:0] core_csr_reg_bp_0_control_tmatch ; 
    reg core_csr_reg_bp_0_control_m ; 
    reg core_csr_reg_bp_0_control_h ; 
    reg core_csr_reg_bp_0_control_s ; 
    reg core_csr_reg_bp_0_control_u ; 
    reg core_csr_reg_bp_0_control_x ; 
    reg core_csr_reg_bp_0_control_w ; 
    reg core_csr_reg_bp_0_control_r ; reg[32:0] core_csr_reg_bp_0_address ; 
    reg core_csr_reg_bp_0_textra_mselect ; reg[47:0] core_csr_reg_bp_0_textra_pad2 ; 
    reg core_csr_reg_bp_0_textra_pad1 ; 
    reg core_csr_reg_bp_0_textra_sselect ; reg[3:0] core_csr_reg_bp_1_control_ttype ; 
    reg core_csr_reg_bp_1_control_dmode ; reg[5:0] core_csr_reg_bp_1_control_maskmax ; reg[39:0] core_csr_reg_bp_1_control_reserved ; 
    reg core_csr_reg_bp_1_control_action ; 
    reg core_csr_reg_bp_1_control_chain ; reg[1:0] core_csr_reg_bp_1_control_zero ; reg[1:0] core_csr_reg_bp_1_control_tmatch ; 
    reg core_csr_reg_bp_1_control_m ; 
    reg core_csr_reg_bp_1_control_h ; 
    reg core_csr_reg_bp_1_control_s ; 
    reg core_csr_reg_bp_1_control_u ; 
    reg core_csr_reg_bp_1_control_x ; 
    reg core_csr_reg_bp_1_control_w ; 
    reg core_csr_reg_bp_1_control_r ; reg[32:0] core_csr_reg_bp_1_address ; 
    reg core_csr_reg_bp_1_textra_mselect ; reg[47:0] core_csr_reg_bp_1_textra_pad2 ; 
    reg core_csr_reg_bp_1_textra_pad1 ; 
    reg core_csr_reg_bp_1_textra_sselect ; 
    reg core_csr_reg_pmp_0_cfg_l ; 
    wire core_csr_pmp_cfg_l = core_csr_reg_pmp_0_cfg_l ; reg[1:0] core_csr_reg_pmp_0_cfg_res ; 
    wire[1:0] core_csr_pmp_cfg_res = core_csr_reg_pmp_0_cfg_res ; reg[1:0] core_csr_reg_pmp_0_cfg_a ; 
    wire[1:0] core_csr_pmp_cfg_a = core_csr_reg_pmp_0_cfg_a ; 
    reg core_csr_reg_pmp_0_cfg_x ; 
    wire core_csr_pmp_cfg_x = core_csr_reg_pmp_0_cfg_x ; 
    reg core_csr_reg_pmp_0_cfg_w ; 
    wire core_csr_pmp_cfg_w = core_csr_reg_pmp_0_cfg_w ; 
    reg core_csr_reg_pmp_0_cfg_r ; 
    wire core_csr_pmp_cfg_r = core_csr_reg_pmp_0_cfg_r ; reg[29:0] core_csr_reg_pmp_0_addr ; 
    wire[29:0] core_csr_pmp_addr = core_csr_reg_pmp_0_addr ; 
    reg core_csr_reg_pmp_1_cfg_l ; 
    wire core_csr_pmp_1_cfg_l = core_csr_reg_pmp_1_cfg_l ; reg[1:0] core_csr_reg_pmp_1_cfg_res ; 
    wire[1:0] core_csr_pmp_1_cfg_res = core_csr_reg_pmp_1_cfg_res ; reg[1:0] core_csr_reg_pmp_1_cfg_a ; 
    wire[1:0] core_csr_pmp_1_cfg_a = core_csr_reg_pmp_1_cfg_a ; 
    reg core_csr_reg_pmp_1_cfg_x ; 
    wire core_csr_pmp_1_cfg_x = core_csr_reg_pmp_1_cfg_x ; 
    reg core_csr_reg_pmp_1_cfg_w ; 
    wire core_csr_pmp_1_cfg_w = core_csr_reg_pmp_1_cfg_w ; 
    reg core_csr_reg_pmp_1_cfg_r ; 
    wire core_csr_pmp_1_cfg_r = core_csr_reg_pmp_1_cfg_r ; reg[29:0] core_csr_reg_pmp_1_addr ; 
    wire[29:0] core_csr_pmp_1_addr = core_csr_reg_pmp_1_addr ; 
    reg core_csr_reg_pmp_2_cfg_l ; 
    wire core_csr_pmp_2_cfg_l = core_csr_reg_pmp_2_cfg_l ; reg[1:0] core_csr_reg_pmp_2_cfg_res ; 
    wire[1:0] core_csr_pmp_2_cfg_res = core_csr_reg_pmp_2_cfg_res ; reg[1:0] core_csr_reg_pmp_2_cfg_a ; 
    wire[1:0] core_csr_pmp_2_cfg_a = core_csr_reg_pmp_2_cfg_a ; 
    reg core_csr_reg_pmp_2_cfg_x ; 
    wire core_csr_pmp_2_cfg_x = core_csr_reg_pmp_2_cfg_x ; 
    reg core_csr_reg_pmp_2_cfg_w ; 
    wire core_csr_pmp_2_cfg_w = core_csr_reg_pmp_2_cfg_w ; 
    reg core_csr_reg_pmp_2_cfg_r ; 
    wire core_csr_pmp_2_cfg_r = core_csr_reg_pmp_2_cfg_r ; reg[29:0] core_csr_reg_pmp_2_addr ; 
    wire[29:0] core_csr_pmp_2_addr = core_csr_reg_pmp_2_addr ; 
    reg core_csr_reg_pmp_3_cfg_l ; 
    wire core_csr_pmp_3_cfg_l = core_csr_reg_pmp_3_cfg_l ; reg[1:0] core_csr_reg_pmp_3_cfg_res ; 
    wire[1:0] core_csr_pmp_3_cfg_res = core_csr_reg_pmp_3_cfg_res ; reg[1:0] core_csr_reg_pmp_3_cfg_a ; 
    wire[1:0] core_csr_pmp_3_cfg_a = core_csr_reg_pmp_3_cfg_a ; 
    reg core_csr_reg_pmp_3_cfg_x ; 
    wire core_csr_pmp_3_cfg_x = core_csr_reg_pmp_3_cfg_x ; 
    reg core_csr_reg_pmp_3_cfg_w ; 
    wire core_csr_pmp_3_cfg_w = core_csr_reg_pmp_3_cfg_w ; 
    reg core_csr_reg_pmp_3_cfg_r ; 
    wire core_csr_pmp_3_cfg_r = core_csr_reg_pmp_3_cfg_r ; reg[29:0] core_csr_reg_pmp_3_addr ; 
    wire[29:0] core_csr_pmp_3_addr = core_csr_reg_pmp_3_addr ; 
    reg core_csr_reg_pmp_4_cfg_l ; 
    wire core_csr_pmp_4_cfg_l = core_csr_reg_pmp_4_cfg_l ; reg[1:0] core_csr_reg_pmp_4_cfg_res ; 
    wire[1:0] core_csr_pmp_4_cfg_res = core_csr_reg_pmp_4_cfg_res ; reg[1:0] core_csr_reg_pmp_4_cfg_a ; 
    wire[1:0] core_csr_pmp_4_cfg_a = core_csr_reg_pmp_4_cfg_a ; 
    reg core_csr_reg_pmp_4_cfg_x ; 
    wire core_csr_pmp_4_cfg_x = core_csr_reg_pmp_4_cfg_x ; 
    reg core_csr_reg_pmp_4_cfg_w ; 
    wire core_csr_pmp_4_cfg_w = core_csr_reg_pmp_4_cfg_w ; 
    reg core_csr_reg_pmp_4_cfg_r ; 
    wire core_csr_pmp_4_cfg_r = core_csr_reg_pmp_4_cfg_r ; reg[29:0] core_csr_reg_pmp_4_addr ; 
    wire[29:0] core_csr_pmp_4_addr = core_csr_reg_pmp_4_addr ; 
    reg core_csr_reg_pmp_5_cfg_l ; 
    wire core_csr_pmp_5_cfg_l = core_csr_reg_pmp_5_cfg_l ; reg[1:0] core_csr_reg_pmp_5_cfg_res ; 
    wire[1:0] core_csr_pmp_5_cfg_res = core_csr_reg_pmp_5_cfg_res ; reg[1:0] core_csr_reg_pmp_5_cfg_a ; 
    wire[1:0] core_csr_pmp_5_cfg_a = core_csr_reg_pmp_5_cfg_a ; 
    reg core_csr_reg_pmp_5_cfg_x ; 
    wire core_csr_pmp_5_cfg_x = core_csr_reg_pmp_5_cfg_x ; 
    reg core_csr_reg_pmp_5_cfg_w ; 
    wire core_csr_pmp_5_cfg_w = core_csr_reg_pmp_5_cfg_w ; 
    reg core_csr_reg_pmp_5_cfg_r ; 
    wire core_csr_pmp_5_cfg_r = core_csr_reg_pmp_5_cfg_r ; reg[29:0] core_csr_reg_pmp_5_addr ; 
    wire[29:0] core_csr_pmp_5_addr = core_csr_reg_pmp_5_addr ; 
    reg core_csr_reg_pmp_6_cfg_l ; 
    wire core_csr_pmp_6_cfg_l = core_csr_reg_pmp_6_cfg_l ; reg[1:0] core_csr_reg_pmp_6_cfg_res ; 
    wire[1:0] core_csr_pmp_6_cfg_res = core_csr_reg_pmp_6_cfg_res ; reg[1:0] core_csr_reg_pmp_6_cfg_a ; 
    wire[1:0] core_csr_pmp_6_cfg_a = core_csr_reg_pmp_6_cfg_a ; 
    reg core_csr_reg_pmp_6_cfg_x ; 
    wire core_csr_pmp_6_cfg_x = core_csr_reg_pmp_6_cfg_x ; 
    reg core_csr_reg_pmp_6_cfg_w ; 
    wire core_csr_pmp_6_cfg_w = core_csr_reg_pmp_6_cfg_w ; 
    reg core_csr_reg_pmp_6_cfg_r ; 
    wire core_csr_pmp_6_cfg_r = core_csr_reg_pmp_6_cfg_r ; reg[29:0] core_csr_reg_pmp_6_addr ; 
    wire[29:0] core_csr_pmp_6_addr = core_csr_reg_pmp_6_addr ; 
    reg core_csr_reg_pmp_7_cfg_l ; 
    wire core_csr_pmp_7_cfg_l = core_csr_reg_pmp_7_cfg_l ; reg[1:0] core_csr_reg_pmp_7_cfg_res ; 
    wire[1:0] core_csr_pmp_7_cfg_res = core_csr_reg_pmp_7_cfg_res ; reg[1:0] core_csr_reg_pmp_7_cfg_a ; 
    wire[1:0] core_csr_pmp_7_cfg_a = core_csr_reg_pmp_7_cfg_a ; 
    reg core_csr_reg_pmp_7_cfg_x ; 
    wire core_csr_pmp_7_cfg_x = core_csr_reg_pmp_7_cfg_x ; 
    reg core_csr_reg_pmp_7_cfg_w ; 
    wire core_csr_pmp_7_cfg_w = core_csr_reg_pmp_7_cfg_w ; 
    reg core_csr_reg_pmp_7_cfg_r ; 
    wire core_csr_pmp_7_cfg_r = core_csr_reg_pmp_7_cfg_r ; reg[29:0] core_csr_reg_pmp_7_addr ; 
    wire[29:0] core_csr_pmp_7_addr = core_csr_reg_pmp_7_addr ; reg[63:0] core_csr_reg_mie ; reg[63:0] core_csr_reg_mideleg ; reg[63:0] core_csr_reg_medeleg ; 
    reg core_csr_reg_mip_zero1 ; 
    wire core_csr_mip_zero1 = core_csr_reg_mip_zero1 ; 
    reg core_csr_reg_mip_debug ; 
    wire core_csr_mip_debug = core_csr_reg_mip_debug ; 
    reg core_csr_reg_mip_rocc ; 
    reg core_csr_reg_mip_sgeip ; 
    wire core_csr_mip_sgeip = core_csr_reg_mip_sgeip ; 
    reg core_csr_reg_mip_meip ; 
    reg core_csr_reg_mip_vseip ; 
    wire core_csr_mip_vseip = core_csr_reg_mip_vseip ; 
    reg core_csr_reg_mip_seip ; 
    wire core_csr_mip_seip = core_csr_reg_mip_seip ; 
    reg core_csr_reg_mip_ueip ; 
    wire core_csr_mip_ueip = core_csr_reg_mip_ueip ; 
    reg core_csr_reg_mip_mtip ; 
    reg core_csr_reg_mip_vstip ; 
    wire core_csr_mip_vstip = core_csr_reg_mip_vstip ; 
    reg core_csr_reg_mip_stip ; 
    wire core_csr_mip_stip = core_csr_reg_mip_stip ; 
    reg core_csr_reg_mip_utip ; 
    wire core_csr_mip_utip = core_csr_reg_mip_utip ; 
    reg core_csr_reg_mip_msip ; 
    reg core_csr_reg_mip_vssip ; 
    wire core_csr_mip_vssip = core_csr_reg_mip_vssip ; 
    reg core_csr_reg_mip_ssip ; 
    wire core_csr_mip_ssip = core_csr_reg_mip_ssip ; 
    reg core_csr_reg_mip_usip ; 
    wire core_csr_mip_usip = core_csr_reg_mip_usip ; reg[33:0] core_csr_reg_mepc ; reg[63:0] core_csr_reg_mcause ; reg[33:0] core_csr_reg_mtval ; reg[39:0] core_csr_reg_mtval2 ; reg[63:0] core_csr_reg_mscratch ; reg[31:0] core_csr_reg_mtvec ; 
    wire[2:0] core_csr_reset_mnstatus_zero3 = core_csr__reset_mnstatus_WIRE_zero3 ; 
    wire core_csr_reset_mnstatus_mpv = core_csr__reset_mnstatus_WIRE_mpv ; 
    wire[2:0] core_csr_reset_mnstatus_zero2 = core_csr__reset_mnstatus_WIRE_zero2 ; 
    wire core_csr_reset_mnstatus_mie = core_csr__reset_mnstatus_WIRE_mie ; 
    wire[2:0] core_csr_reset_mnstatus_zero1 = core_csr__reset_mnstatus_WIRE_zero1 ; reg[63:0] core_csr_reg_mnscratch ; reg[33:0] core_csr_reg_mnepc ; reg[63:0] core_csr_reg_mncause ; reg[1:0] core_csr_reg_mnstatus_mpp ; 
    wire[1:0] core_csr_read_mnstatus_mpp = core_csr_reg_mnstatus_mpp ; reg[2:0] core_csr_reg_mnstatus_zero3 ; 
    reg core_csr_reg_mnstatus_mpv ; 
    wire core_csr_read_mnstatus_mpv = core_csr_reg_mnstatus_mpv ; reg[2:0] core_csr_reg_mnstatus_zero2 ; 
    reg core_csr_reg_mnstatus_mie ; reg[2:0] core_csr_reg_mnstatus_zero1 ; 
    reg core_csr_reg_rnmie ; 
    wire core_csr_read_mnstatus_mie = core_csr_reg_rnmie ; 
    reg core_csr_reg_menvcfg_stce ; 
    reg core_csr_reg_menvcfg_pbmte ; reg[53:0] core_csr_reg_menvcfg_zero54 ; 
    reg core_csr_reg_menvcfg_cbze ; 
    reg core_csr_reg_menvcfg_cbcfe ; reg[1:0] core_csr_reg_menvcfg_cbie ; reg[2:0] core_csr_reg_menvcfg_zero3 ; 
    reg core_csr_reg_menvcfg_fiom ; 
    reg core_csr_reg_senvcfg_stce ; 
    reg core_csr_reg_senvcfg_pbmte ; reg[53:0] core_csr_reg_senvcfg_zero54 ; 
    reg core_csr_reg_senvcfg_cbze ; 
    reg core_csr_reg_senvcfg_cbcfe ; reg[1:0] core_csr_reg_senvcfg_cbie ; reg[2:0] core_csr_reg_senvcfg_zero3 ; 
    reg core_csr_reg_senvcfg_fiom ; 
    reg core_csr_reg_henvcfg_stce ; 
    reg core_csr_reg_henvcfg_pbmte ; reg[53:0] core_csr_reg_henvcfg_zero54 ; 
    reg core_csr_reg_henvcfg_cbze ; 
    reg core_csr_reg_henvcfg_cbcfe ; reg[1:0] core_csr_reg_henvcfg_cbie ; reg[2:0] core_csr_reg_henvcfg_zero3 ; 
    reg core_csr_reg_henvcfg_fiom ; reg[31:0] core_csr_reg_mcounteren ; reg[31:0] core_csr_reg_scounteren ; reg[63:0] core_csr_reg_hideleg ; reg[63:0] core_csr_reg_hedeleg ; reg[31:0] core_csr_reg_hcounteren ; reg[29:0] core_csr_reg_hstatus_zero6 ; reg[1:0] core_csr_reg_hstatus_vsxl ; reg[8:0] core_csr_reg_hstatus_zero5 ; 
    reg core_csr_reg_hstatus_vtsr ; 
    reg core_csr_reg_hstatus_vtw ; 
    reg core_csr_reg_hstatus_vtvm ; reg[1:0] core_csr_reg_hstatus_zero3 ; reg[5:0] core_csr_reg_hstatus_vgein ; reg[1:0] core_csr_reg_hstatus_zero2 ; 
    reg core_csr_reg_hstatus_hu ; 
    reg core_csr_reg_hstatus_spvp ; 
    reg core_csr_reg_hstatus_spv ; 
    reg core_csr_reg_hstatus_gva ; 
    reg core_csr_reg_hstatus_vsbe ; reg[4:0] core_csr_reg_hstatus_zero1 ; reg[3:0] core_csr_reg_hgatp_mode ; reg[15:0] core_csr_reg_hgatp_asid ; reg[43:0] core_csr_reg_hgatp_ppn ; reg[39:0] core_csr_reg_htval ; 
    wire[1:0] core_csr_read_hvip_lo_lo_lo ={ core_csr_reg_mip_ssip , core_csr_reg_mip_usip }; 
    wire[1:0] core_csr_read_hvip_lo_lo_hi ={ core_csr_reg_mip_msip , core_csr_reg_mip_vssip }; 
    wire[3:0] core_csr_read_hvip_lo_lo ={ core_csr_read_hvip_lo_lo_hi , core_csr_read_hvip_lo_lo_lo }; 
    wire[1:0] core_csr_read_hvip_lo_hi_lo ={ core_csr_reg_mip_stip , core_csr_reg_mip_utip }; 
    wire[1:0] core_csr_read_hvip_lo_hi_hi ={ core_csr_reg_mip_mtip , core_csr_reg_mip_vstip }; 
    wire[3:0] core_csr_read_hvip_lo_hi ={ core_csr_read_hvip_lo_hi_hi , core_csr_read_hvip_lo_hi_lo }; 
    wire[7:0] core_csr_read_hvip_lo ={ core_csr_read_hvip_lo_hi , core_csr_read_hvip_lo_lo }; 
    wire[1:0] core_csr_read_hvip_hi_lo_lo ={ core_csr_reg_mip_seip , core_csr_reg_mip_ueip }; 
    wire[1:0] core_csr_read_hvip_hi_lo_hi ={ core_csr_reg_mip_meip , core_csr_reg_mip_vseip }; 
    wire[3:0] core_csr_read_hvip_hi_lo ={ core_csr_read_hvip_hi_lo_hi , core_csr_read_hvip_hi_lo_lo }; 
    wire[1:0] core_csr_read_hvip_hi_hi_lo ={ core_csr_reg_mip_rocc , core_csr_reg_mip_sgeip }; 
    wire[1:0] core_csr_read_hvip_hi_hi_hi ={ core_csr_reg_mip_zero1 , core_csr_reg_mip_debug }; 
    wire[3:0] core_csr_read_hvip_hi_hi ={ core_csr_read_hvip_hi_hi_hi , core_csr_read_hvip_hi_hi_lo }; 
    wire[7:0] core_csr_read_hvip_hi ={ core_csr_read_hvip_hi_hi , core_csr_read_hvip_hi_lo }; 
    wire[15:0] core_csr_read_hvip ={ core_csr_read_hvip_hi , core_csr_read_hvip_lo }& core_csr_hs_delegable_interrupts ; 
    wire[63:0] core_csr_read_hie = core_csr_reg_mie &{48'h0, core_csr_hs_delegable_interrupts }; reg[33:0] core_csr_reg_vstvec ; 
    wire[33:0] core_csr__GEN = core_csr_reg_vstvec &~{26'h0, core_csr_reg_vstvec [0] ? 8'hFE:8'h2}; 
    wire[63:0] core_csr_read_vstvec ={ core_csr__GEN [33] ? 30'h3FFFFFFF:30'h0, core_csr__GEN }; 
    reg core_csr_reg_vsstatus_debug ; 
    reg core_csr_reg_vsstatus_cease ; 
    reg core_csr_reg_vsstatus_wfi ; reg[31:0] core_csr_reg_vsstatus_isa ; reg[1:0] core_csr_reg_vsstatus_dprv ; 
    reg core_csr_reg_vsstatus_dv ; reg[1:0] core_csr_reg_vsstatus_prv ; 
    reg core_csr_reg_vsstatus_v ; 
    reg core_csr_reg_vsstatus_sd ; reg[22:0] core_csr_reg_vsstatus_zero2 ; 
    reg core_csr_reg_vsstatus_mpv ; 
    reg core_csr_reg_vsstatus_gva ; 
    reg core_csr_reg_vsstatus_mbe ; 
    reg core_csr_reg_vsstatus_sbe ; reg[1:0] core_csr_reg_vsstatus_sxl ; reg[1:0] core_csr_reg_vsstatus_uxl ; 
    reg core_csr_reg_vsstatus_sd_rv32 ; reg[7:0] core_csr_reg_vsstatus_zero1 ; 
    reg core_csr_reg_vsstatus_tsr ; 
    reg core_csr_reg_vsstatus_tw ; 
    reg core_csr_reg_vsstatus_tvm ; 
    reg core_csr_reg_vsstatus_mxr ; 
    reg core_csr_reg_vsstatus_sum ; 
    reg core_csr_reg_vsstatus_mprv ; reg[1:0] core_csr_reg_vsstatus_xs ; 
    wire[1:0] core_csr__io_gstatus_xs_output = core_csr_reg_vsstatus_xs ; reg[1:0] core_csr_reg_vsstatus_fs ; 
    wire[1:0] core_csr__io_gstatus_fs_output = core_csr_reg_vsstatus_fs ; reg[1:0] core_csr_reg_vsstatus_mpp ; reg[1:0] core_csr_reg_vsstatus_vs ; 
    wire[1:0] core_csr__io_gstatus_vs_output = core_csr_reg_vsstatus_vs ; 
    reg core_csr_reg_vsstatus_spp ; 
    reg core_csr_reg_vsstatus_mpie ; 
    reg core_csr_reg_vsstatus_ube ; 
    reg core_csr_reg_vsstatus_spie ; 
    reg core_csr_reg_vsstatus_upie ; 
    reg core_csr_reg_vsstatus_mie ; 
    reg core_csr_reg_vsstatus_hie ; 
    reg core_csr_reg_vsstatus_sie ; 
    reg core_csr_reg_vsstatus_uie ; reg[63:0] core_csr_reg_vsscratch ; reg[33:0] core_csr_reg_vsepc ; reg[63:0] core_csr_reg_vscause ; reg[33:0] core_csr_reg_vstval ; reg[3:0] core_csr_reg_vsatp_mode ; reg[15:0] core_csr_reg_vsatp_asid ; reg[43:0] core_csr_reg_vsatp_ppn ; reg[33:0] core_csr_reg_sepc ; reg[63:0] core_csr_reg_scause ; reg[33:0] core_csr_reg_stval ; reg[63:0] core_csr_reg_sscratch ; reg[32:0] core_csr_reg_stvec ; reg[3:0] core_csr_reg_satp_mode ; reg[15:0] core_csr_reg_satp_asid ; reg[43:0] core_csr_reg_satp_ppn ; 
    reg core_csr_reg_wfi ; 
    wire core_csr__io_status_wfi_output = core_csr_reg_wfi ; reg[4:0] core_csr_reg_fflags ; reg[2:0] core_csr_reg_frm ; reg[2:0] core_csr_reg_mcountinhibit ; 
    wire core_csr_x3 = core_csr_reg_mcountinhibit [2]; reg[5:0] core_csr_small_0 ; 
    wire[6:0] core_csr_nextSmall ={1'h0, core_csr_small_0 }+{6'h0, core_csr_io_retire }; 
    wire core_csr__GEN_0 = core_csr_x3 ==1'h0; 
    wire[5:0] core_csr__GEN_1 = core_csr__GEN_0  ?  core_csr_nextSmall [5:0]: core_csr_small_0 ; reg[57:0] core_csr_large_0 ; 
    wire core_csr__GEN_2 = core_csr_nextSmall [6]& core_csr_x3 ==1'h0; 
    wire[58:0] core_csr__GEN_3 ={1'h0, core_csr_large_0 }+59'h1; 
    wire[57:0] core_csr__GEN_4 = core_csr__GEN_2  ?  core_csr__GEN_3 [57:0]: core_csr_large_0 ; 
    wire[63:0] core_csr_value ={ core_csr_large_0 , core_csr_small_0 }; 
    wire core_csr__io_csr_stall_output ; 
    wire core_csr_x10 = core_csr__io_csr_stall_output ==1'h0; 
    wire core_csr_x11 = core_csr_reg_mcountinhibit [0]; reg[5:0] core_csr_small_1 ; 
    wire[6:0] core_csr_nextSmall_1 ={1'h0, core_csr_small_1 }+{6'h0, core_csr_x10 }; 
    wire core_csr__GEN_5 = core_csr_x11 ==1'h0; 
    wire[5:0] core_csr__GEN_6 = core_csr__GEN_5  ?  core_csr_nextSmall_1 [5:0]: core_csr_small_1 ; reg[57:0] core_csr_large_1 ; 
    wire core_csr__GEN_7 = core_csr_nextSmall_1 [6]& core_csr_x11 ==1'h0; 
    wire[58:0] core_csr__GEN_8 ={1'h0, core_csr_large_1 }+59'h1; 
    wire[57:0] core_csr__GEN_9 = core_csr__GEN_7  ?  core_csr__GEN_8 [57:0]: core_csr_large_1 ; 
    wire[63:0] core_csr_value_1 ={ core_csr_large_1 , core_csr_small_1 }; 
    wire[1:0] core_csr_read_mip_lo_lo_lo ={ core_csr_mip_ssip , core_csr_mip_usip }; 
    wire[1:0] core_csr_read_mip_lo_lo_hi ={ core_csr_mip_msip , core_csr_mip_vssip }; 
    wire[3:0] core_csr_read_mip_lo_lo ={ core_csr_read_mip_lo_lo_hi , core_csr_read_mip_lo_lo_lo }; 
    wire[1:0] core_csr_read_mip_lo_hi_lo ={ core_csr_mip_stip , core_csr_mip_utip }; 
    wire[1:0] core_csr_read_mip_lo_hi_hi ={ core_csr_mip_mtip , core_csr_mip_vstip }; 
    wire[3:0] core_csr_read_mip_lo_hi ={ core_csr_read_mip_lo_hi_hi , core_csr_read_mip_lo_hi_lo }; 
    wire[7:0] core_csr_read_mip_lo ={ core_csr_read_mip_lo_hi , core_csr_read_mip_lo_lo }; 
    wire[1:0] core_csr_read_mip_hi_lo_lo ={ core_csr_mip_seip , core_csr_mip_ueip }; 
    wire[1:0] core_csr_read_mip_hi_lo_hi ={ core_csr_mip_meip , core_csr_mip_vseip }; 
    wire[3:0] core_csr_read_mip_hi_lo ={ core_csr_read_mip_hi_lo_hi , core_csr_read_mip_hi_lo_lo }; 
    wire[1:0] core_csr_read_mip_hi_hi_lo ={ core_csr_mip_rocc , core_csr_mip_sgeip }; 
    wire[1:0] core_csr_read_mip_hi_hi_hi ={ core_csr_mip_zero1 , core_csr_mip_debug }; 
    wire[3:0] core_csr_read_mip_hi_hi ={ core_csr_read_mip_hi_hi_hi , core_csr_read_mip_hi_hi_lo }; 
    wire[7:0] core_csr_read_mip_hi ={ core_csr_read_mip_hi_hi , core_csr_read_mip_hi_lo }; 
    wire[15:0] core_csr_read_mip ={ core_csr_read_mip_hi , core_csr_read_mip_lo }& core_csr_supported_interrupts ; 
    wire[15:0] core_csr_read_hip = core_csr_read_mip & core_csr_hs_delegable_interrupts ; 
    wire[63:0] core_csr_pending_interrupts ={48'h0, core_csr_read_mip }& core_csr_reg_mie |64'h0; 
    wire[14:0] core_csr_d_interrupts ={ core_csr_io_interrupts_debug ,14'h0}; 
    wire[63:0] core_csr_m_interrupts = core_csr_reg_rnmie &( core_csr_reg_mstatus_prv <=2'h1| core_csr_reg_mstatus_mie ) ? ~(~ core_csr_pending_interrupts | core_csr_read_mideleg ):64'h0; 
    wire[63:0] core_csr_s_interrupts = core_csr_reg_rnmie &( core_csr_reg_mstatus_v | core_csr_reg_mstatus_prv <2'h1| core_csr_reg_mstatus_prv ==2'h1& core_csr_reg_mstatus_sie ) ?  core_csr_pending_interrupts & core_csr_read_mideleg &~ core_csr_read_hideleg :64'h0; 
    wire[63:0] core_csr_vs_interrupts = core_csr_reg_rnmie & core_csr_reg_mstatus_v &( core_csr_reg_mstatus_prv <2'h1| core_csr_reg_mstatus_prv ==2'h1& core_csr_reg_vsstatus_sie ) ?  core_csr_pending_interrupts & core_csr_read_hideleg :64'h0; 
    wire core_csr_anyInterrupt = core_csr_d_interrupts [14]| core_csr_d_interrupts [13]| core_csr_d_interrupts [12]| core_csr_d_interrupts [11]| core_csr_d_interrupts [3]| core_csr_d_interrupts [7]| core_csr_d_interrupts [9]| core_csr_d_interrupts [1]| core_csr_d_interrupts [5]| core_csr_d_interrupts [10]| core_csr_d_interrupts [2]| core_csr_d_interrupts [6]| core_csr_d_interrupts [8]| core_csr_d_interrupts [0]| core_csr_d_interrupts [4]| core_csr_m_interrupts [15]| core_csr_m_interrupts [14]| core_csr_m_interrupts [13]| core_csr_m_interrupts [12]| core_csr_m_interrupts [11]| core_csr_m_interrupts [3]| core_csr_m_interrupts [7]| core_csr_m_interrupts [9]| core_csr_m_interrupts [1]| core_csr_m_interrupts [5]| core_csr_m_interrupts [10]| core_csr_m_interrupts [2]| core_csr_m_interrupts [6]| core_csr_m_interrupts [8]| core_csr_m_interrupts [0]| core_csr_m_interrupts [4]| core_csr_s_interrupts [15]| core_csr_s_interrupts [14]| core_csr_s_interrupts [13]| core_csr_s_interrupts [12]| core_csr_s_interrupts [11]| core_csr_s_interrupts [3]| core_csr_s_interrupts [7]| core_csr_s_interrupts [9]| core_csr_s_interrupts [1]| core_csr_s_interrupts [5]| core_csr_s_interrupts [10]| core_csr_s_interrupts [2]| core_csr_s_interrupts [6]| core_csr_s_interrupts [8]| core_csr_s_interrupts [0]| core_csr_s_interrupts [4]| core_csr_vs_interrupts [15]| core_csr_vs_interrupts [14]| core_csr_vs_interrupts [13]| core_csr_vs_interrupts [12]| core_csr_vs_interrupts [11]| core_csr_vs_interrupts [3]| core_csr_vs_interrupts [7]| core_csr_vs_interrupts [9]| core_csr_vs_interrupts [1]| core_csr_vs_interrupts [5]| core_csr_vs_interrupts [10]| core_csr_vs_interrupts [2]| core_csr_vs_interrupts [6]| core_csr_vs_interrupts [8]| core_csr_vs_interrupts [0]| core_csr_vs_interrupts [4]; 
    wire[3:0] core_csr_whichInterrupt = core_csr_d_interrupts [14] ? 4'hE: core_csr_d_interrupts [13] ? 4'hD: core_csr_d_interrupts [12] ? 4'hC: core_csr_d_interrupts [11] ? 4'hB: core_csr_d_interrupts [3] ? 4'h3: core_csr_d_interrupts [7] ? 4'h7: core_csr_d_interrupts [9] ? 4'h9: core_csr_d_interrupts [1] ? 4'h1: core_csr_d_interrupts [5] ? 4'h5: core_csr_d_interrupts [10] ? 4'hA: core_csr_d_interrupts [2] ? 4'h2: core_csr_d_interrupts [6] ? 4'h6: core_csr_d_interrupts [8] ? 4'h8: core_csr_d_interrupts [0] ? 4'h0: core_csr_d_interrupts [4] ? 4'h4: core_csr_m_interrupts [15] ? 4'hF: core_csr_m_interrupts [14] ? 4'hE: core_csr_m_interrupts [13] ? 4'hD: core_csr_m_interrupts [12] ? 4'hC: core_csr_m_interrupts [11] ? 4'hB: core_csr_m_interrupts [3] ? 4'h3: core_csr_m_interrupts [7] ? 4'h7: core_csr_m_interrupts [9] ? 4'h9: core_csr_m_interrupts [1] ? 4'h1: core_csr_m_interrupts [5] ? 4'h5: core_csr_m_interrupts [10] ? 4'hA: core_csr_m_interrupts [2] ? 4'h2: core_csr_m_interrupts [6] ? 4'h6: core_csr_m_interrupts [8] ? 4'h8: core_csr_m_interrupts [0] ? 4'h0: core_csr_m_interrupts [4] ? 4'h4: core_csr_s_interrupts [15] ? 4'hF: core_csr_s_interrupts [14] ? 4'hE: core_csr_s_interrupts [13] ? 4'hD: core_csr_s_interrupts [12] ? 4'hC: core_csr_s_interrupts [11] ? 4'hB: core_csr_s_interrupts [3] ? 4'h3: core_csr_s_interrupts [7] ? 4'h7: core_csr_s_interrupts [9] ? 4'h9: core_csr_s_interrupts [1] ? 4'h1: core_csr_s_interrupts [5] ? 4'h5: core_csr_s_interrupts [10] ? 4'hA: core_csr_s_interrupts [2] ? 4'h2: core_csr_s_interrupts [6] ? 4'h6: core_csr_s_interrupts [8] ? 4'h8: core_csr_s_interrupts [0] ? 4'h0: core_csr_s_interrupts [4] ? 4'h4: core_csr_vs_interrupts [15] ? 4'hF: core_csr_vs_interrupts [14] ? 4'hE: core_csr_vs_interrupts [13] ? 4'hD: core_csr_vs_interrupts [12] ? 4'hC: core_csr_vs_interrupts [11] ? 4'hB: core_csr_vs_interrupts [3] ? 4'h3: core_csr_vs_interrupts [7] ? 4'h7: core_csr_vs_interrupts [9] ? 4'h9: core_csr_vs_interrupts [1] ? 4'h1: core_csr_vs_interrupts [5] ? 4'h5: core_csr_vs_interrupts [10] ? 4'hA: core_csr_vs_interrupts [2] ? 4'h2: core_csr_vs_interrupts [6] ? 4'h6: core_csr_vs_interrupts [8] ? 4'h8:{1'h0, core_csr_vs_interrupts [0] ? 3'h0:3'h4}; 
    wire[64:0] core_csr__GEN_10 ={61'h0, core_csr_whichInterrupt }+65'h8000000000000000; 
    wire[63:0] core_csr_interruptCause = core_csr__GEN_10 [63:0]; 
    wire core_csr__io_singleStep_output ; 
    wire core_csr__io_status_cease_output ; 
    wire[30:0] core_csr_pmp_mask_base ={ core_csr_pmp_addr , core_csr_pmp_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_11 ={1'h0, core_csr_pmp_mask_base }+32'h1; 
    wire[32:0] core_csr__GEN_12 ={ core_csr_pmp_mask_base &~( core_csr__GEN_11 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_mask = core_csr__GEN_12 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_1 ={ core_csr_pmp_1_addr , core_csr_pmp_1_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_13 ={1'h0, core_csr_pmp_mask_base_1 }+32'h1; 
    wire[32:0] core_csr__GEN_14 ={ core_csr_pmp_mask_base_1 &~( core_csr__GEN_13 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_1_mask = core_csr__GEN_14 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_2 ={ core_csr_pmp_2_addr , core_csr_pmp_2_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_15 ={1'h0, core_csr_pmp_mask_base_2 }+32'h1; 
    wire[32:0] core_csr__GEN_16 ={ core_csr_pmp_mask_base_2 &~( core_csr__GEN_15 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_2_mask = core_csr__GEN_16 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_3 ={ core_csr_pmp_3_addr , core_csr_pmp_3_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_17 ={1'h0, core_csr_pmp_mask_base_3 }+32'h1; 
    wire[32:0] core_csr__GEN_18 ={ core_csr_pmp_mask_base_3 &~( core_csr__GEN_17 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_3_mask = core_csr__GEN_18 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_4 ={ core_csr_pmp_4_addr , core_csr_pmp_4_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_19 ={1'h0, core_csr_pmp_mask_base_4 }+32'h1; 
    wire[32:0] core_csr__GEN_20 ={ core_csr_pmp_mask_base_4 &~( core_csr__GEN_19 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_4_mask = core_csr__GEN_20 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_5 ={ core_csr_pmp_5_addr , core_csr_pmp_5_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_21 ={1'h0, core_csr_pmp_mask_base_5 }+32'h1; 
    wire[32:0] core_csr__GEN_22 ={ core_csr_pmp_mask_base_5 &~( core_csr__GEN_21 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_5_mask = core_csr__GEN_22 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_6 ={ core_csr_pmp_6_addr , core_csr_pmp_6_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_23 ={1'h0, core_csr_pmp_mask_base_6 }+32'h1; 
    wire[32:0] core_csr__GEN_24 ={ core_csr_pmp_mask_base_6 &~( core_csr__GEN_23 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_6_mask = core_csr__GEN_24 [31:0]; 
    wire[30:0] core_csr_pmp_mask_base_7 ={ core_csr_pmp_7_addr , core_csr_pmp_7_cfg_a [0]}; 
    wire[31:0] core_csr__GEN_25 ={1'h0, core_csr_pmp_mask_base_7 }+32'h1; 
    wire[32:0] core_csr__GEN_26 ={ core_csr_pmp_mask_base_7 &~( core_csr__GEN_25 [30:0]),2'h3}; 
    wire[31:0] core_csr_pmp_7_mask = core_csr__GEN_26 [31:0]; reg[63:0] core_csr_reg_misa ; 
    wire[1:0] core_csr_read_mstatus_lo_lo_lo_lo ={ core_csr__io_status_sie_output , core_csr__io_status_uie_output }; 
    wire[1:0] core_csr_read_mstatus_lo_lo_lo_hi ={ core_csr__io_status_mie_output , core_csr__io_status_hie_output }; 
    wire[3:0] core_csr_read_mstatus_lo_lo_lo ={ core_csr_read_mstatus_lo_lo_lo_hi , core_csr_read_mstatus_lo_lo_lo_lo }; 
    wire[1:0] core_csr_read_mstatus_lo_lo_hi_lo ={ core_csr__io_status_spie_output , core_csr__io_status_upie_output }; 
    wire[1:0] core_csr_read_mstatus_lo_lo_hi_hi_hi ={ core_csr__io_status_spp_output , core_csr__io_status_mpie_output }; 
    wire[2:0] core_csr_read_mstatus_lo_lo_hi_hi ={ core_csr_read_mstatus_lo_lo_hi_hi_hi , core_csr__io_status_ube_output }; 
    wire[4:0] core_csr_read_mstatus_lo_lo_hi ={ core_csr_read_mstatus_lo_lo_hi_hi , core_csr_read_mstatus_lo_lo_hi_lo }; 
    wire[8:0] core_csr_read_mstatus_lo_lo ={ core_csr_read_mstatus_lo_lo_hi , core_csr_read_mstatus_lo_lo_lo }; 
    wire[3:0] core_csr_read_mstatus_lo_hi_lo_lo ={ core_csr__io_status_mpp_output , core_csr__io_status_vs_output }; 
    wire[3:0] core_csr_read_mstatus_lo_hi_lo_hi ={ core_csr__io_status_xs_output , core_csr__io_status_fs_output }; 
    wire[7:0] core_csr_read_mstatus_lo_hi_lo ={ core_csr_read_mstatus_lo_hi_lo_hi , core_csr_read_mstatus_lo_hi_lo_lo }; 
    wire[1:0] core_csr_read_mstatus_lo_hi_hi_lo ={ core_csr__io_status_sum_output , core_csr__io_status_mprv_output }; 
    wire[1:0] core_csr_read_mstatus_lo_hi_hi_hi_hi ={ core_csr__io_status_tw_output , core_csr__io_status_tvm_output }; 
    wire[2:0] core_csr_read_mstatus_lo_hi_hi_hi ={ core_csr_read_mstatus_lo_hi_hi_hi_hi , core_csr__io_status_mxr_output }; 
    wire[4:0] core_csr_read_mstatus_lo_hi_hi ={ core_csr_read_mstatus_lo_hi_hi_hi , core_csr_read_mstatus_lo_hi_hi_lo }; 
    wire[12:0] core_csr_read_mstatus_lo_hi ={ core_csr_read_mstatus_lo_hi_hi , core_csr_read_mstatus_lo_hi_lo }; 
    wire[21:0] core_csr_read_mstatus_lo ={ core_csr_read_mstatus_lo_hi , core_csr_read_mstatus_lo_lo }; 
    wire[8:0] core_csr_read_mstatus_hi_lo_lo_lo ={ core_csr__io_status_zero1_output , core_csr__io_status_tsr_output }; 
    wire[1:0] core_csr__io_status_uxl_output =2'h0; 
    wire[2:0] core_csr_read_mstatus_hi_lo_lo_hi ={ core_csr__io_status_uxl_output , core_csr__io_status_sd_rv32_output }; 
    wire[11:0] core_csr_read_mstatus_hi_lo_lo ={ core_csr_read_mstatus_hi_lo_lo_hi , core_csr_read_mstatus_hi_lo_lo_lo }; 
    wire[1:0] core_csr__io_status_sxl_output =2'h0; 
    wire[2:0] core_csr_read_mstatus_hi_lo_hi_lo ={ core_csr__io_status_sbe_output , core_csr__io_status_sxl_output }; 
    wire[1:0] core_csr_read_mstatus_hi_lo_hi_hi_hi ={ core_csr__io_status_mpv_output , core_csr__io_status_gva_output }; 
    wire[2:0] core_csr_read_mstatus_hi_lo_hi_hi ={ core_csr_read_mstatus_hi_lo_hi_hi_hi , core_csr__io_status_mbe_output }; 
    wire[5:0] core_csr_read_mstatus_hi_lo_hi ={ core_csr_read_mstatus_hi_lo_hi_hi , core_csr_read_mstatus_hi_lo_hi_lo }; 
    wire[17:0] core_csr_read_mstatus_hi_lo ={ core_csr_read_mstatus_hi_lo_hi , core_csr_read_mstatus_hi_lo_lo }; 
    wire core_csr__io_status_sd_output ; 
    wire[23:0] core_csr_read_mstatus_hi_hi_lo_lo ={ core_csr__io_status_sd_output , core_csr__io_status_zero2_output }; 
    wire core_csr__io_status_dv_output ; 
    wire[2:0] core_csr_read_mstatus_hi_hi_lo_hi_hi ={ core_csr__io_status_dv_output , core_csr__io_status_prv_output }; 
    wire[3:0] core_csr_read_mstatus_hi_hi_lo_hi ={ core_csr_read_mstatus_hi_hi_lo_hi_hi , core_csr__io_status_v_output }; 
    wire[27:0] core_csr_read_mstatus_hi_hi_lo ={ core_csr_read_mstatus_hi_hi_lo_hi , core_csr_read_mstatus_hi_hi_lo_lo }; 
    wire[31:0] core_csr__io_status_isa_output ; 
    wire[1:0] core_csr__io_status_dprv_output ; 
    wire[33:0] core_csr_read_mstatus_hi_hi_hi_lo ={ core_csr__io_status_isa_output , core_csr__io_status_dprv_output }; 
    wire[1:0] core_csr_read_mstatus_hi_hi_hi_hi_hi ={ core_csr__io_status_debug_output , core_csr__io_status_cease_output }; 
    wire[2:0] core_csr_read_mstatus_hi_hi_hi_hi ={ core_csr_read_mstatus_hi_hi_hi_hi_hi , core_csr__io_status_wfi_output }; 
    wire[36:0] core_csr_read_mstatus_hi_hi_hi ={ core_csr_read_mstatus_hi_hi_hi_hi , core_csr_read_mstatus_hi_hi_hi_lo }; 
    wire[64:0] core_csr_read_mstatus_hi_hi ={ core_csr_read_mstatus_hi_hi_hi , core_csr_read_mstatus_hi_hi_lo }; 
    wire[82:0] core_csr_read_mstatus_hi ={ core_csr_read_mstatus_hi_hi , core_csr_read_mstatus_hi_lo }; 
    wire[104:0] core_csr__GEN_27 ={ core_csr_read_mstatus_hi , core_csr_read_mstatus_lo }; 
    wire[63:0] core_csr_read_mstatus = core_csr__GEN_27 [63:0]; 
    wire[63:0] core_csr_read_mtvec ={32'h0, core_csr_reg_mtvec &~{24'h0, core_csr_reg_mtvec [0] ? 8'hFE:8'h2}}; 
    wire[32:0] core_csr__GEN_28 = core_csr_reg_stvec &~{25'h0, core_csr_reg_stvec [0] ? 8'hFE:8'h2}; 
    wire[63:0] core_csr_read_stvec ={ core_csr__GEN_28 [32] ? 31'h7FFFFFFF:31'h0, core_csr__GEN_28 }; reg[3:0] core_csr_casez_tmp ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_0 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_0  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_0  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_1 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_1  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_1  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_2 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_2  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_2  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_3 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_3  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_3  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_4 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_4  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_4  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_5 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_5  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_5  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_6 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_6  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_6  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_7 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_7  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_7  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_8 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_8  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_8  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_9 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_9  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_9  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_10 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_10  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_10  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_11 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_11  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_11  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_12 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_12  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_12  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_13 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_13  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_13  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_14 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_14  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_14  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_15 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_15  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_15  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_16 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_16  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_16  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_17 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_17  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_17  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_18 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_18  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_18  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_19 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_19  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_19  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_20 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_20  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_20  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_21 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_21  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_21  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_22 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_22  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_22  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_23 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_23  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_23  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_24 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_24  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_24  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_25 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_25  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_25  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_26 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_26  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_26  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_27 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_27  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_27  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_28 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_28  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_28  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_29 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_29  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_29  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_30 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_30  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_30  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_31 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_31  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_31  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_32 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_32  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_32  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_33 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_33  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_33  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_34 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_34  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_34  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_35 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_35  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_35  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_36 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_36  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_36  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_37 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_37  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_37  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_38 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_38  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_38  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[1:0] core_csr_lo_lo_hi_4 ={ core_csr_casez_tmp_11 , core_csr_casez_tmp_32 }; reg[3:0] core_csr_casez_tmp_39 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_39  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_39  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_40 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_40  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_40  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_41 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_41  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_41  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_42 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_42  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_42  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_43 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_43  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_43  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_44 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_44  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_44  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_45 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_45  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_45  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_46 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_46  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_46  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_47 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_47  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_47  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_48 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_48  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_48  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_49 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_49  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_49  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_50 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_50  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_50  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_51 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_51  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_51  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_52 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_52  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_52  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_53 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_53  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_53  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_54 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_54  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_54  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_55 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_55  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_55  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_56 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_56  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_56  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_57 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_57  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_57  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_58 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_58  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_58  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[2:0] core_csr_lo_lo_4 ={ core_csr_lo_lo_hi_4 , core_csr_casez_tmp_53 }; reg[3:0] core_csr_casez_tmp_59 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_59  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_59  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_60 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_60  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_60  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_61 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_61  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_61  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_62 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_62  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_62  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_63 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_63  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_63  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_64 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_64  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_64  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_65 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_65  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_65  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_66 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_66  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_66  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_67 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_67  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_67  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_68 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_68  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_68  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_69 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_69  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_69  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_70 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_70  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_70  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_71 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_71  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_71  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_72 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_72  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_72  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_73 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_73  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_73  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_74 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_74  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_74  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_75 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_75  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_75  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_76 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_76  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_76  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_77 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_77  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_77  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_78 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_78  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_78  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_79 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_79  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_79  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_80 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_80  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_80  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_81 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_81  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_81  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_82 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_82  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_82  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_83 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_83  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_83  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_84 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_84  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_84  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_85 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_85  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_85  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_86 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_86  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_86  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_87 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_87  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_87  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_88 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_88  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_88  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_89 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_89  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_89  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_90 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_90  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_90  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_91 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_91  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_91  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_92 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_92  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_92  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_93 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_93  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_93  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_94 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_94  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_94  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_95 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_95  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_95  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_96 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_96  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_96  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_97 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_97  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_97  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_98 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_98  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_98  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[1:0] core_csr_lo_hi_lo_4 ={ core_csr_casez_tmp_69 , core_csr_casez_tmp_90 }; reg[3:0] core_csr_casez_tmp_99 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_99  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_99  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_100 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_100  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_100  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_101 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_101  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_101  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_102 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_102  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_102  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_103 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_103  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_103  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_104 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_104  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_104  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_105 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_105  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_105  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_106 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_106  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_106  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_107 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_107  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_107  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_108 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_108  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_108  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_109 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_109  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_109  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_110 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_110  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_110  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_111 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_111  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_111  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_112 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_112  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_112  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_113 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_113  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_113  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_114 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_114  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_114  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_115 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_115  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_115  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_116 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_116  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_116  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_117 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_117  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_117  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_118 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_118  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_118  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_119 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_119  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_119  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_120 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_120  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_120  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_121 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_121  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_121  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_122 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_122  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_122  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_123 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_123  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_123  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_124 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_124  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_124  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_125 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_125  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_125  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_126 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_126  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_126  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_127 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_127  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_127  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_128 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_128  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_128  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_129 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_129  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_129  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_130 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_130  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_130  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_131 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_131  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_131  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_132 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_132  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_132  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_133 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_133  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_133  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_134 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_134  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_134  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_135 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_135  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_135  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_136 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_136  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_136  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_137 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_137  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_137  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_138 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_138  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_138  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[1:0] core_csr_lo_hi_hi_4 ={ core_csr_casez_tmp_107 , core_csr_casez_tmp_128 }; 
    wire[3:0] core_csr_lo_hi_4 ={ core_csr_lo_hi_hi_4 , core_csr_lo_hi_lo_4 }; 
    wire[6:0] core_csr_lo_4 ={ core_csr_lo_hi_4 , core_csr_lo_lo_4 }; reg[3:0] core_csr_casez_tmp_139 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_139  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_139  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_140 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_140  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_140  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_141 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_141  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_141  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_142 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_142  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_142  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_143 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_143  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_143  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_144 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_144  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_144  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_145 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_145  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_145  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_146 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_146  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_146  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_147 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_147  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_147  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_148 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_148  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_148  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_149 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_149  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_149  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_150 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_150  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_150  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_151 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_151  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_151  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_152 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_152  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_152  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_153 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_153  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_153  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_154 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_154  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_154  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_155 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_155  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_155  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_156 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_156  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_156  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_157 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_157  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_157  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_158 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_158  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_158  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_159 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_159  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_159  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_160 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_160  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_160  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_161 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_161  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_161  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_162 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_162  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_162  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_163 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_163  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_163  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_164 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_164  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_164  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_165 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_165  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_165  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_166 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_166  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_166  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_167 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_167  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_167  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_168 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_168  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_168  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_169 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_169  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_169  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_170 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_170  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_170  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_171 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_171  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_171  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_172 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_172  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_172  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_173 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_173  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_173  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_174 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_174  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_174  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_175 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_175  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_175  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_176 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_176  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_176  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_177 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_177  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_177  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_178 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_178  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_178  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[3:0] core_csr_hi_lo_lo_4 ={ core_csr_casez_tmp_145 , core_csr_casez_tmp_166 }; reg[3:0] core_csr_casez_tmp_179 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_179  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_179  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_180 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_180  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_180  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_181 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_181  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_181  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_182 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_182  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_182  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_183 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_183  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_183  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_184 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_184  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_184  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_185 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_185  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_185  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_186 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_186  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_186  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_187 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_187  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_187  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_188 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_188  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_188  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_189 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_189  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_189  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_190 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_190  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_190  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_191 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_191  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_191  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_192 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_192  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_192  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_193 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_193  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_193  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_194 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_194  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_194  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_195 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_195  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_195  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_196 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_196  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_196  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_197 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_197  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_197  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_198 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_198  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_198  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_199 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_199  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_199  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_200 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_200  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_200  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_201 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_201  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_201  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_202 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_202  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_202  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_203 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_203  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_203  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_204 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_204  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_204  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_205 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_205  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_205  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_206 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_206  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_206  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_207 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_207  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_207  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_208 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_208  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_208  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_209 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_209  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_209  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_210 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_210  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_210  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_211 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_211  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_211  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_212 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_212  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_212  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_213 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_213  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_213  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_214 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_214  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_214  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_215 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_215  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_215  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_216 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_216  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_216  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_217 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_217  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_217  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_218 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_218  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_218  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[1:0] core_csr_hi_lo_hi_4 ={ core_csr_casez_tmp_183 , core_csr_casez_tmp_204 }; 
    wire[5:0] core_csr_hi_lo_4 ={ core_csr_hi_lo_hi_4 , core_csr_hi_lo_lo_4 }; reg[3:0] core_csr_casez_tmp_219 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_219  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_219  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_220 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_220  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_220  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_221 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_221  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_221  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_222 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_222  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_222  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_223 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_223  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_223  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_224 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_224  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_224  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_225 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_225  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_225  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_226 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_226  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_226  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_227 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_227  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_227  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_228 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_228  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_228  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_229 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_229  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_229  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_230 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_230  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_230  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_231 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_231  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_231  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_232 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_232  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_232  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_233 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_233  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_233  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_234 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_234  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_234  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_235 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_235  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_235  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_236 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_236  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_236  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_237 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_237  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_237  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_238 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_238  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_238  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_239 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_239  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_239  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_240 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_240  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_240  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_241 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_241  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_241  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_242 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_242  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_242  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_243 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_243  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_243  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_244 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_244  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_244  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_245 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_245  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_245  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_246 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_246  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_246  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_247 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_247  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_247  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_248 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_248  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_248  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_249 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_249  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_249  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_250 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_250  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_250  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_251 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_251  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_251  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_252 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_252  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_252  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_253 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_253  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_253  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_254 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_254  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_254  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_255 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_255  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_255  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_256 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_256  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_256  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_257 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_257  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_257  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_258 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_258  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_258  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[45:0] core_csr_hi_hi_lo_4 ={ core_csr_casez_tmp_221 , core_csr_casez_tmp_242 }; reg[3:0] core_csr_casez_tmp_259 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_259  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_259  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_260 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_260  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_260  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_261 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_261  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_261  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_262 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_262  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_262  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_263 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_263  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_263  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_264 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_264  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_264  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_265 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_265  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_265  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_266 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_266  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_266  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_267 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_267  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_267  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_268 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_268  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_268  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_269 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_269  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_269  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_270 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_270  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_270  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_271 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_271  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_271  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_272 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_272  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_272  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_273 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_273  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_273  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_274 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_274  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_274  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_275 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_275  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_275  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_276 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_276  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_276  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_277 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_277  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_277  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_278 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_278  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_278  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_279 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_279  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_279  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_280 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_280  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_280  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_281 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_281  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_281  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_282 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_282  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_282  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_283 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_283  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_283  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_284 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_284  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_284  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_285 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_285  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_285  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_286 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_286  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_286  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_287 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_287  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_287  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_288 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_288  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_288  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_289 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_289  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_289  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_290 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_290  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_290  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_291 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_291  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_291  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_292 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_292  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_292  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_293 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_293  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_293  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_294 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_294  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_294  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_295 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_295  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_295  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_296 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_296  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_296  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_297 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_297  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_297  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_298 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_298  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_298  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[4:0] core_csr_hi_hi_hi_4 ={ core_csr_casez_tmp_259 , core_csr_casez_tmp_280 }; 
    wire[50:0] core_csr_hi_hi_4 ={ core_csr_hi_hi_hi_4 , core_csr_hi_hi_lo_4 }; 
    wire[56:0] core_csr_hi_4 ={ core_csr_hi_hi_4 , core_csr_hi_lo_4 }; reg[3:0] core_csr_casez_tmp_299 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_299  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_299  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_300 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_300  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_300  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_301 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_301  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_301  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_302 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_302  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_302  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_303 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_303  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_303  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_304 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_304  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_304  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_305 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_305  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_305  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_306 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_306  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_306  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_307 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_307  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_307  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_308 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_308  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_308  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_309 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_309  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_309  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_310 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_310  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_310  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_311 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_311  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_311  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_312 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_312  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_312  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_313 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_313  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_313  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_314 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_314  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_314  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_315 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_315  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_315  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_316 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_316  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_316  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_317 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_317  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_317  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_318 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_318  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_318  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_319 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_319  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_319  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_320 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_320  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_320  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_321 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_321  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_321  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_322 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_322  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_322  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_323 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_323  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_323  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_324 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_324  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_324  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_325 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_325  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_325  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_326 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_326  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_326  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_327 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_327  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_327  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_328 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_328  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_328  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_329 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_329  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_329  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_330 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_330  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_330  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_331 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_331  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_331  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_332 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_332  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_332  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_333 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_333  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_333  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_334 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_334  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_334  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_335 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_335  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_335  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_336 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_336  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_336  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_337 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_337  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_337  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_338 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_338  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_338  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_339 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_339  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_339  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_340 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_340  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_340  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_341 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_341  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_341  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_342 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_342  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_342  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_343 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_343  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_343  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_344 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_344  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_344  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_345 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_345  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_345  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_346 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_346  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_346  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_347 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_347  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_347  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_348 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_348  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_348  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_349 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_349  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_349  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_350 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_350  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_350  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_351 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_351  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_351  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_352 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_352  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_352  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_353 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_353  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_353  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_354 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_354  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_354  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_355 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_355  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_355  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_356 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_356  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_356  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_357 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_357  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_357  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_358 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_358  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_358  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_359 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_359  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_359  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_360 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_360  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_360  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_361 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_361  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_361  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_362 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_362  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_362  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_363 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_363  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_363  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_364 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_364  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_364  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_365 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_365  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_365  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_366 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_366  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_366  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_367 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_367  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_367  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_368 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_368  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_368  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_369 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_369  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_369  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_370 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_370  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_370  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_371 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_371  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_371  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_372 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_372  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_372  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_373 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_373  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_373  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_374 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_374  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_374  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_375 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_375  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_375  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_376 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_376  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_376  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_377 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_377  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_377  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    wire core_csr_lo_hi_5 = core_csr_casez_tmp_377 ; 
    reg core_csr_casez_tmp_378 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_378  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_378  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_379 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_379  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_379  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_380 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_380  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_380  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_381 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_381  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_381  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_382 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_382  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_382  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_383 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_383  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_383  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_384 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_384  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_384  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_385 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_385  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_385  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_386 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_386  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_386  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_387 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_387  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_387  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_388 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_388  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_388  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_389 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_389  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_389  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_390 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_390  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_390  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_391 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_391  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_391  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_392 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_392  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_392  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_393 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_393  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_393  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_394 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_394  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_394  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_395 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_395  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_395  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_396 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_396  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_396  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_397 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_397  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_397  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_398 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_398  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_398  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[1:0] core_csr_lo_5 ={ core_csr_lo_hi_5 , core_csr_casez_tmp_398 }; reg[3:0] core_csr_casez_tmp_399 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_399  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_399  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_400 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_400  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_400  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_401 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_401  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_401  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_402 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_402  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_402  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_403 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_403  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_403  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_404 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_404  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_404  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_405 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_405  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_405  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_406 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_406  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_406  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_407 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_407  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_407  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_408 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_408  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_408  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_409 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_409  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_409  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_410 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_410  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_410  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_411 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_411  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_411  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_412 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_412  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_412  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_413 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_413  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_413  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_414 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_414  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_414  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_415 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_415  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_415  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_416 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_416  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_416  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_417 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_417  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_417  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_418 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_418  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_418  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_419 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_419  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_419  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_420 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_420  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_420  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_421 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_421  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_421  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_422 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_422  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_422  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_423 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_423  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_423  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_424 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_424  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_424  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_425 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_425  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_425  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_426 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_426  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_426  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_427 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_427  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_427  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_428 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_428  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_428  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_429 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_429  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_429  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_430 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_430  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_430  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_431 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_431  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_431  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_432 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_432  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_432  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_433 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_433  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_433  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_434 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_434  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_434  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_435 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_435  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_435  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
    wire core_csr_hi_hi_5 = core_csr_casez_tmp_435 ; reg[47:0] core_csr_casez_tmp_436 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_436  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_436  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_437 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_437  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_437  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_438 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_438  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_438  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
  reg[3:0] core_csr_casez_tmp_439 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_439  = core_csr_reg_bp_0_control_ttype ;
              default : 
                  core_csr_casez_tmp_439  = core_csr_reg_bp_1_control_ttype ;endcase
         end
    reg core_csr_casez_tmp_440 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_440  = core_csr_reg_bp_0_control_dmode ;
              default : 
                  core_csr_casez_tmp_440  = core_csr_reg_bp_1_control_dmode ;endcase
         end
  reg[5:0] core_csr_casez_tmp_441 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_441  = core_csr_reg_bp_0_control_maskmax ;
              default : 
                  core_csr_casez_tmp_441  = core_csr_reg_bp_1_control_maskmax ;endcase
         end
  reg[39:0] core_csr_casez_tmp_442 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_442  = core_csr_reg_bp_0_control_reserved ;
              default : 
                  core_csr_casez_tmp_442  = core_csr_reg_bp_1_control_reserved ;endcase
         end
    reg core_csr_casez_tmp_443 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_443  = core_csr_reg_bp_0_control_action ;
              default : 
                  core_csr_casez_tmp_443  = core_csr_reg_bp_1_control_action ;endcase
         end
    reg core_csr_casez_tmp_444 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_444  = core_csr_reg_bp_0_control_chain ;
              default : 
                  core_csr_casez_tmp_444  = core_csr_reg_bp_1_control_chain ;endcase
         end
  reg[1:0] core_csr_casez_tmp_445 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_445  = core_csr_reg_bp_0_control_zero ;
              default : 
                  core_csr_casez_tmp_445  = core_csr_reg_bp_1_control_zero ;endcase
         end
  reg[1:0] core_csr_casez_tmp_446 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_446  = core_csr_reg_bp_0_control_tmatch ;
              default : 
                  core_csr_casez_tmp_446  = core_csr_reg_bp_1_control_tmatch ;endcase
         end
    reg core_csr_casez_tmp_447 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_447  = core_csr_reg_bp_0_control_m ;
              default : 
                  core_csr_casez_tmp_447  = core_csr_reg_bp_1_control_m ;endcase
         end
    reg core_csr_casez_tmp_448 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_448  = core_csr_reg_bp_0_control_h ;
              default : 
                  core_csr_casez_tmp_448  = core_csr_reg_bp_1_control_h ;endcase
         end
    reg core_csr_casez_tmp_449 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_449  = core_csr_reg_bp_0_control_s ;
              default : 
                  core_csr_casez_tmp_449  = core_csr_reg_bp_1_control_s ;endcase
         end
    reg core_csr_casez_tmp_450 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_450  = core_csr_reg_bp_0_control_u ;
              default : 
                  core_csr_casez_tmp_450  = core_csr_reg_bp_1_control_u ;endcase
         end
    reg core_csr_casez_tmp_451 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_451  = core_csr_reg_bp_0_control_x ;
              default : 
                  core_csr_casez_tmp_451  = core_csr_reg_bp_1_control_x ;endcase
         end
    reg core_csr_casez_tmp_452 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_452  = core_csr_reg_bp_0_control_w ;
              default : 
                  core_csr_casez_tmp_452  = core_csr_reg_bp_1_control_w ;endcase
         end
    reg core_csr_casez_tmp_453 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_453  = core_csr_reg_bp_0_control_r ;
              default : 
                  core_csr_casez_tmp_453  = core_csr_reg_bp_1_control_r ;endcase
         end
  reg[32:0] core_csr_casez_tmp_454 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_454  = core_csr_reg_bp_0_address ;
              default : 
                  core_csr_casez_tmp_454  = core_csr_reg_bp_1_address ;endcase
         end
    reg core_csr_casez_tmp_455 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_455  = core_csr_reg_bp_0_textra_mselect ;
              default : 
                  core_csr_casez_tmp_455  = core_csr_reg_bp_1_textra_mselect ;endcase
         end
  reg[47:0] core_csr_casez_tmp_456 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_456  = core_csr_reg_bp_0_textra_pad2 ;
              default : 
                  core_csr_casez_tmp_456  = core_csr_reg_bp_1_textra_pad2 ;endcase
         end
    reg core_csr_casez_tmp_457 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_457  = core_csr_reg_bp_0_textra_pad1 ;
              default : 
                  core_csr_casez_tmp_457  = core_csr_reg_bp_1_textra_pad1 ;endcase
         end
    reg core_csr_casez_tmp_458 ; 
  always @(*)
         begin 
             casez ( core_csr_reg_tselect )
              1 'b0: 
                  core_csr_casez_tmp_458  = core_csr_reg_bp_0_textra_sselect ;
              default : 
                  core_csr_casez_tmp_458  = core_csr_reg_bp_1_textra_sselect ;endcase
         end
    wire[48:0] core_csr_hi_5 ={ core_csr_hi_hi_5 , core_csr_casez_tmp_456 }; 
    wire[33:0] core_csr__GEN_29 =~(~ core_csr_reg_mepc |{32'h0, core_csr_reg_misa [2] ? 2'h1:2'h3}); 
    wire[2:0] core_csr_lo_lo_hi_5 ={ core_csr_reg_dcsr_zero1 , core_csr_reg_dcsr_step }; 
    wire[4:0] core_csr_lo_lo_5 ={ core_csr_lo_lo_hi_5 , core_csr_reg_dcsr_prv }; 
    wire[3:0] core_csr_lo_hi_lo_5 ={ core_csr_reg_dcsr_cause , core_csr_reg_dcsr_v }; 
    wire[1:0] core_csr_lo_hi_hi_5 ={ core_csr_reg_dcsr_stopcycle , core_csr_reg_dcsr_stoptime }; 
    wire[5:0] core_csr_lo_hi_6 ={ core_csr_lo_hi_hi_5 , core_csr_lo_hi_lo_5 }; 
    wire[10:0] core_csr_lo_6 ={ core_csr_lo_hi_6 , core_csr_lo_lo_5 }; 
    wire[1:0] core_csr_hi_lo_lo_5 ={ core_csr_reg_dcsr_ebreaku , core_csr_reg_dcsr_zero2 }; 
    wire[1:0] core_csr_hi_lo_hi_5 ={ core_csr_reg_dcsr_ebreakh , core_csr_reg_dcsr_ebreaks }; 
    wire[3:0] core_csr_hi_lo_5 ={ core_csr_hi_lo_hi_5 , core_csr_hi_lo_lo_5 }; 
    wire[12:0] core_csr_hi_hi_lo_5 ={ core_csr_reg_dcsr_zero3 , core_csr_reg_dcsr_ebreakm }; 
    wire[3:0] core_csr_hi_hi_hi_5 ={ core_csr_reg_dcsr_xdebugver , core_csr_reg_dcsr_zero4 }; 
    wire[16:0] core_csr_hi_hi_6 ={ core_csr_hi_hi_hi_5 , core_csr_hi_hi_lo_5 }; 
    wire[20:0] core_csr_hi_6 ={ core_csr_hi_hi_6 , core_csr_hi_lo_5 }; 
    wire[33:0] core_csr__GEN_30 =~(~ core_csr_reg_dpc |{32'h0, core_csr_reg_misa [2] ? 2'h1:2'h3}); 
    wire[2:0] core_csr_read_mnstatus_zero3 = core_csr__read_mnstatus_WIRE_zero3 ; 
    wire[2:0] core_csr_read_mnstatus_zero2 = core_csr__read_mnstatus_WIRE_zero2 ; 
    wire[2:0] core_csr_read_mnstatus_zero1 = core_csr__read_mnstatus_WIRE_zero1 ; 
    wire[7:0] core_csr_read_fcsr ={ core_csr_reg_frm , core_csr_reg_fflags }; 
    wire core_csr_sie_mask_sgeip_mask_zero1 = core_csr__sie_mask_sgeip_mask_WIRE_zero1 ; 
    wire core_csr_sie_mask_sgeip_mask_debug = core_csr__sie_mask_sgeip_mask_WIRE_debug ; 
    wire core_csr_sie_mask_sgeip_mask_rocc = core_csr__sie_mask_sgeip_mask_WIRE_rocc ; 
    wire core_csr_sie_mask_sgeip_mask_meip = core_csr__sie_mask_sgeip_mask_WIRE_meip ; 
    wire core_csr_sie_mask_sgeip_mask_vseip = core_csr__sie_mask_sgeip_mask_WIRE_vseip ; 
    wire core_csr_sie_mask_sgeip_mask_seip = core_csr__sie_mask_sgeip_mask_WIRE_seip ; 
    wire core_csr_sie_mask_sgeip_mask_ueip = core_csr__sie_mask_sgeip_mask_WIRE_ueip ; 
    wire core_csr_sie_mask_sgeip_mask_mtip = core_csr__sie_mask_sgeip_mask_WIRE_mtip ; 
    wire core_csr_sie_mask_sgeip_mask_vstip = core_csr__sie_mask_sgeip_mask_WIRE_vstip ; 
    wire core_csr_sie_mask_sgeip_mask_stip = core_csr__sie_mask_sgeip_mask_WIRE_stip ; 
    wire core_csr_sie_mask_sgeip_mask_utip = core_csr__sie_mask_sgeip_mask_WIRE_utip ; 
    wire core_csr_sie_mask_sgeip_mask_msip = core_csr__sie_mask_sgeip_mask_WIRE_msip ; 
    wire core_csr_sie_mask_sgeip_mask_vssip = core_csr__sie_mask_sgeip_mask_WIRE_vssip ; 
    wire core_csr_sie_mask_sgeip_mask_ssip = core_csr__sie_mask_sgeip_mask_WIRE_ssip ; 
    wire core_csr_sie_mask_sgeip_mask_usip = core_csr__sie_mask_sgeip_mask_WIRE_usip ; 
    wire[1:0] core_csr_sie_mask_lo_lo_lo ={ core_csr_sie_mask_sgeip_mask_ssip , core_csr_sie_mask_sgeip_mask_usip }; 
    wire[1:0] core_csr_sie_mask_lo_lo_hi ={ core_csr_sie_mask_sgeip_mask_msip , core_csr_sie_mask_sgeip_mask_vssip }; 
    wire[3:0] core_csr_sie_mask_lo_lo ={ core_csr_sie_mask_lo_lo_hi , core_csr_sie_mask_lo_lo_lo }; 
    wire[1:0] core_csr_sie_mask_lo_hi_lo ={ core_csr_sie_mask_sgeip_mask_stip , core_csr_sie_mask_sgeip_mask_utip }; 
    wire[1:0] core_csr_sie_mask_lo_hi_hi ={ core_csr_sie_mask_sgeip_mask_mtip , core_csr_sie_mask_sgeip_mask_vstip }; 
    wire[3:0] core_csr_sie_mask_lo_hi ={ core_csr_sie_mask_lo_hi_hi , core_csr_sie_mask_lo_hi_lo }; 
    wire[7:0] core_csr_sie_mask_lo ={ core_csr_sie_mask_lo_hi , core_csr_sie_mask_lo_lo }; 
    wire[1:0] core_csr_sie_mask_hi_lo_lo ={ core_csr_sie_mask_sgeip_mask_seip , core_csr_sie_mask_sgeip_mask_ueip }; 
    wire[1:0] core_csr_sie_mask_hi_lo_hi ={ core_csr_sie_mask_sgeip_mask_meip , core_csr_sie_mask_sgeip_mask_vseip }; 
    wire[3:0] core_csr_sie_mask_hi_lo ={ core_csr_sie_mask_hi_lo_hi , core_csr_sie_mask_hi_lo_lo }; 
    wire[1:0] core_csr_sie_mask_hi_hi_lo ={ core_csr_sie_mask_sgeip_mask_rocc , core_csr_sie_mask_sgeip_mask_sgeip }; 
    wire[1:0] core_csr_sie_mask_hi_hi_hi ={ core_csr_sie_mask_sgeip_mask_zero1 , core_csr_sie_mask_sgeip_mask_debug }; 
    wire[3:0] core_csr_sie_mask_hi_hi ={ core_csr_sie_mask_hi_hi_hi , core_csr_sie_mask_hi_hi_lo }; 
    wire[7:0] core_csr_sie_mask_hi ={ core_csr_sie_mask_hi_hi , core_csr_sie_mask_hi_lo }; 
    wire[63:0] core_csr_sie_mask = core_csr_read_mideleg &{48'h0,~( core_csr_hs_delegable_interrupts |{ core_csr_sie_mask_hi , core_csr_sie_mask_lo })}; 
    wire[1:0] core_csr_lo_hi_7 ={ core_csr_reg_pmp_0_cfg_x , core_csr_reg_pmp_0_cfg_w }; 
    wire[2:0] core_csr_lo_7 ={ core_csr_lo_hi_7 , core_csr_reg_pmp_0_cfg_r }; 
    wire[2:0] core_csr_hi_hi_7 ={ core_csr_reg_pmp_0_cfg_l , core_csr_reg_pmp_0_cfg_res }; 
    wire[4:0] core_csr_hi_7 ={ core_csr_hi_hi_7 , core_csr_reg_pmp_0_cfg_a }; 
    wire[1:0] core_csr_lo_hi_8 ={ core_csr_reg_pmp_1_cfg_x , core_csr_reg_pmp_1_cfg_w }; 
    wire[2:0] core_csr_lo_8 ={ core_csr_lo_hi_8 , core_csr_reg_pmp_1_cfg_r }; 
    wire[2:0] core_csr_hi_hi_8 ={ core_csr_reg_pmp_1_cfg_l , core_csr_reg_pmp_1_cfg_res }; 
    wire[4:0] core_csr_hi_8 ={ core_csr_hi_hi_8 , core_csr_reg_pmp_1_cfg_a }; 
    wire[1:0] core_csr_lo_hi_9 ={ core_csr_reg_pmp_2_cfg_x , core_csr_reg_pmp_2_cfg_w }; 
    wire[2:0] core_csr_lo_9 ={ core_csr_lo_hi_9 , core_csr_reg_pmp_2_cfg_r }; 
    wire[2:0] core_csr_hi_hi_9 ={ core_csr_reg_pmp_2_cfg_l , core_csr_reg_pmp_2_cfg_res }; 
    wire[4:0] core_csr_hi_9 ={ core_csr_hi_hi_9 , core_csr_reg_pmp_2_cfg_a }; 
    wire[1:0] core_csr_lo_hi_10 ={ core_csr_reg_pmp_3_cfg_x , core_csr_reg_pmp_3_cfg_w }; 
    wire[2:0] core_csr_lo_10 ={ core_csr_lo_hi_10 , core_csr_reg_pmp_3_cfg_r }; 
    wire[2:0] core_csr_hi_hi_10 ={ core_csr_reg_pmp_3_cfg_l , core_csr_reg_pmp_3_cfg_res }; 
    wire[4:0] core_csr_hi_10 ={ core_csr_hi_hi_10 , core_csr_reg_pmp_3_cfg_a }; 
    wire[1:0] core_csr_lo_hi_11 ={ core_csr_reg_pmp_4_cfg_x , core_csr_reg_pmp_4_cfg_w }; 
    wire[2:0] core_csr_lo_11 ={ core_csr_lo_hi_11 , core_csr_reg_pmp_4_cfg_r }; 
    wire[2:0] core_csr_hi_hi_11 ={ core_csr_reg_pmp_4_cfg_l , core_csr_reg_pmp_4_cfg_res }; 
    wire[4:0] core_csr_hi_11 ={ core_csr_hi_hi_11 , core_csr_reg_pmp_4_cfg_a }; 
    wire[1:0] core_csr_lo_hi_12 ={ core_csr_reg_pmp_5_cfg_x , core_csr_reg_pmp_5_cfg_w }; 
    wire[2:0] core_csr_lo_12 ={ core_csr_lo_hi_12 , core_csr_reg_pmp_5_cfg_r }; 
    wire[2:0] core_csr_hi_hi_12 ={ core_csr_reg_pmp_5_cfg_l , core_csr_reg_pmp_5_cfg_res }; 
    wire[4:0] core_csr_hi_12 ={ core_csr_hi_hi_12 , core_csr_reg_pmp_5_cfg_a }; 
    wire[1:0] core_csr_lo_hi_13 ={ core_csr_reg_pmp_6_cfg_x , core_csr_reg_pmp_6_cfg_w }; 
    wire[2:0] core_csr_lo_13 ={ core_csr_lo_hi_13 , core_csr_reg_pmp_6_cfg_r }; 
    wire[2:0] core_csr_hi_hi_13 ={ core_csr_reg_pmp_6_cfg_l , core_csr_reg_pmp_6_cfg_res }; 
    wire[4:0] core_csr_hi_13 ={ core_csr_hi_hi_13 , core_csr_reg_pmp_6_cfg_a }; 
    wire[1:0] core_csr_lo_hi_14 ={ core_csr_reg_pmp_7_cfg_x , core_csr_reg_pmp_7_cfg_w }; 
    wire[2:0] core_csr_lo_14 ={ core_csr_lo_hi_14 , core_csr_reg_pmp_7_cfg_r }; 
    wire[2:0] core_csr_hi_hi_14 ={ core_csr_reg_pmp_7_cfg_l , core_csr_reg_pmp_7_cfg_res }; 
    wire[4:0] core_csr_hi_14 ={ core_csr_hi_hi_14 , core_csr_reg_pmp_7_cfg_a }; 
    wire[15:0] core_csr_lo_lo_6 ={{ core_csr_hi_8 , core_csr_lo_8 },{ core_csr_hi_7 , core_csr_lo_7 }}; 
    wire[15:0] core_csr_lo_hi_15 ={{ core_csr_hi_10 , core_csr_lo_10 },{ core_csr_hi_9 , core_csr_lo_9 }}; 
    wire[31:0] core_csr_lo_15 ={ core_csr_lo_hi_15 , core_csr_lo_lo_6 }; 
    wire[15:0] core_csr_hi_lo_6 ={{ core_csr_hi_12 , core_csr_lo_12 },{ core_csr_hi_11 , core_csr_lo_11 }}; 
    wire[15:0] core_csr_hi_hi_15 ={{ core_csr_hi_14 , core_csr_lo_14 },{ core_csr_hi_13 , core_csr_lo_13 }}; 
    wire[31:0] core_csr_hi_15 ={ core_csr_hi_hi_15 , core_csr_hi_lo_6 }; 
    wire[1:0] core_csr_lo_hi_16 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_16 ={ core_csr_lo_hi_16 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_16 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_16 ={ core_csr_hi_hi_16 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_17 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_17 ={ core_csr_lo_hi_17 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_17 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_17 ={ core_csr_hi_hi_17 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_18 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_18 ={ core_csr_lo_hi_18 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_18 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_18 ={ core_csr_hi_hi_18 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_19 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_19 ={ core_csr_lo_hi_19 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_19 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_19 ={ core_csr_hi_hi_19 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_20 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_20 ={ core_csr_lo_hi_20 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_20 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_20 ={ core_csr_hi_hi_20 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_21 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_21 ={ core_csr_lo_hi_21 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_21 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_21 ={ core_csr_hi_hi_21 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_22 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_22 ={ core_csr_lo_hi_22 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_22 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_22 ={ core_csr_hi_hi_22 , core_csr_read_pmp_15_cfg_a }; 
    wire[1:0] core_csr_lo_hi_23 ={ core_csr_read_pmp_15_cfg_x , core_csr_read_pmp_15_cfg_w }; 
    wire[2:0] core_csr_lo_23 ={ core_csr_lo_hi_23 , core_csr_read_pmp_15_cfg_r }; 
    wire[2:0] core_csr_hi_hi_23 ={ core_csr_read_pmp_15_cfg_l , core_csr_read_pmp_15_cfg_res }; 
    wire[4:0] core_csr_hi_23 ={ core_csr_hi_hi_23 , core_csr_read_pmp_15_cfg_a }; 
    wire[15:0] core_csr_lo_lo_7 ={{ core_csr_hi_17 , core_csr_lo_17 },{ core_csr_hi_16 , core_csr_lo_16 }}; 
    wire[15:0] core_csr_lo_hi_24 ={{ core_csr_hi_19 , core_csr_lo_19 },{ core_csr_hi_18 , core_csr_lo_18 }}; 
    wire[31:0] core_csr_lo_24 ={ core_csr_lo_hi_24 , core_csr_lo_lo_7 }; 
    wire[15:0] core_csr_hi_lo_7 ={{ core_csr_hi_21 , core_csr_lo_21 },{ core_csr_hi_20 , core_csr_lo_20 }}; 
    wire[15:0] core_csr_hi_hi_24 ={{ core_csr_hi_23 , core_csr_lo_23 },{ core_csr_hi_22 , core_csr_lo_22 }}; 
    wire[31:0] core_csr_hi_24 ={ core_csr_hi_hi_24 , core_csr_hi_lo_7 }; reg[63:0] core_csr_reg_custom_0 ; 
    wire core_csr_reg_custom_read =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'h7C1; reg[63:0] core_csr_reg_custom_1 ; 
    wire core_csr_reg_custom_read_1 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF12; reg[63:0] core_csr_reg_custom_2 ; 
    wire core_csr_reg_custom_read_2 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF11; reg[63:0] core_csr_reg_custom_3 ; 
    wire core_csr_reg_custom_read_3 =(| core_csr_io_rw_cmd )& core_csr_io_rw_addr ==12'hF13; 
    wire core_csr__io_rw_stall_output = core_csr_reg_custom_read_3 & core_csr_io_customCSRs_3_stall  ? 1'h1: core_csr_reg_custom_read_2 & core_csr_io_customCSRs_2_stall  ? 1'h1: core_csr_reg_custom_read_1 & core_csr_io_customCSRs_1_stall  ? 1'h1: core_csr_reg_custom_read & core_csr_io_customCSRs_0_stall ; 
    wire[12:0] core_csr_addr ={ core_csr__io_status_v_output , core_csr_io_rw_addr }; 
    wire[11:0] core_csr_decoded_decoded_plaInput ; 
    wire[11:0] core_csr_decoded_decoded_invInputs =~ core_csr_decoded_decoded_plaInput ; 
    wire[131:0] core_csr_decoded_decoded_invMatrixOutputs ; 
    wire core_csr_decoded_decoded_andMatrixInput_0 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi ={ core_csr_decoded_decoded_andMatrixInput_9 , core_csr_decoded_decoded_andMatrixInput_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo ={ core_csr_decoded_decoded_lo_lo_hi , core_csr_decoded_decoded_andMatrixInput_11 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi ={ core_csr_decoded_decoded_andMatrixInput_6 , core_csr_decoded_decoded_andMatrixInput_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi ={ core_csr_decoded_decoded_lo_hi_hi , core_csr_decoded_decoded_andMatrixInput_8 }; 
    wire[5:0] core_csr_decoded_decoded_lo ={ core_csr_decoded_decoded_lo_hi , core_csr_decoded_decoded_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi ={ core_csr_decoded_decoded_andMatrixInput_3 , core_csr_decoded_decoded_andMatrixInput_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo ={ core_csr_decoded_decoded_hi_lo_hi , core_csr_decoded_decoded_andMatrixInput_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi ={ core_csr_decoded_decoded_andMatrixInput_0 , core_csr_decoded_decoded_andMatrixInput_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi ={ core_csr_decoded_decoded_hi_hi_hi , core_csr_decoded_decoded_andMatrixInput_2 }; 
    wire[5:0] core_csr_decoded_decoded_hi ={ core_csr_decoded_decoded_hi_hi , core_csr_decoded_decoded_hi_lo }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_1 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_1 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_1 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_1 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_1 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_1 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_1 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_1 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_1 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_1 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_1 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_1 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_9_1 , core_csr_decoded_decoded_andMatrixInput_10_1 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_1 ={ core_csr_decoded_decoded_lo_lo_hi_1 , core_csr_decoded_decoded_andMatrixInput_11_1 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_6_1 , core_csr_decoded_decoded_andMatrixInput_7_1 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_1 ={ core_csr_decoded_decoded_lo_hi_hi_1 , core_csr_decoded_decoded_andMatrixInput_8_1 }; 
    wire[5:0] core_csr_decoded_decoded_lo_1 ={ core_csr_decoded_decoded_lo_hi_1 , core_csr_decoded_decoded_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_3_1 , core_csr_decoded_decoded_andMatrixInput_4_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_1 ={ core_csr_decoded_decoded_hi_lo_hi_1 , core_csr_decoded_decoded_andMatrixInput_5_1 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_1 ={ core_csr_decoded_decoded_andMatrixInput_0_1 , core_csr_decoded_decoded_andMatrixInput_1_1 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_1 ={ core_csr_decoded_decoded_hi_hi_hi_1 , core_csr_decoded_decoded_andMatrixInput_2_1 }; 
    wire[5:0] core_csr_decoded_decoded_hi_1 ={ core_csr_decoded_decoded_hi_hi_1 , core_csr_decoded_decoded_hi_lo_1 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_2 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_2 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_2 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_2 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_2 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_2 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_2 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_2 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_2 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_2 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_2 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_2 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_9_2 , core_csr_decoded_decoded_andMatrixInput_10_2 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_2 ={ core_csr_decoded_decoded_lo_lo_hi_2 , core_csr_decoded_decoded_andMatrixInput_11_2 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_6_2 , core_csr_decoded_decoded_andMatrixInput_7_2 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_2 ={ core_csr_decoded_decoded_lo_hi_hi_2 , core_csr_decoded_decoded_andMatrixInput_8_2 }; 
    wire[5:0] core_csr_decoded_decoded_lo_2 ={ core_csr_decoded_decoded_lo_hi_2 , core_csr_decoded_decoded_lo_lo_2 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_3_2 , core_csr_decoded_decoded_andMatrixInput_4_2 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_2 ={ core_csr_decoded_decoded_hi_lo_hi_2 , core_csr_decoded_decoded_andMatrixInput_5_2 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_2 ={ core_csr_decoded_decoded_andMatrixInput_0_2 , core_csr_decoded_decoded_andMatrixInput_1_2 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_2 ={ core_csr_decoded_decoded_hi_hi_hi_2 , core_csr_decoded_decoded_andMatrixInput_2_2 }; 
    wire[5:0] core_csr_decoded_decoded_hi_2 ={ core_csr_decoded_decoded_hi_hi_2 , core_csr_decoded_decoded_hi_lo_2 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_3 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_3 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_3 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_3 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_3 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_3 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_3 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_3 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_3 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_3 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_3 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_3 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_9_3 , core_csr_decoded_decoded_andMatrixInput_10_3 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_3 ={ core_csr_decoded_decoded_lo_lo_hi_3 , core_csr_decoded_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_6_3 , core_csr_decoded_decoded_andMatrixInput_7_3 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_3 ={ core_csr_decoded_decoded_lo_hi_hi_3 , core_csr_decoded_decoded_andMatrixInput_8_3 }; 
    wire[5:0] core_csr_decoded_decoded_lo_3 ={ core_csr_decoded_decoded_lo_hi_3 , core_csr_decoded_decoded_lo_lo_3 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_3_3 , core_csr_decoded_decoded_andMatrixInput_4_3 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_3 ={ core_csr_decoded_decoded_hi_lo_hi_3 , core_csr_decoded_decoded_andMatrixInput_5_3 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_3 ={ core_csr_decoded_decoded_andMatrixInput_0_3 , core_csr_decoded_decoded_andMatrixInput_1_3 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_3 ={ core_csr_decoded_decoded_hi_hi_hi_3 , core_csr_decoded_decoded_andMatrixInput_2_3 }; 
    wire[5:0] core_csr_decoded_decoded_hi_3 ={ core_csr_decoded_decoded_hi_hi_3 , core_csr_decoded_decoded_hi_lo_3 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_4 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_4 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_4 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_4 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_4 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_4 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_4 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_4 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_4 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_4 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_4 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_4 ={ core_csr_decoded_decoded_andMatrixInput_9_4 , core_csr_decoded_decoded_andMatrixInput_10_4 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_6_4 , core_csr_decoded_decoded_andMatrixInput_7_4 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_4 ={ core_csr_decoded_decoded_lo_hi_hi_4 , core_csr_decoded_decoded_andMatrixInput_8_4 }; 
    wire[4:0] core_csr_decoded_decoded_lo_4 ={ core_csr_decoded_decoded_lo_hi_4 , core_csr_decoded_decoded_lo_lo_4 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_3_4 , core_csr_decoded_decoded_andMatrixInput_4_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_4 ={ core_csr_decoded_decoded_hi_lo_hi_4 , core_csr_decoded_decoded_andMatrixInput_5_4 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_0_4 , core_csr_decoded_decoded_andMatrixInput_1_4 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_4 ={ core_csr_decoded_decoded_hi_hi_hi_4 , core_csr_decoded_decoded_andMatrixInput_2_4 }; 
    wire[5:0] core_csr_decoded_decoded_hi_4 ={ core_csr_decoded_decoded_hi_hi_4 , core_csr_decoded_decoded_hi_lo_4 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_5 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_5 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_5 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_5 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_5 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_5 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_5 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_5 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_5 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_5 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_5 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_5 ={ core_csr_decoded_decoded_andMatrixInput_9_5 , core_csr_decoded_decoded_andMatrixInput_10_5 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_6_5 , core_csr_decoded_decoded_andMatrixInput_7_5 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_5 ={ core_csr_decoded_decoded_lo_hi_hi_5 , core_csr_decoded_decoded_andMatrixInput_8_5 }; 
    wire[4:0] core_csr_decoded_decoded_lo_5 ={ core_csr_decoded_decoded_lo_hi_5 , core_csr_decoded_decoded_lo_lo_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_3_5 , core_csr_decoded_decoded_andMatrixInput_4_5 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_5 ={ core_csr_decoded_decoded_hi_lo_hi_5 , core_csr_decoded_decoded_andMatrixInput_5_5 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_0_5 , core_csr_decoded_decoded_andMatrixInput_1_5 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_5 ={ core_csr_decoded_decoded_hi_hi_hi_5 , core_csr_decoded_decoded_andMatrixInput_2_5 }; 
    wire[5:0] core_csr_decoded_decoded_hi_5 ={ core_csr_decoded_decoded_hi_hi_5 , core_csr_decoded_decoded_hi_lo_5 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_6 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_6 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_6 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_6 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_6 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_6 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_6 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_6 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_6 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_6 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_6 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_4 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_4 ={ core_csr_decoded_decoded_andMatrixInput_9_6 , core_csr_decoded_decoded_andMatrixInput_10_6 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_6 ={ core_csr_decoded_decoded_lo_lo_hi_4 , core_csr_decoded_decoded_andMatrixInput_11_4 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_6_6 , core_csr_decoded_decoded_andMatrixInput_7_6 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_6 ={ core_csr_decoded_decoded_lo_hi_hi_6 , core_csr_decoded_decoded_andMatrixInput_8_6 }; 
    wire[5:0] core_csr_decoded_decoded_lo_6 ={ core_csr_decoded_decoded_lo_hi_6 , core_csr_decoded_decoded_lo_lo_6 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_3_6 , core_csr_decoded_decoded_andMatrixInput_4_6 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_6 ={ core_csr_decoded_decoded_hi_lo_hi_6 , core_csr_decoded_decoded_andMatrixInput_5_6 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_0_6 , core_csr_decoded_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_6 ={ core_csr_decoded_decoded_hi_hi_hi_6 , core_csr_decoded_decoded_andMatrixInput_2_6 }; 
    wire[5:0] core_csr_decoded_decoded_hi_6 ={ core_csr_decoded_decoded_hi_hi_6 , core_csr_decoded_decoded_hi_lo_6 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_7 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_7 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_7 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_7 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_7 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_7 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_7 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_7 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_7 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_7 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_7 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_5 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_5 ={ core_csr_decoded_decoded_andMatrixInput_9_7 , core_csr_decoded_decoded_andMatrixInput_10_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_7 ={ core_csr_decoded_decoded_lo_lo_hi_5 , core_csr_decoded_decoded_andMatrixInput_11_5 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_6_7 , core_csr_decoded_decoded_andMatrixInput_7_7 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_7 ={ core_csr_decoded_decoded_lo_hi_hi_7 , core_csr_decoded_decoded_andMatrixInput_8_7 }; 
    wire[5:0] core_csr_decoded_decoded_lo_7 ={ core_csr_decoded_decoded_lo_hi_7 , core_csr_decoded_decoded_lo_lo_7 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_3_7 , core_csr_decoded_decoded_andMatrixInput_4_7 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_7 ={ core_csr_decoded_decoded_hi_lo_hi_7 , core_csr_decoded_decoded_andMatrixInput_5_7 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_0_7 , core_csr_decoded_decoded_andMatrixInput_1_7 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_7 ={ core_csr_decoded_decoded_hi_hi_hi_7 , core_csr_decoded_decoded_andMatrixInput_2_7 }; 
    wire[5:0] core_csr_decoded_decoded_hi_7 ={ core_csr_decoded_decoded_hi_hi_7 , core_csr_decoded_decoded_hi_lo_7 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_8 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_8 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_8 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_8 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_8 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_8 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_8 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_8 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_8 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_8 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_8 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_6 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_6 ={ core_csr_decoded_decoded_andMatrixInput_9_8 , core_csr_decoded_decoded_andMatrixInput_10_8 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_8 ={ core_csr_decoded_decoded_lo_lo_hi_6 , core_csr_decoded_decoded_andMatrixInput_11_6 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_6_8 , core_csr_decoded_decoded_andMatrixInput_7_8 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_8 ={ core_csr_decoded_decoded_lo_hi_hi_8 , core_csr_decoded_decoded_andMatrixInput_8_8 }; 
    wire[5:0] core_csr_decoded_decoded_lo_8 ={ core_csr_decoded_decoded_lo_hi_8 , core_csr_decoded_decoded_lo_lo_8 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_3_8 , core_csr_decoded_decoded_andMatrixInput_4_8 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_8 ={ core_csr_decoded_decoded_hi_lo_hi_8 , core_csr_decoded_decoded_andMatrixInput_5_8 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_0_8 , core_csr_decoded_decoded_andMatrixInput_1_8 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_8 ={ core_csr_decoded_decoded_hi_hi_hi_8 , core_csr_decoded_decoded_andMatrixInput_2_8 }; 
    wire[5:0] core_csr_decoded_decoded_hi_8 ={ core_csr_decoded_decoded_hi_hi_8 , core_csr_decoded_decoded_hi_lo_8 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_9 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_9 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_9 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_9 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_9 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_9 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_9 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_9 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_9 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_9 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_9 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_7 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_7 ={ core_csr_decoded_decoded_andMatrixInput_9_9 , core_csr_decoded_decoded_andMatrixInput_10_9 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_9 ={ core_csr_decoded_decoded_lo_lo_hi_7 , core_csr_decoded_decoded_andMatrixInput_11_7 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_6_9 , core_csr_decoded_decoded_andMatrixInput_7_9 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_9 ={ core_csr_decoded_decoded_lo_hi_hi_9 , core_csr_decoded_decoded_andMatrixInput_8_9 }; 
    wire[5:0] core_csr_decoded_decoded_lo_9 ={ core_csr_decoded_decoded_lo_hi_9 , core_csr_decoded_decoded_lo_lo_9 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_3_9 , core_csr_decoded_decoded_andMatrixInput_4_9 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_9 ={ core_csr_decoded_decoded_hi_lo_hi_9 , core_csr_decoded_decoded_andMatrixInput_5_9 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_0_9 , core_csr_decoded_decoded_andMatrixInput_1_9 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_9 ={ core_csr_decoded_decoded_hi_hi_hi_9 , core_csr_decoded_decoded_andMatrixInput_2_9 }; 
    wire[5:0] core_csr_decoded_decoded_hi_9 ={ core_csr_decoded_decoded_hi_hi_9 , core_csr_decoded_decoded_hi_lo_9 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_10 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_10 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_10 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_10 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_10 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_10 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_10 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_10 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_10 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_10 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_10 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_8 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_8 ={ core_csr_decoded_decoded_andMatrixInput_9_10 , core_csr_decoded_decoded_andMatrixInput_10_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_10 ={ core_csr_decoded_decoded_lo_lo_hi_8 , core_csr_decoded_decoded_andMatrixInput_11_8 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_6_10 , core_csr_decoded_decoded_andMatrixInput_7_10 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_10 ={ core_csr_decoded_decoded_lo_hi_hi_10 , core_csr_decoded_decoded_andMatrixInput_8_10 }; 
    wire[5:0] core_csr_decoded_decoded_lo_10 ={ core_csr_decoded_decoded_lo_hi_10 , core_csr_decoded_decoded_lo_lo_10 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_3_10 , core_csr_decoded_decoded_andMatrixInput_4_10 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_10 ={ core_csr_decoded_decoded_hi_lo_hi_10 , core_csr_decoded_decoded_andMatrixInput_5_10 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_0_10 , core_csr_decoded_decoded_andMatrixInput_1_10 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_10 ={ core_csr_decoded_decoded_hi_hi_hi_10 , core_csr_decoded_decoded_andMatrixInput_2_10 }; 
    wire[5:0] core_csr_decoded_decoded_hi_10 ={ core_csr_decoded_decoded_hi_hi_10 , core_csr_decoded_decoded_hi_lo_10 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_11 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_11 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_11 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_11 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_11 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_11 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_11 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_11 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_11 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_11 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_11 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_9 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_9 ={ core_csr_decoded_decoded_andMatrixInput_9_11 , core_csr_decoded_decoded_andMatrixInput_10_11 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_11 ={ core_csr_decoded_decoded_lo_lo_hi_9 , core_csr_decoded_decoded_andMatrixInput_11_9 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_6_11 , core_csr_decoded_decoded_andMatrixInput_7_11 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_11 ={ core_csr_decoded_decoded_lo_hi_hi_11 , core_csr_decoded_decoded_andMatrixInput_8_11 }; 
    wire[5:0] core_csr_decoded_decoded_lo_11 ={ core_csr_decoded_decoded_lo_hi_11 , core_csr_decoded_decoded_lo_lo_11 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_3_11 , core_csr_decoded_decoded_andMatrixInput_4_11 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_11 ={ core_csr_decoded_decoded_hi_lo_hi_11 , core_csr_decoded_decoded_andMatrixInput_5_11 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_0_11 , core_csr_decoded_decoded_andMatrixInput_1_11 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_11 ={ core_csr_decoded_decoded_hi_hi_hi_11 , core_csr_decoded_decoded_andMatrixInput_2_11 }; 
    wire[5:0] core_csr_decoded_decoded_hi_11 ={ core_csr_decoded_decoded_hi_hi_11 , core_csr_decoded_decoded_hi_lo_11 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_12 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_12 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_12 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_12 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_12 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_12 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_12 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_12 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_12 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_12 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_12 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_10 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_10 ={ core_csr_decoded_decoded_andMatrixInput_9_12 , core_csr_decoded_decoded_andMatrixInput_10_12 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_12 ={ core_csr_decoded_decoded_lo_lo_hi_10 , core_csr_decoded_decoded_andMatrixInput_11_10 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_6_12 , core_csr_decoded_decoded_andMatrixInput_7_12 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_12 ={ core_csr_decoded_decoded_lo_hi_hi_12 , core_csr_decoded_decoded_andMatrixInput_8_12 }; 
    wire[5:0] core_csr_decoded_decoded_lo_12 ={ core_csr_decoded_decoded_lo_hi_12 , core_csr_decoded_decoded_lo_lo_12 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_3_12 , core_csr_decoded_decoded_andMatrixInput_4_12 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_12 ={ core_csr_decoded_decoded_hi_lo_hi_12 , core_csr_decoded_decoded_andMatrixInput_5_12 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_0_12 , core_csr_decoded_decoded_andMatrixInput_1_12 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_12 ={ core_csr_decoded_decoded_hi_hi_hi_12 , core_csr_decoded_decoded_andMatrixInput_2_12 }; 
    wire[5:0] core_csr_decoded_decoded_hi_12 ={ core_csr_decoded_decoded_hi_hi_12 , core_csr_decoded_decoded_hi_lo_12 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_13 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_13 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_13 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_13 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_13 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_13 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_13 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_13 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_13 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_13 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_13 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_11 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_11 ={ core_csr_decoded_decoded_andMatrixInput_9_13 , core_csr_decoded_decoded_andMatrixInput_10_13 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_13 ={ core_csr_decoded_decoded_lo_lo_hi_11 , core_csr_decoded_decoded_andMatrixInput_11_11 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_6_13 , core_csr_decoded_decoded_andMatrixInput_7_13 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_13 ={ core_csr_decoded_decoded_lo_hi_hi_13 , core_csr_decoded_decoded_andMatrixInput_8_13 }; 
    wire[5:0] core_csr_decoded_decoded_lo_13 ={ core_csr_decoded_decoded_lo_hi_13 , core_csr_decoded_decoded_lo_lo_13 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_3_13 , core_csr_decoded_decoded_andMatrixInput_4_13 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_13 ={ core_csr_decoded_decoded_hi_lo_hi_13 , core_csr_decoded_decoded_andMatrixInput_5_13 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_0_13 , core_csr_decoded_decoded_andMatrixInput_1_13 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_13 ={ core_csr_decoded_decoded_hi_hi_hi_13 , core_csr_decoded_decoded_andMatrixInput_2_13 }; 
    wire[5:0] core_csr_decoded_decoded_hi_13 ={ core_csr_decoded_decoded_hi_hi_13 , core_csr_decoded_decoded_hi_lo_13 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_14 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_14 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_14 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_14 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_14 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_14 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_14 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_14 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_14 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_14 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_14 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_12 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_12 ={ core_csr_decoded_decoded_andMatrixInput_9_14 , core_csr_decoded_decoded_andMatrixInput_10_14 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_14 ={ core_csr_decoded_decoded_lo_lo_hi_12 , core_csr_decoded_decoded_andMatrixInput_11_12 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_6_14 , core_csr_decoded_decoded_andMatrixInput_7_14 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_14 ={ core_csr_decoded_decoded_lo_hi_hi_14 , core_csr_decoded_decoded_andMatrixInput_8_14 }; 
    wire[5:0] core_csr_decoded_decoded_lo_14 ={ core_csr_decoded_decoded_lo_hi_14 , core_csr_decoded_decoded_lo_lo_14 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_3_14 , core_csr_decoded_decoded_andMatrixInput_4_14 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_14 ={ core_csr_decoded_decoded_hi_lo_hi_14 , core_csr_decoded_decoded_andMatrixInput_5_14 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_0_14 , core_csr_decoded_decoded_andMatrixInput_1_14 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_14 ={ core_csr_decoded_decoded_hi_hi_hi_14 , core_csr_decoded_decoded_andMatrixInput_2_14 }; 
    wire[5:0] core_csr_decoded_decoded_hi_14 ={ core_csr_decoded_decoded_hi_hi_14 , core_csr_decoded_decoded_hi_lo_14 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_15 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_15 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_15 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_15 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_15 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_15 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_15 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_15 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_15 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_15 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_15 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_13 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_13 ={ core_csr_decoded_decoded_andMatrixInput_9_15 , core_csr_decoded_decoded_andMatrixInput_10_15 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_15 ={ core_csr_decoded_decoded_lo_lo_hi_13 , core_csr_decoded_decoded_andMatrixInput_11_13 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_6_15 , core_csr_decoded_decoded_andMatrixInput_7_15 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_15 ={ core_csr_decoded_decoded_lo_hi_hi_15 , core_csr_decoded_decoded_andMatrixInput_8_15 }; 
    wire[5:0] core_csr_decoded_decoded_lo_15 ={ core_csr_decoded_decoded_lo_hi_15 , core_csr_decoded_decoded_lo_lo_15 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_3_15 , core_csr_decoded_decoded_andMatrixInput_4_15 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_15 ={ core_csr_decoded_decoded_hi_lo_hi_15 , core_csr_decoded_decoded_andMatrixInput_5_15 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_0_15 , core_csr_decoded_decoded_andMatrixInput_1_15 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_15 ={ core_csr_decoded_decoded_hi_hi_hi_15 , core_csr_decoded_decoded_andMatrixInput_2_15 }; 
    wire[5:0] core_csr_decoded_decoded_hi_15 ={ core_csr_decoded_decoded_hi_hi_15 , core_csr_decoded_decoded_hi_lo_15 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_16 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_16 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_16 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_16 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_16 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_16 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_16 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_16 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_16 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_16 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_16 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_14 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_14 ={ core_csr_decoded_decoded_andMatrixInput_9_16 , core_csr_decoded_decoded_andMatrixInput_10_16 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_16 ={ core_csr_decoded_decoded_lo_lo_hi_14 , core_csr_decoded_decoded_andMatrixInput_11_14 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_6_16 , core_csr_decoded_decoded_andMatrixInput_7_16 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_16 ={ core_csr_decoded_decoded_lo_hi_hi_16 , core_csr_decoded_decoded_andMatrixInput_8_16 }; 
    wire[5:0] core_csr_decoded_decoded_lo_16 ={ core_csr_decoded_decoded_lo_hi_16 , core_csr_decoded_decoded_lo_lo_16 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_3_16 , core_csr_decoded_decoded_andMatrixInput_4_16 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_16 ={ core_csr_decoded_decoded_hi_lo_hi_16 , core_csr_decoded_decoded_andMatrixInput_5_16 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_0_16 , core_csr_decoded_decoded_andMatrixInput_1_16 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_16 ={ core_csr_decoded_decoded_hi_hi_hi_16 , core_csr_decoded_decoded_andMatrixInput_2_16 }; 
    wire[5:0] core_csr_decoded_decoded_hi_16 ={ core_csr_decoded_decoded_hi_hi_16 , core_csr_decoded_decoded_hi_lo_16 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_17 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_17 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_17 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_17 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_17 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_17 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_17 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_17 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_17 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_17 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_17 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_15 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_15 ={ core_csr_decoded_decoded_andMatrixInput_9_17 , core_csr_decoded_decoded_andMatrixInput_10_17 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_17 ={ core_csr_decoded_decoded_lo_lo_hi_15 , core_csr_decoded_decoded_andMatrixInput_11_15 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_6_17 , core_csr_decoded_decoded_andMatrixInput_7_17 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_17 ={ core_csr_decoded_decoded_lo_hi_hi_17 , core_csr_decoded_decoded_andMatrixInput_8_17 }; 
    wire[5:0] core_csr_decoded_decoded_lo_17 ={ core_csr_decoded_decoded_lo_hi_17 , core_csr_decoded_decoded_lo_lo_17 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_3_17 , core_csr_decoded_decoded_andMatrixInput_4_17 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_17 ={ core_csr_decoded_decoded_hi_lo_hi_17 , core_csr_decoded_decoded_andMatrixInput_5_17 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_0_17 , core_csr_decoded_decoded_andMatrixInput_1_17 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_17 ={ core_csr_decoded_decoded_hi_hi_hi_17 , core_csr_decoded_decoded_andMatrixInput_2_17 }; 
    wire[5:0] core_csr_decoded_decoded_hi_17 ={ core_csr_decoded_decoded_hi_hi_17 , core_csr_decoded_decoded_hi_lo_17 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_18 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_18 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_18 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_18 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_18 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_18 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_18 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_18 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_18 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_18 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_18 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_16 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_16 ={ core_csr_decoded_decoded_andMatrixInput_9_18 , core_csr_decoded_decoded_andMatrixInput_10_18 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_18 ={ core_csr_decoded_decoded_lo_lo_hi_16 , core_csr_decoded_decoded_andMatrixInput_11_16 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_6_18 , core_csr_decoded_decoded_andMatrixInput_7_18 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_18 ={ core_csr_decoded_decoded_lo_hi_hi_18 , core_csr_decoded_decoded_andMatrixInput_8_18 }; 
    wire[5:0] core_csr_decoded_decoded_lo_18 ={ core_csr_decoded_decoded_lo_hi_18 , core_csr_decoded_decoded_lo_lo_18 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_3_18 , core_csr_decoded_decoded_andMatrixInput_4_18 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_18 ={ core_csr_decoded_decoded_hi_lo_hi_18 , core_csr_decoded_decoded_andMatrixInput_5_18 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_0_18 , core_csr_decoded_decoded_andMatrixInput_1_18 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_18 ={ core_csr_decoded_decoded_hi_hi_hi_18 , core_csr_decoded_decoded_andMatrixInput_2_18 }; 
    wire[5:0] core_csr_decoded_decoded_hi_18 ={ core_csr_decoded_decoded_hi_hi_18 , core_csr_decoded_decoded_hi_lo_18 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_19 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_19 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_19 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_19 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_19 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_19 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_19 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_19 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_19 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_19 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_19 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_17 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_17 ={ core_csr_decoded_decoded_andMatrixInput_9_19 , core_csr_decoded_decoded_andMatrixInput_10_19 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_19 ={ core_csr_decoded_decoded_lo_lo_hi_17 , core_csr_decoded_decoded_andMatrixInput_11_17 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_6_19 , core_csr_decoded_decoded_andMatrixInput_7_19 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_19 ={ core_csr_decoded_decoded_lo_hi_hi_19 , core_csr_decoded_decoded_andMatrixInput_8_19 }; 
    wire[5:0] core_csr_decoded_decoded_lo_19 ={ core_csr_decoded_decoded_lo_hi_19 , core_csr_decoded_decoded_lo_lo_19 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_3_19 , core_csr_decoded_decoded_andMatrixInput_4_19 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_19 ={ core_csr_decoded_decoded_hi_lo_hi_19 , core_csr_decoded_decoded_andMatrixInput_5_19 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_0_19 , core_csr_decoded_decoded_andMatrixInput_1_19 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_19 ={ core_csr_decoded_decoded_hi_hi_hi_19 , core_csr_decoded_decoded_andMatrixInput_2_19 }; 
    wire[5:0] core_csr_decoded_decoded_hi_19 ={ core_csr_decoded_decoded_hi_hi_19 , core_csr_decoded_decoded_hi_lo_19 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_20 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_20 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_20 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_20 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_20 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_20 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_20 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_20 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_20 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_20 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_20 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_18 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_18 ={ core_csr_decoded_decoded_andMatrixInput_9_20 , core_csr_decoded_decoded_andMatrixInput_10_20 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_20 ={ core_csr_decoded_decoded_lo_lo_hi_18 , core_csr_decoded_decoded_andMatrixInput_11_18 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_6_20 , core_csr_decoded_decoded_andMatrixInput_7_20 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_20 ={ core_csr_decoded_decoded_lo_hi_hi_20 , core_csr_decoded_decoded_andMatrixInput_8_20 }; 
    wire[5:0] core_csr_decoded_decoded_lo_20 ={ core_csr_decoded_decoded_lo_hi_20 , core_csr_decoded_decoded_lo_lo_20 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_3_20 , core_csr_decoded_decoded_andMatrixInput_4_20 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_20 ={ core_csr_decoded_decoded_hi_lo_hi_20 , core_csr_decoded_decoded_andMatrixInput_5_20 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_0_20 , core_csr_decoded_decoded_andMatrixInput_1_20 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_20 ={ core_csr_decoded_decoded_hi_hi_hi_20 , core_csr_decoded_decoded_andMatrixInput_2_20 }; 
    wire[5:0] core_csr_decoded_decoded_hi_20 ={ core_csr_decoded_decoded_hi_hi_20 , core_csr_decoded_decoded_hi_lo_20 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_21 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_21 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_21 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_21 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_21 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_21 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_21 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_21 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_21 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_21 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_21 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_19 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_19 ={ core_csr_decoded_decoded_andMatrixInput_9_21 , core_csr_decoded_decoded_andMatrixInput_10_21 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_21 ={ core_csr_decoded_decoded_lo_lo_hi_19 , core_csr_decoded_decoded_andMatrixInput_11_19 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_6_21 , core_csr_decoded_decoded_andMatrixInput_7_21 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_21 ={ core_csr_decoded_decoded_lo_hi_hi_21 , core_csr_decoded_decoded_andMatrixInput_8_21 }; 
    wire[5:0] core_csr_decoded_decoded_lo_21 ={ core_csr_decoded_decoded_lo_hi_21 , core_csr_decoded_decoded_lo_lo_21 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_3_21 , core_csr_decoded_decoded_andMatrixInput_4_21 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_21 ={ core_csr_decoded_decoded_hi_lo_hi_21 , core_csr_decoded_decoded_andMatrixInput_5_21 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_0_21 , core_csr_decoded_decoded_andMatrixInput_1_21 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_21 ={ core_csr_decoded_decoded_hi_hi_hi_21 , core_csr_decoded_decoded_andMatrixInput_2_21 }; 
    wire[5:0] core_csr_decoded_decoded_hi_21 ={ core_csr_decoded_decoded_hi_hi_21 , core_csr_decoded_decoded_hi_lo_21 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_22 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_22 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_22 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_22 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_22 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_22 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_22 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_22 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_22 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_22 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_22 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_20 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_20 ={ core_csr_decoded_decoded_andMatrixInput_9_22 , core_csr_decoded_decoded_andMatrixInput_10_22 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_22 ={ core_csr_decoded_decoded_lo_lo_hi_20 , core_csr_decoded_decoded_andMatrixInput_11_20 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_6_22 , core_csr_decoded_decoded_andMatrixInput_7_22 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_22 ={ core_csr_decoded_decoded_lo_hi_hi_22 , core_csr_decoded_decoded_andMatrixInput_8_22 }; 
    wire[5:0] core_csr_decoded_decoded_lo_22 ={ core_csr_decoded_decoded_lo_hi_22 , core_csr_decoded_decoded_lo_lo_22 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_3_22 , core_csr_decoded_decoded_andMatrixInput_4_22 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_22 ={ core_csr_decoded_decoded_hi_lo_hi_22 , core_csr_decoded_decoded_andMatrixInput_5_22 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_0_22 , core_csr_decoded_decoded_andMatrixInput_1_22 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_22 ={ core_csr_decoded_decoded_hi_hi_hi_22 , core_csr_decoded_decoded_andMatrixInput_2_22 }; 
    wire[5:0] core_csr_decoded_decoded_hi_22 ={ core_csr_decoded_decoded_hi_hi_22 , core_csr_decoded_decoded_hi_lo_22 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_23 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_23 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_23 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_23 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_23 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_23 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_23 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_23 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_23 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_23 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_23 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_21 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_21 ={ core_csr_decoded_decoded_andMatrixInput_9_23 , core_csr_decoded_decoded_andMatrixInput_10_23 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_23 ={ core_csr_decoded_decoded_lo_lo_hi_21 , core_csr_decoded_decoded_andMatrixInput_11_21 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_6_23 , core_csr_decoded_decoded_andMatrixInput_7_23 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_23 ={ core_csr_decoded_decoded_lo_hi_hi_23 , core_csr_decoded_decoded_andMatrixInput_8_23 }; 
    wire[5:0] core_csr_decoded_decoded_lo_23 ={ core_csr_decoded_decoded_lo_hi_23 , core_csr_decoded_decoded_lo_lo_23 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_3_23 , core_csr_decoded_decoded_andMatrixInput_4_23 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_23 ={ core_csr_decoded_decoded_hi_lo_hi_23 , core_csr_decoded_decoded_andMatrixInput_5_23 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_0_23 , core_csr_decoded_decoded_andMatrixInput_1_23 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_23 ={ core_csr_decoded_decoded_hi_hi_hi_23 , core_csr_decoded_decoded_andMatrixInput_2_23 }; 
    wire[5:0] core_csr_decoded_decoded_hi_23 ={ core_csr_decoded_decoded_hi_hi_23 , core_csr_decoded_decoded_hi_lo_23 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_24 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_24 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_24 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_24 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_24 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_24 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_24 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_24 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_24 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_24 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_24 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_22 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_22 ={ core_csr_decoded_decoded_andMatrixInput_9_24 , core_csr_decoded_decoded_andMatrixInput_10_24 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_24 ={ core_csr_decoded_decoded_lo_lo_hi_22 , core_csr_decoded_decoded_andMatrixInput_11_22 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_6_24 , core_csr_decoded_decoded_andMatrixInput_7_24 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_24 ={ core_csr_decoded_decoded_lo_hi_hi_24 , core_csr_decoded_decoded_andMatrixInput_8_24 }; 
    wire[5:0] core_csr_decoded_decoded_lo_24 ={ core_csr_decoded_decoded_lo_hi_24 , core_csr_decoded_decoded_lo_lo_24 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_3_24 , core_csr_decoded_decoded_andMatrixInput_4_24 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_24 ={ core_csr_decoded_decoded_hi_lo_hi_24 , core_csr_decoded_decoded_andMatrixInput_5_24 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_0_24 , core_csr_decoded_decoded_andMatrixInput_1_24 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_24 ={ core_csr_decoded_decoded_hi_hi_hi_24 , core_csr_decoded_decoded_andMatrixInput_2_24 }; 
    wire[5:0] core_csr_decoded_decoded_hi_24 ={ core_csr_decoded_decoded_hi_hi_24 , core_csr_decoded_decoded_hi_lo_24 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_25 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_25 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_25 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_25 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_25 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_25 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_25 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_25 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_25 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_25 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_25 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_23 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_23 ={ core_csr_decoded_decoded_andMatrixInput_9_25 , core_csr_decoded_decoded_andMatrixInput_10_25 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_25 ={ core_csr_decoded_decoded_lo_lo_hi_23 , core_csr_decoded_decoded_andMatrixInput_11_23 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_6_25 , core_csr_decoded_decoded_andMatrixInput_7_25 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_25 ={ core_csr_decoded_decoded_lo_hi_hi_25 , core_csr_decoded_decoded_andMatrixInput_8_25 }; 
    wire[5:0] core_csr_decoded_decoded_lo_25 ={ core_csr_decoded_decoded_lo_hi_25 , core_csr_decoded_decoded_lo_lo_25 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_3_25 , core_csr_decoded_decoded_andMatrixInput_4_25 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_25 ={ core_csr_decoded_decoded_hi_lo_hi_25 , core_csr_decoded_decoded_andMatrixInput_5_25 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_0_25 , core_csr_decoded_decoded_andMatrixInput_1_25 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_25 ={ core_csr_decoded_decoded_hi_hi_hi_25 , core_csr_decoded_decoded_andMatrixInput_2_25 }; 
    wire[5:0] core_csr_decoded_decoded_hi_25 ={ core_csr_decoded_decoded_hi_hi_25 , core_csr_decoded_decoded_hi_lo_25 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_26 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_26 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_26 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_26 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_26 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_26 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_26 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_26 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_26 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_26 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_26 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_24 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_24 ={ core_csr_decoded_decoded_andMatrixInput_9_26 , core_csr_decoded_decoded_andMatrixInput_10_26 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_26 ={ core_csr_decoded_decoded_lo_lo_hi_24 , core_csr_decoded_decoded_andMatrixInput_11_24 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_6_26 , core_csr_decoded_decoded_andMatrixInput_7_26 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_26 ={ core_csr_decoded_decoded_lo_hi_hi_26 , core_csr_decoded_decoded_andMatrixInput_8_26 }; 
    wire[5:0] core_csr_decoded_decoded_lo_26 ={ core_csr_decoded_decoded_lo_hi_26 , core_csr_decoded_decoded_lo_lo_26 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_3_26 , core_csr_decoded_decoded_andMatrixInput_4_26 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_26 ={ core_csr_decoded_decoded_hi_lo_hi_26 , core_csr_decoded_decoded_andMatrixInput_5_26 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_0_26 , core_csr_decoded_decoded_andMatrixInput_1_26 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_26 ={ core_csr_decoded_decoded_hi_hi_hi_26 , core_csr_decoded_decoded_andMatrixInput_2_26 }; 
    wire[5:0] core_csr_decoded_decoded_hi_26 ={ core_csr_decoded_decoded_hi_hi_26 , core_csr_decoded_decoded_hi_lo_26 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_27 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_27 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_27 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_27 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_27 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_27 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_27 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_27 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_27 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_27 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_27 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_25 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_25 ={ core_csr_decoded_decoded_andMatrixInput_9_27 , core_csr_decoded_decoded_andMatrixInput_10_27 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_27 ={ core_csr_decoded_decoded_lo_lo_hi_25 , core_csr_decoded_decoded_andMatrixInput_11_25 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_6_27 , core_csr_decoded_decoded_andMatrixInput_7_27 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_27 ={ core_csr_decoded_decoded_lo_hi_hi_27 , core_csr_decoded_decoded_andMatrixInput_8_27 }; 
    wire[5:0] core_csr_decoded_decoded_lo_27 ={ core_csr_decoded_decoded_lo_hi_27 , core_csr_decoded_decoded_lo_lo_27 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_3_27 , core_csr_decoded_decoded_andMatrixInput_4_27 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_27 ={ core_csr_decoded_decoded_hi_lo_hi_27 , core_csr_decoded_decoded_andMatrixInput_5_27 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_0_27 , core_csr_decoded_decoded_andMatrixInput_1_27 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_27 ={ core_csr_decoded_decoded_hi_hi_hi_27 , core_csr_decoded_decoded_andMatrixInput_2_27 }; 
    wire[5:0] core_csr_decoded_decoded_hi_27 ={ core_csr_decoded_decoded_hi_hi_27 , core_csr_decoded_decoded_hi_lo_27 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_28 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_28 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_28 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_28 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_28 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_28 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_28 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_28 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_28 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_28 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_28 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_26 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_26 ={ core_csr_decoded_decoded_andMatrixInput_9_28 , core_csr_decoded_decoded_andMatrixInput_10_28 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_28 ={ core_csr_decoded_decoded_lo_lo_hi_26 , core_csr_decoded_decoded_andMatrixInput_11_26 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_6_28 , core_csr_decoded_decoded_andMatrixInput_7_28 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_28 ={ core_csr_decoded_decoded_lo_hi_hi_28 , core_csr_decoded_decoded_andMatrixInput_8_28 }; 
    wire[5:0] core_csr_decoded_decoded_lo_28 ={ core_csr_decoded_decoded_lo_hi_28 , core_csr_decoded_decoded_lo_lo_28 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_3_28 , core_csr_decoded_decoded_andMatrixInput_4_28 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_28 ={ core_csr_decoded_decoded_hi_lo_hi_28 , core_csr_decoded_decoded_andMatrixInput_5_28 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_0_28 , core_csr_decoded_decoded_andMatrixInput_1_28 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_28 ={ core_csr_decoded_decoded_hi_hi_hi_28 , core_csr_decoded_decoded_andMatrixInput_2_28 }; 
    wire[5:0] core_csr_decoded_decoded_hi_28 ={ core_csr_decoded_decoded_hi_hi_28 , core_csr_decoded_decoded_hi_lo_28 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_29 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_29 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_29 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_29 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_29 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_29 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_29 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_29 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_29 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_29 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_29 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_27 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_27 ={ core_csr_decoded_decoded_andMatrixInput_9_29 , core_csr_decoded_decoded_andMatrixInput_10_29 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_29 ={ core_csr_decoded_decoded_lo_lo_hi_27 , core_csr_decoded_decoded_andMatrixInput_11_27 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_6_29 , core_csr_decoded_decoded_andMatrixInput_7_29 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_29 ={ core_csr_decoded_decoded_lo_hi_hi_29 , core_csr_decoded_decoded_andMatrixInput_8_29 }; 
    wire[5:0] core_csr_decoded_decoded_lo_29 ={ core_csr_decoded_decoded_lo_hi_29 , core_csr_decoded_decoded_lo_lo_29 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_3_29 , core_csr_decoded_decoded_andMatrixInput_4_29 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_29 ={ core_csr_decoded_decoded_hi_lo_hi_29 , core_csr_decoded_decoded_andMatrixInput_5_29 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_0_29 , core_csr_decoded_decoded_andMatrixInput_1_29 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_29 ={ core_csr_decoded_decoded_hi_hi_hi_29 , core_csr_decoded_decoded_andMatrixInput_2_29 }; 
    wire[5:0] core_csr_decoded_decoded_hi_29 ={ core_csr_decoded_decoded_hi_hi_29 , core_csr_decoded_decoded_hi_lo_29 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_30 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_30 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_30 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_30 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_30 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_30 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_30 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_30 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_30 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_30 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_30 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_28 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_28 ={ core_csr_decoded_decoded_andMatrixInput_9_30 , core_csr_decoded_decoded_andMatrixInput_10_30 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_30 ={ core_csr_decoded_decoded_lo_lo_hi_28 , core_csr_decoded_decoded_andMatrixInput_11_28 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_6_30 , core_csr_decoded_decoded_andMatrixInput_7_30 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_30 ={ core_csr_decoded_decoded_lo_hi_hi_30 , core_csr_decoded_decoded_andMatrixInput_8_30 }; 
    wire[5:0] core_csr_decoded_decoded_lo_30 ={ core_csr_decoded_decoded_lo_hi_30 , core_csr_decoded_decoded_lo_lo_30 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_3_30 , core_csr_decoded_decoded_andMatrixInput_4_30 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_30 ={ core_csr_decoded_decoded_hi_lo_hi_30 , core_csr_decoded_decoded_andMatrixInput_5_30 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_0_30 , core_csr_decoded_decoded_andMatrixInput_1_30 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_30 ={ core_csr_decoded_decoded_hi_hi_hi_30 , core_csr_decoded_decoded_andMatrixInput_2_30 }; 
    wire[5:0] core_csr_decoded_decoded_hi_30 ={ core_csr_decoded_decoded_hi_hi_30 , core_csr_decoded_decoded_hi_lo_30 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_31 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_31 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_31 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_31 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_31 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_31 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_31 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_31 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_31 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_31 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_31 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_29 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_29 ={ core_csr_decoded_decoded_andMatrixInput_9_31 , core_csr_decoded_decoded_andMatrixInput_10_31 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_31 ={ core_csr_decoded_decoded_lo_lo_hi_29 , core_csr_decoded_decoded_andMatrixInput_11_29 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_6_31 , core_csr_decoded_decoded_andMatrixInput_7_31 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_31 ={ core_csr_decoded_decoded_lo_hi_hi_31 , core_csr_decoded_decoded_andMatrixInput_8_31 }; 
    wire[5:0] core_csr_decoded_decoded_lo_31 ={ core_csr_decoded_decoded_lo_hi_31 , core_csr_decoded_decoded_lo_lo_31 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_3_31 , core_csr_decoded_decoded_andMatrixInput_4_31 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_31 ={ core_csr_decoded_decoded_hi_lo_hi_31 , core_csr_decoded_decoded_andMatrixInput_5_31 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_0_31 , core_csr_decoded_decoded_andMatrixInput_1_31 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_31 ={ core_csr_decoded_decoded_hi_hi_hi_31 , core_csr_decoded_decoded_andMatrixInput_2_31 }; 
    wire[5:0] core_csr_decoded_decoded_hi_31 ={ core_csr_decoded_decoded_hi_hi_31 , core_csr_decoded_decoded_hi_lo_31 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_32 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_32 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_32 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_32 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_32 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_32 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_32 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_32 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_32 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_32 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_32 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_30 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_30 ={ core_csr_decoded_decoded_andMatrixInput_9_32 , core_csr_decoded_decoded_andMatrixInput_10_32 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_32 ={ core_csr_decoded_decoded_lo_lo_hi_30 , core_csr_decoded_decoded_andMatrixInput_11_30 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_6_32 , core_csr_decoded_decoded_andMatrixInput_7_32 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_32 ={ core_csr_decoded_decoded_lo_hi_hi_32 , core_csr_decoded_decoded_andMatrixInput_8_32 }; 
    wire[5:0] core_csr_decoded_decoded_lo_32 ={ core_csr_decoded_decoded_lo_hi_32 , core_csr_decoded_decoded_lo_lo_32 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_3_32 , core_csr_decoded_decoded_andMatrixInput_4_32 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_32 ={ core_csr_decoded_decoded_hi_lo_hi_32 , core_csr_decoded_decoded_andMatrixInput_5_32 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_0_32 , core_csr_decoded_decoded_andMatrixInput_1_32 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_32 ={ core_csr_decoded_decoded_hi_hi_hi_32 , core_csr_decoded_decoded_andMatrixInput_2_32 }; 
    wire[5:0] core_csr_decoded_decoded_hi_32 ={ core_csr_decoded_decoded_hi_hi_32 , core_csr_decoded_decoded_hi_lo_32 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_33 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_33 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_33 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_33 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_33 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_33 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_33 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_33 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_33 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_33 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_33 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_31 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_31 ={ core_csr_decoded_decoded_andMatrixInput_9_33 , core_csr_decoded_decoded_andMatrixInput_10_33 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_33 ={ core_csr_decoded_decoded_lo_lo_hi_31 , core_csr_decoded_decoded_andMatrixInput_11_31 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_6_33 , core_csr_decoded_decoded_andMatrixInput_7_33 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_33 ={ core_csr_decoded_decoded_lo_hi_hi_33 , core_csr_decoded_decoded_andMatrixInput_8_33 }; 
    wire[5:0] core_csr_decoded_decoded_lo_33 ={ core_csr_decoded_decoded_lo_hi_33 , core_csr_decoded_decoded_lo_lo_33 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_3_33 , core_csr_decoded_decoded_andMatrixInput_4_33 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_33 ={ core_csr_decoded_decoded_hi_lo_hi_33 , core_csr_decoded_decoded_andMatrixInput_5_33 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_0_33 , core_csr_decoded_decoded_andMatrixInput_1_33 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_33 ={ core_csr_decoded_decoded_hi_hi_hi_33 , core_csr_decoded_decoded_andMatrixInput_2_33 }; 
    wire[5:0] core_csr_decoded_decoded_hi_33 ={ core_csr_decoded_decoded_hi_hi_33 , core_csr_decoded_decoded_hi_lo_33 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_34 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_34 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_34 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_34 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_34 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_34 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_34 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_34 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_34 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_34 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_34 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_32 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_32 ={ core_csr_decoded_decoded_andMatrixInput_9_34 , core_csr_decoded_decoded_andMatrixInput_10_34 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_34 ={ core_csr_decoded_decoded_lo_lo_hi_32 , core_csr_decoded_decoded_andMatrixInput_11_32 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_6_34 , core_csr_decoded_decoded_andMatrixInput_7_34 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_34 ={ core_csr_decoded_decoded_lo_hi_hi_34 , core_csr_decoded_decoded_andMatrixInput_8_34 }; 
    wire[5:0] core_csr_decoded_decoded_lo_34 ={ core_csr_decoded_decoded_lo_hi_34 , core_csr_decoded_decoded_lo_lo_34 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_3_34 , core_csr_decoded_decoded_andMatrixInput_4_34 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_34 ={ core_csr_decoded_decoded_hi_lo_hi_34 , core_csr_decoded_decoded_andMatrixInput_5_34 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_0_34 , core_csr_decoded_decoded_andMatrixInput_1_34 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_34 ={ core_csr_decoded_decoded_hi_hi_hi_34 , core_csr_decoded_decoded_andMatrixInput_2_34 }; 
    wire[5:0] core_csr_decoded_decoded_hi_34 ={ core_csr_decoded_decoded_hi_hi_34 , core_csr_decoded_decoded_hi_lo_34 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_35 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_35 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_35 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_35 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_35 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_35 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_35 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_35 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_35 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_35 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_35 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_33 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_33 ={ core_csr_decoded_decoded_andMatrixInput_9_35 , core_csr_decoded_decoded_andMatrixInput_10_35 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_35 ={ core_csr_decoded_decoded_lo_lo_hi_33 , core_csr_decoded_decoded_andMatrixInput_11_33 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_6_35 , core_csr_decoded_decoded_andMatrixInput_7_35 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_35 ={ core_csr_decoded_decoded_lo_hi_hi_35 , core_csr_decoded_decoded_andMatrixInput_8_35 }; 
    wire[5:0] core_csr_decoded_decoded_lo_35 ={ core_csr_decoded_decoded_lo_hi_35 , core_csr_decoded_decoded_lo_lo_35 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_3_35 , core_csr_decoded_decoded_andMatrixInput_4_35 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_35 ={ core_csr_decoded_decoded_hi_lo_hi_35 , core_csr_decoded_decoded_andMatrixInput_5_35 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_0_35 , core_csr_decoded_decoded_andMatrixInput_1_35 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_35 ={ core_csr_decoded_decoded_hi_hi_hi_35 , core_csr_decoded_decoded_andMatrixInput_2_35 }; 
    wire[5:0] core_csr_decoded_decoded_hi_35 ={ core_csr_decoded_decoded_hi_hi_35 , core_csr_decoded_decoded_hi_lo_35 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_36 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_36 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_36 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_36 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_36 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_36 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_36 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_36 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_36 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_36 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_36 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_34 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_34 ={ core_csr_decoded_decoded_andMatrixInput_9_36 , core_csr_decoded_decoded_andMatrixInput_10_36 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_36 ={ core_csr_decoded_decoded_lo_lo_hi_34 , core_csr_decoded_decoded_andMatrixInput_11_34 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_6_36 , core_csr_decoded_decoded_andMatrixInput_7_36 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_36 ={ core_csr_decoded_decoded_lo_hi_hi_36 , core_csr_decoded_decoded_andMatrixInput_8_36 }; 
    wire[5:0] core_csr_decoded_decoded_lo_36 ={ core_csr_decoded_decoded_lo_hi_36 , core_csr_decoded_decoded_lo_lo_36 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_3_36 , core_csr_decoded_decoded_andMatrixInput_4_36 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_36 ={ core_csr_decoded_decoded_hi_lo_hi_36 , core_csr_decoded_decoded_andMatrixInput_5_36 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_0_36 , core_csr_decoded_decoded_andMatrixInput_1_36 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_36 ={ core_csr_decoded_decoded_hi_hi_hi_36 , core_csr_decoded_decoded_andMatrixInput_2_36 }; 
    wire[5:0] core_csr_decoded_decoded_hi_36 ={ core_csr_decoded_decoded_hi_hi_36 , core_csr_decoded_decoded_hi_lo_36 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_37 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_37 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_37 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_37 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_37 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_37 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_37 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_37 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_37 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_37 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_37 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_35 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_35 ={ core_csr_decoded_decoded_andMatrixInput_9_37 , core_csr_decoded_decoded_andMatrixInput_10_37 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_37 ={ core_csr_decoded_decoded_lo_lo_hi_35 , core_csr_decoded_decoded_andMatrixInput_11_35 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_6_37 , core_csr_decoded_decoded_andMatrixInput_7_37 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_37 ={ core_csr_decoded_decoded_lo_hi_hi_37 , core_csr_decoded_decoded_andMatrixInput_8_37 }; 
    wire[5:0] core_csr_decoded_decoded_lo_37 ={ core_csr_decoded_decoded_lo_hi_37 , core_csr_decoded_decoded_lo_lo_37 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_3_37 , core_csr_decoded_decoded_andMatrixInput_4_37 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_37 ={ core_csr_decoded_decoded_hi_lo_hi_37 , core_csr_decoded_decoded_andMatrixInput_5_37 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_0_37 , core_csr_decoded_decoded_andMatrixInput_1_37 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_37 ={ core_csr_decoded_decoded_hi_hi_hi_37 , core_csr_decoded_decoded_andMatrixInput_2_37 }; 
    wire[5:0] core_csr_decoded_decoded_hi_37 ={ core_csr_decoded_decoded_hi_hi_37 , core_csr_decoded_decoded_hi_lo_37 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_38 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_38 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_38 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_38 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_38 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_38 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_38 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_38 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_38 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_38 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_38 ={ core_csr_decoded_decoded_andMatrixInput_8_38 , core_csr_decoded_decoded_andMatrixInput_9_38 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_5_38 , core_csr_decoded_decoded_andMatrixInput_6_38 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_38 ={ core_csr_decoded_decoded_lo_hi_hi_38 , core_csr_decoded_decoded_andMatrixInput_7_38 }; 
    wire[4:0] core_csr_decoded_decoded_lo_38 ={ core_csr_decoded_decoded_lo_hi_38 , core_csr_decoded_decoded_lo_lo_38 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_38 ={ core_csr_decoded_decoded_andMatrixInput_3_38 , core_csr_decoded_decoded_andMatrixInput_4_38 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_0_38 , core_csr_decoded_decoded_andMatrixInput_1_38 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_38 ={ core_csr_decoded_decoded_hi_hi_hi_38 , core_csr_decoded_decoded_andMatrixInput_2_38 }; 
    wire[4:0] core_csr_decoded_decoded_hi_38 ={ core_csr_decoded_decoded_hi_hi_38 , core_csr_decoded_decoded_hi_lo_38 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_39 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_39 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_39 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_39 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_39 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_39 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_39 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_39 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_39 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_39 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_38 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_39 ={ core_csr_decoded_decoded_andMatrixInput_9_39 , core_csr_decoded_decoded_andMatrixInput_10_38 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_6_39 , core_csr_decoded_decoded_andMatrixInput_7_39 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_39 ={ core_csr_decoded_decoded_lo_hi_hi_39 , core_csr_decoded_decoded_andMatrixInput_8_39 }; 
    wire[4:0] core_csr_decoded_decoded_lo_39 ={ core_csr_decoded_decoded_lo_hi_39 , core_csr_decoded_decoded_lo_lo_39 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_3_39 , core_csr_decoded_decoded_andMatrixInput_4_39 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_39 ={ core_csr_decoded_decoded_hi_lo_hi_38 , core_csr_decoded_decoded_andMatrixInput_5_39 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_0_39 , core_csr_decoded_decoded_andMatrixInput_1_39 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_39 ={ core_csr_decoded_decoded_hi_hi_hi_39 , core_csr_decoded_decoded_andMatrixInput_2_39 }; 
    wire[5:0] core_csr_decoded_decoded_hi_39 ={ core_csr_decoded_decoded_hi_hi_39 , core_csr_decoded_decoded_hi_lo_39 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_40 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_40 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_40 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_40 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_40 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_40 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_40 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_40 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_40 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_40 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_39 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_40 ={ core_csr_decoded_decoded_andMatrixInput_9_40 , core_csr_decoded_decoded_andMatrixInput_10_39 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_6_40 , core_csr_decoded_decoded_andMatrixInput_7_40 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_40 ={ core_csr_decoded_decoded_lo_hi_hi_40 , core_csr_decoded_decoded_andMatrixInput_8_40 }; 
    wire[4:0] core_csr_decoded_decoded_lo_40 ={ core_csr_decoded_decoded_lo_hi_40 , core_csr_decoded_decoded_lo_lo_40 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_3_40 , core_csr_decoded_decoded_andMatrixInput_4_40 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_40 ={ core_csr_decoded_decoded_hi_lo_hi_39 , core_csr_decoded_decoded_andMatrixInput_5_40 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_0_40 , core_csr_decoded_decoded_andMatrixInput_1_40 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_40 ={ core_csr_decoded_decoded_hi_hi_hi_40 , core_csr_decoded_decoded_andMatrixInput_2_40 }; 
    wire[5:0] core_csr_decoded_decoded_hi_40 ={ core_csr_decoded_decoded_hi_hi_40 , core_csr_decoded_decoded_hi_lo_40 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_41 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_41 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_41 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_41 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_41 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_41 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_41 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_41 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_41 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_41 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_40 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_36 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_36 ={ core_csr_decoded_decoded_andMatrixInput_9_41 , core_csr_decoded_decoded_andMatrixInput_10_40 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_41 ={ core_csr_decoded_decoded_lo_lo_hi_36 , core_csr_decoded_decoded_andMatrixInput_11_36 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_6_41 , core_csr_decoded_decoded_andMatrixInput_7_41 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_41 ={ core_csr_decoded_decoded_lo_hi_hi_41 , core_csr_decoded_decoded_andMatrixInput_8_41 }; 
    wire[5:0] core_csr_decoded_decoded_lo_41 ={ core_csr_decoded_decoded_lo_hi_41 , core_csr_decoded_decoded_lo_lo_41 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_3_41 , core_csr_decoded_decoded_andMatrixInput_4_41 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_41 ={ core_csr_decoded_decoded_hi_lo_hi_40 , core_csr_decoded_decoded_andMatrixInput_5_41 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_0_41 , core_csr_decoded_decoded_andMatrixInput_1_41 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_41 ={ core_csr_decoded_decoded_hi_hi_hi_41 , core_csr_decoded_decoded_andMatrixInput_2_41 }; 
    wire[5:0] core_csr_decoded_decoded_hi_41 ={ core_csr_decoded_decoded_hi_hi_41 , core_csr_decoded_decoded_hi_lo_41 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_42 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_42 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_42 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_42 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_42 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_42 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_42 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_42 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_42 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_42 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_41 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_37 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_37 ={ core_csr_decoded_decoded_andMatrixInput_9_42 , core_csr_decoded_decoded_andMatrixInput_10_41 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_42 ={ core_csr_decoded_decoded_lo_lo_hi_37 , core_csr_decoded_decoded_andMatrixInput_11_37 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_6_42 , core_csr_decoded_decoded_andMatrixInput_7_42 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_42 ={ core_csr_decoded_decoded_lo_hi_hi_42 , core_csr_decoded_decoded_andMatrixInput_8_42 }; 
    wire[5:0] core_csr_decoded_decoded_lo_42 ={ core_csr_decoded_decoded_lo_hi_42 , core_csr_decoded_decoded_lo_lo_42 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_3_42 , core_csr_decoded_decoded_andMatrixInput_4_42 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_42 ={ core_csr_decoded_decoded_hi_lo_hi_41 , core_csr_decoded_decoded_andMatrixInput_5_42 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_0_42 , core_csr_decoded_decoded_andMatrixInput_1_42 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_42 ={ core_csr_decoded_decoded_hi_hi_hi_42 , core_csr_decoded_decoded_andMatrixInput_2_42 }; 
    wire[5:0] core_csr_decoded_decoded_hi_42 ={ core_csr_decoded_decoded_hi_hi_42 , core_csr_decoded_decoded_hi_lo_42 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_43 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_43 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_43 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_43 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_43 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_43 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_43 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_43 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_43 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_43 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_42 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_38 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_38 ={ core_csr_decoded_decoded_andMatrixInput_9_43 , core_csr_decoded_decoded_andMatrixInput_10_42 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_43 ={ core_csr_decoded_decoded_lo_lo_hi_38 , core_csr_decoded_decoded_andMatrixInput_11_38 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_6_43 , core_csr_decoded_decoded_andMatrixInput_7_43 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_43 ={ core_csr_decoded_decoded_lo_hi_hi_43 , core_csr_decoded_decoded_andMatrixInput_8_43 }; 
    wire[5:0] core_csr_decoded_decoded_lo_43 ={ core_csr_decoded_decoded_lo_hi_43 , core_csr_decoded_decoded_lo_lo_43 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_3_43 , core_csr_decoded_decoded_andMatrixInput_4_43 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_43 ={ core_csr_decoded_decoded_hi_lo_hi_42 , core_csr_decoded_decoded_andMatrixInput_5_43 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_0_43 , core_csr_decoded_decoded_andMatrixInput_1_43 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_43 ={ core_csr_decoded_decoded_hi_hi_hi_43 , core_csr_decoded_decoded_andMatrixInput_2_43 }; 
    wire[5:0] core_csr_decoded_decoded_hi_43 ={ core_csr_decoded_decoded_hi_hi_43 , core_csr_decoded_decoded_hi_lo_43 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_44 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_44 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_44 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_44 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_44 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_44 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_44 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_44 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_44 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_44 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_43 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_39 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_39 ={ core_csr_decoded_decoded_andMatrixInput_9_44 , core_csr_decoded_decoded_andMatrixInput_10_43 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_44 ={ core_csr_decoded_decoded_lo_lo_hi_39 , core_csr_decoded_decoded_andMatrixInput_11_39 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_6_44 , core_csr_decoded_decoded_andMatrixInput_7_44 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_44 ={ core_csr_decoded_decoded_lo_hi_hi_44 , core_csr_decoded_decoded_andMatrixInput_8_44 }; 
    wire[5:0] core_csr_decoded_decoded_lo_44 ={ core_csr_decoded_decoded_lo_hi_44 , core_csr_decoded_decoded_lo_lo_44 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_3_44 , core_csr_decoded_decoded_andMatrixInput_4_44 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_44 ={ core_csr_decoded_decoded_hi_lo_hi_43 , core_csr_decoded_decoded_andMatrixInput_5_44 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_0_44 , core_csr_decoded_decoded_andMatrixInput_1_44 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_44 ={ core_csr_decoded_decoded_hi_hi_hi_44 , core_csr_decoded_decoded_andMatrixInput_2_44 }; 
    wire[5:0] core_csr_decoded_decoded_hi_44 ={ core_csr_decoded_decoded_hi_hi_44 , core_csr_decoded_decoded_hi_lo_44 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_45 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_45 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_45 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_45 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_45 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_45 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_45 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_45 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_45 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_45 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_44 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_40 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_40 ={ core_csr_decoded_decoded_andMatrixInput_9_45 , core_csr_decoded_decoded_andMatrixInput_10_44 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_45 ={ core_csr_decoded_decoded_lo_lo_hi_40 , core_csr_decoded_decoded_andMatrixInput_11_40 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_6_45 , core_csr_decoded_decoded_andMatrixInput_7_45 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_45 ={ core_csr_decoded_decoded_lo_hi_hi_45 , core_csr_decoded_decoded_andMatrixInput_8_45 }; 
    wire[5:0] core_csr_decoded_decoded_lo_45 ={ core_csr_decoded_decoded_lo_hi_45 , core_csr_decoded_decoded_lo_lo_45 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_3_45 , core_csr_decoded_decoded_andMatrixInput_4_45 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_45 ={ core_csr_decoded_decoded_hi_lo_hi_44 , core_csr_decoded_decoded_andMatrixInput_5_45 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_0_45 , core_csr_decoded_decoded_andMatrixInput_1_45 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_45 ={ core_csr_decoded_decoded_hi_hi_hi_45 , core_csr_decoded_decoded_andMatrixInput_2_45 }; 
    wire[5:0] core_csr_decoded_decoded_hi_45 ={ core_csr_decoded_decoded_hi_hi_45 , core_csr_decoded_decoded_hi_lo_45 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_46 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_46 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_46 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_46 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_46 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_46 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_46 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_46 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_46 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_46 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_45 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_41 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_41 ={ core_csr_decoded_decoded_andMatrixInput_9_46 , core_csr_decoded_decoded_andMatrixInput_10_45 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_46 ={ core_csr_decoded_decoded_lo_lo_hi_41 , core_csr_decoded_decoded_andMatrixInput_11_41 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_6_46 , core_csr_decoded_decoded_andMatrixInput_7_46 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_46 ={ core_csr_decoded_decoded_lo_hi_hi_46 , core_csr_decoded_decoded_andMatrixInput_8_46 }; 
    wire[5:0] core_csr_decoded_decoded_lo_46 ={ core_csr_decoded_decoded_lo_hi_46 , core_csr_decoded_decoded_lo_lo_46 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_3_46 , core_csr_decoded_decoded_andMatrixInput_4_46 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_46 ={ core_csr_decoded_decoded_hi_lo_hi_45 , core_csr_decoded_decoded_andMatrixInput_5_46 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_0_46 , core_csr_decoded_decoded_andMatrixInput_1_46 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_46 ={ core_csr_decoded_decoded_hi_hi_hi_46 , core_csr_decoded_decoded_andMatrixInput_2_46 }; 
    wire[5:0] core_csr_decoded_decoded_hi_46 ={ core_csr_decoded_decoded_hi_hi_46 , core_csr_decoded_decoded_hi_lo_46 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_47 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_47 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_47 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_47 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_47 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_47 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_47 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_47 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_47 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_47 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_46 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_42 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_42 ={ core_csr_decoded_decoded_andMatrixInput_9_47 , core_csr_decoded_decoded_andMatrixInput_10_46 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_47 ={ core_csr_decoded_decoded_lo_lo_hi_42 , core_csr_decoded_decoded_andMatrixInput_11_42 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_6_47 , core_csr_decoded_decoded_andMatrixInput_7_47 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_47 ={ core_csr_decoded_decoded_lo_hi_hi_47 , core_csr_decoded_decoded_andMatrixInput_8_47 }; 
    wire[5:0] core_csr_decoded_decoded_lo_47 ={ core_csr_decoded_decoded_lo_hi_47 , core_csr_decoded_decoded_lo_lo_47 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_3_47 , core_csr_decoded_decoded_andMatrixInput_4_47 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_47 ={ core_csr_decoded_decoded_hi_lo_hi_46 , core_csr_decoded_decoded_andMatrixInput_5_47 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_0_47 , core_csr_decoded_decoded_andMatrixInput_1_47 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_47 ={ core_csr_decoded_decoded_hi_hi_hi_47 , core_csr_decoded_decoded_andMatrixInput_2_47 }; 
    wire[5:0] core_csr_decoded_decoded_hi_47 ={ core_csr_decoded_decoded_hi_hi_47 , core_csr_decoded_decoded_hi_lo_47 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_48 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_48 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_48 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_48 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_48 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_48 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_48 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_48 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_48 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_48 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_47 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_43 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_43 ={ core_csr_decoded_decoded_andMatrixInput_9_48 , core_csr_decoded_decoded_andMatrixInput_10_47 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_48 ={ core_csr_decoded_decoded_lo_lo_hi_43 , core_csr_decoded_decoded_andMatrixInput_11_43 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_6_48 , core_csr_decoded_decoded_andMatrixInput_7_48 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_48 ={ core_csr_decoded_decoded_lo_hi_hi_48 , core_csr_decoded_decoded_andMatrixInput_8_48 }; 
    wire[5:0] core_csr_decoded_decoded_lo_48 ={ core_csr_decoded_decoded_lo_hi_48 , core_csr_decoded_decoded_lo_lo_48 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_3_48 , core_csr_decoded_decoded_andMatrixInput_4_48 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_48 ={ core_csr_decoded_decoded_hi_lo_hi_47 , core_csr_decoded_decoded_andMatrixInput_5_48 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_0_48 , core_csr_decoded_decoded_andMatrixInput_1_48 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_48 ={ core_csr_decoded_decoded_hi_hi_hi_48 , core_csr_decoded_decoded_andMatrixInput_2_48 }; 
    wire[5:0] core_csr_decoded_decoded_hi_48 ={ core_csr_decoded_decoded_hi_hi_48 , core_csr_decoded_decoded_hi_lo_48 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_49 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_49 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_49 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_49 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_49 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_49 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_49 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_49 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_49 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_49 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_48 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_44 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_44 ={ core_csr_decoded_decoded_andMatrixInput_9_49 , core_csr_decoded_decoded_andMatrixInput_10_48 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_49 ={ core_csr_decoded_decoded_lo_lo_hi_44 , core_csr_decoded_decoded_andMatrixInput_11_44 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_6_49 , core_csr_decoded_decoded_andMatrixInput_7_49 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_49 ={ core_csr_decoded_decoded_lo_hi_hi_49 , core_csr_decoded_decoded_andMatrixInput_8_49 }; 
    wire[5:0] core_csr_decoded_decoded_lo_49 ={ core_csr_decoded_decoded_lo_hi_49 , core_csr_decoded_decoded_lo_lo_49 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_3_49 , core_csr_decoded_decoded_andMatrixInput_4_49 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_49 ={ core_csr_decoded_decoded_hi_lo_hi_48 , core_csr_decoded_decoded_andMatrixInput_5_49 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_0_49 , core_csr_decoded_decoded_andMatrixInput_1_49 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_49 ={ core_csr_decoded_decoded_hi_hi_hi_49 , core_csr_decoded_decoded_andMatrixInput_2_49 }; 
    wire[5:0] core_csr_decoded_decoded_hi_49 ={ core_csr_decoded_decoded_hi_hi_49 , core_csr_decoded_decoded_hi_lo_49 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_50 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_50 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_50 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_50 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_50 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_50 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_50 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_50 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_50 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_50 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_49 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_45 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_45 ={ core_csr_decoded_decoded_andMatrixInput_9_50 , core_csr_decoded_decoded_andMatrixInput_10_49 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_50 ={ core_csr_decoded_decoded_lo_lo_hi_45 , core_csr_decoded_decoded_andMatrixInput_11_45 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_6_50 , core_csr_decoded_decoded_andMatrixInput_7_50 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_50 ={ core_csr_decoded_decoded_lo_hi_hi_50 , core_csr_decoded_decoded_andMatrixInput_8_50 }; 
    wire[5:0] core_csr_decoded_decoded_lo_50 ={ core_csr_decoded_decoded_lo_hi_50 , core_csr_decoded_decoded_lo_lo_50 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_3_50 , core_csr_decoded_decoded_andMatrixInput_4_50 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_50 ={ core_csr_decoded_decoded_hi_lo_hi_49 , core_csr_decoded_decoded_andMatrixInput_5_50 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_0_50 , core_csr_decoded_decoded_andMatrixInput_1_50 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_50 ={ core_csr_decoded_decoded_hi_hi_hi_50 , core_csr_decoded_decoded_andMatrixInput_2_50 }; 
    wire[5:0] core_csr_decoded_decoded_hi_50 ={ core_csr_decoded_decoded_hi_hi_50 , core_csr_decoded_decoded_hi_lo_50 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_51 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_51 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_51 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_51 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_51 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_51 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_51 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_51 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_51 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_51 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_50 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_46 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_46 ={ core_csr_decoded_decoded_andMatrixInput_9_51 , core_csr_decoded_decoded_andMatrixInput_10_50 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_51 ={ core_csr_decoded_decoded_lo_lo_hi_46 , core_csr_decoded_decoded_andMatrixInput_11_46 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_6_51 , core_csr_decoded_decoded_andMatrixInput_7_51 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_51 ={ core_csr_decoded_decoded_lo_hi_hi_51 , core_csr_decoded_decoded_andMatrixInput_8_51 }; 
    wire[5:0] core_csr_decoded_decoded_lo_51 ={ core_csr_decoded_decoded_lo_hi_51 , core_csr_decoded_decoded_lo_lo_51 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_3_51 , core_csr_decoded_decoded_andMatrixInput_4_51 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_51 ={ core_csr_decoded_decoded_hi_lo_hi_50 , core_csr_decoded_decoded_andMatrixInput_5_51 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_0_51 , core_csr_decoded_decoded_andMatrixInput_1_51 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_51 ={ core_csr_decoded_decoded_hi_hi_hi_51 , core_csr_decoded_decoded_andMatrixInput_2_51 }; 
    wire[5:0] core_csr_decoded_decoded_hi_51 ={ core_csr_decoded_decoded_hi_hi_51 , core_csr_decoded_decoded_hi_lo_51 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_52 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_52 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_52 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_52 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_52 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_52 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_52 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_52 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_52 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_52 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_51 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_47 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_47 ={ core_csr_decoded_decoded_andMatrixInput_9_52 , core_csr_decoded_decoded_andMatrixInput_10_51 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_52 ={ core_csr_decoded_decoded_lo_lo_hi_47 , core_csr_decoded_decoded_andMatrixInput_11_47 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_6_52 , core_csr_decoded_decoded_andMatrixInput_7_52 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_52 ={ core_csr_decoded_decoded_lo_hi_hi_52 , core_csr_decoded_decoded_andMatrixInput_8_52 }; 
    wire[5:0] core_csr_decoded_decoded_lo_52 ={ core_csr_decoded_decoded_lo_hi_52 , core_csr_decoded_decoded_lo_lo_52 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_3_52 , core_csr_decoded_decoded_andMatrixInput_4_52 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_52 ={ core_csr_decoded_decoded_hi_lo_hi_51 , core_csr_decoded_decoded_andMatrixInput_5_52 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_0_52 , core_csr_decoded_decoded_andMatrixInput_1_52 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_52 ={ core_csr_decoded_decoded_hi_hi_hi_52 , core_csr_decoded_decoded_andMatrixInput_2_52 }; 
    wire[5:0] core_csr_decoded_decoded_hi_52 ={ core_csr_decoded_decoded_hi_hi_52 , core_csr_decoded_decoded_hi_lo_52 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_53 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_53 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_53 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_53 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_53 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_53 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_53 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_53 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_53 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_53 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_52 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_48 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_48 ={ core_csr_decoded_decoded_andMatrixInput_9_53 , core_csr_decoded_decoded_andMatrixInput_10_52 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_53 ={ core_csr_decoded_decoded_lo_lo_hi_48 , core_csr_decoded_decoded_andMatrixInput_11_48 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_6_53 , core_csr_decoded_decoded_andMatrixInput_7_53 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_53 ={ core_csr_decoded_decoded_lo_hi_hi_53 , core_csr_decoded_decoded_andMatrixInput_8_53 }; 
    wire[5:0] core_csr_decoded_decoded_lo_53 ={ core_csr_decoded_decoded_lo_hi_53 , core_csr_decoded_decoded_lo_lo_53 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_3_53 , core_csr_decoded_decoded_andMatrixInput_4_53 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_53 ={ core_csr_decoded_decoded_hi_lo_hi_52 , core_csr_decoded_decoded_andMatrixInput_5_53 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_0_53 , core_csr_decoded_decoded_andMatrixInput_1_53 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_53 ={ core_csr_decoded_decoded_hi_hi_hi_53 , core_csr_decoded_decoded_andMatrixInput_2_53 }; 
    wire[5:0] core_csr_decoded_decoded_hi_53 ={ core_csr_decoded_decoded_hi_hi_53 , core_csr_decoded_decoded_hi_lo_53 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_54 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_54 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_54 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_54 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_54 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_54 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_54 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_54 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_54 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_54 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_53 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_49 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_49 ={ core_csr_decoded_decoded_andMatrixInput_9_54 , core_csr_decoded_decoded_andMatrixInput_10_53 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_54 ={ core_csr_decoded_decoded_lo_lo_hi_49 , core_csr_decoded_decoded_andMatrixInput_11_49 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_6_54 , core_csr_decoded_decoded_andMatrixInput_7_54 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_54 ={ core_csr_decoded_decoded_lo_hi_hi_54 , core_csr_decoded_decoded_andMatrixInput_8_54 }; 
    wire[5:0] core_csr_decoded_decoded_lo_54 ={ core_csr_decoded_decoded_lo_hi_54 , core_csr_decoded_decoded_lo_lo_54 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_3_54 , core_csr_decoded_decoded_andMatrixInput_4_54 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_54 ={ core_csr_decoded_decoded_hi_lo_hi_53 , core_csr_decoded_decoded_andMatrixInput_5_54 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_0_54 , core_csr_decoded_decoded_andMatrixInput_1_54 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_54 ={ core_csr_decoded_decoded_hi_hi_hi_54 , core_csr_decoded_decoded_andMatrixInput_2_54 }; 
    wire[5:0] core_csr_decoded_decoded_hi_54 ={ core_csr_decoded_decoded_hi_hi_54 , core_csr_decoded_decoded_hi_lo_54 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_55 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_55 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_55 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_55 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_55 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_55 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_55 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_55 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_55 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_55 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_54 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_50 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_50 ={ core_csr_decoded_decoded_andMatrixInput_9_55 , core_csr_decoded_decoded_andMatrixInput_10_54 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_55 ={ core_csr_decoded_decoded_lo_lo_hi_50 , core_csr_decoded_decoded_andMatrixInput_11_50 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_6_55 , core_csr_decoded_decoded_andMatrixInput_7_55 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_55 ={ core_csr_decoded_decoded_lo_hi_hi_55 , core_csr_decoded_decoded_andMatrixInput_8_55 }; 
    wire[5:0] core_csr_decoded_decoded_lo_55 ={ core_csr_decoded_decoded_lo_hi_55 , core_csr_decoded_decoded_lo_lo_55 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_3_55 , core_csr_decoded_decoded_andMatrixInput_4_55 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_55 ={ core_csr_decoded_decoded_hi_lo_hi_54 , core_csr_decoded_decoded_andMatrixInput_5_55 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_0_55 , core_csr_decoded_decoded_andMatrixInput_1_55 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_55 ={ core_csr_decoded_decoded_hi_hi_hi_55 , core_csr_decoded_decoded_andMatrixInput_2_55 }; 
    wire[5:0] core_csr_decoded_decoded_hi_55 ={ core_csr_decoded_decoded_hi_hi_55 , core_csr_decoded_decoded_hi_lo_55 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_56 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_56 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_56 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_56 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_56 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_56 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_56 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_56 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_56 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_56 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_55 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_51 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_51 ={ core_csr_decoded_decoded_andMatrixInput_9_56 , core_csr_decoded_decoded_andMatrixInput_10_55 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_56 ={ core_csr_decoded_decoded_lo_lo_hi_51 , core_csr_decoded_decoded_andMatrixInput_11_51 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_6_56 , core_csr_decoded_decoded_andMatrixInput_7_56 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_56 ={ core_csr_decoded_decoded_lo_hi_hi_56 , core_csr_decoded_decoded_andMatrixInput_8_56 }; 
    wire[5:0] core_csr_decoded_decoded_lo_56 ={ core_csr_decoded_decoded_lo_hi_56 , core_csr_decoded_decoded_lo_lo_56 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_3_56 , core_csr_decoded_decoded_andMatrixInput_4_56 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_56 ={ core_csr_decoded_decoded_hi_lo_hi_55 , core_csr_decoded_decoded_andMatrixInput_5_56 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_0_56 , core_csr_decoded_decoded_andMatrixInput_1_56 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_56 ={ core_csr_decoded_decoded_hi_hi_hi_56 , core_csr_decoded_decoded_andMatrixInput_2_56 }; 
    wire[5:0] core_csr_decoded_decoded_hi_56 ={ core_csr_decoded_decoded_hi_hi_56 , core_csr_decoded_decoded_hi_lo_56 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_57 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_57 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_57 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_57 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_57 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_57 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_57 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_57 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_57 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_57 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_56 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_52 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_52 ={ core_csr_decoded_decoded_andMatrixInput_9_57 , core_csr_decoded_decoded_andMatrixInput_10_56 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_57 ={ core_csr_decoded_decoded_lo_lo_hi_52 , core_csr_decoded_decoded_andMatrixInput_11_52 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_6_57 , core_csr_decoded_decoded_andMatrixInput_7_57 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_57 ={ core_csr_decoded_decoded_lo_hi_hi_57 , core_csr_decoded_decoded_andMatrixInput_8_57 }; 
    wire[5:0] core_csr_decoded_decoded_lo_57 ={ core_csr_decoded_decoded_lo_hi_57 , core_csr_decoded_decoded_lo_lo_57 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_3_57 , core_csr_decoded_decoded_andMatrixInput_4_57 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_57 ={ core_csr_decoded_decoded_hi_lo_hi_56 , core_csr_decoded_decoded_andMatrixInput_5_57 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_0_57 , core_csr_decoded_decoded_andMatrixInput_1_57 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_57 ={ core_csr_decoded_decoded_hi_hi_hi_57 , core_csr_decoded_decoded_andMatrixInput_2_57 }; 
    wire[5:0] core_csr_decoded_decoded_hi_57 ={ core_csr_decoded_decoded_hi_hi_57 , core_csr_decoded_decoded_hi_lo_57 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_58 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_58 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_58 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_58 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_58 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_58 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_58 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_58 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_58 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_58 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_57 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_53 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_53 ={ core_csr_decoded_decoded_andMatrixInput_9_58 , core_csr_decoded_decoded_andMatrixInput_10_57 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_58 ={ core_csr_decoded_decoded_lo_lo_hi_53 , core_csr_decoded_decoded_andMatrixInput_11_53 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_6_58 , core_csr_decoded_decoded_andMatrixInput_7_58 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_58 ={ core_csr_decoded_decoded_lo_hi_hi_58 , core_csr_decoded_decoded_andMatrixInput_8_58 }; 
    wire[5:0] core_csr_decoded_decoded_lo_58 ={ core_csr_decoded_decoded_lo_hi_58 , core_csr_decoded_decoded_lo_lo_58 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_3_58 , core_csr_decoded_decoded_andMatrixInput_4_58 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_58 ={ core_csr_decoded_decoded_hi_lo_hi_57 , core_csr_decoded_decoded_andMatrixInput_5_58 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_0_58 , core_csr_decoded_decoded_andMatrixInput_1_58 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_58 ={ core_csr_decoded_decoded_hi_hi_hi_58 , core_csr_decoded_decoded_andMatrixInput_2_58 }; 
    wire[5:0] core_csr_decoded_decoded_hi_58 ={ core_csr_decoded_decoded_hi_hi_58 , core_csr_decoded_decoded_hi_lo_58 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_59 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_59 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_59 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_59 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_59 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_59 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_59 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_59 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_59 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_59 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_58 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_54 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_54 ={ core_csr_decoded_decoded_andMatrixInput_9_59 , core_csr_decoded_decoded_andMatrixInput_10_58 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_59 ={ core_csr_decoded_decoded_lo_lo_hi_54 , core_csr_decoded_decoded_andMatrixInput_11_54 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_6_59 , core_csr_decoded_decoded_andMatrixInput_7_59 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_59 ={ core_csr_decoded_decoded_lo_hi_hi_59 , core_csr_decoded_decoded_andMatrixInput_8_59 }; 
    wire[5:0] core_csr_decoded_decoded_lo_59 ={ core_csr_decoded_decoded_lo_hi_59 , core_csr_decoded_decoded_lo_lo_59 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_3_59 , core_csr_decoded_decoded_andMatrixInput_4_59 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_59 ={ core_csr_decoded_decoded_hi_lo_hi_58 , core_csr_decoded_decoded_andMatrixInput_5_59 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_0_59 , core_csr_decoded_decoded_andMatrixInput_1_59 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_59 ={ core_csr_decoded_decoded_hi_hi_hi_59 , core_csr_decoded_decoded_andMatrixInput_2_59 }; 
    wire[5:0] core_csr_decoded_decoded_hi_59 ={ core_csr_decoded_decoded_hi_hi_59 , core_csr_decoded_decoded_hi_lo_59 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_60 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_60 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_60 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_60 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_60 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_60 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_60 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_60 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_60 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_60 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_59 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_55 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_55 ={ core_csr_decoded_decoded_andMatrixInput_9_60 , core_csr_decoded_decoded_andMatrixInput_10_59 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_60 ={ core_csr_decoded_decoded_lo_lo_hi_55 , core_csr_decoded_decoded_andMatrixInput_11_55 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_6_60 , core_csr_decoded_decoded_andMatrixInput_7_60 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_60 ={ core_csr_decoded_decoded_lo_hi_hi_60 , core_csr_decoded_decoded_andMatrixInput_8_60 }; 
    wire[5:0] core_csr_decoded_decoded_lo_60 ={ core_csr_decoded_decoded_lo_hi_60 , core_csr_decoded_decoded_lo_lo_60 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_3_60 , core_csr_decoded_decoded_andMatrixInput_4_60 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_60 ={ core_csr_decoded_decoded_hi_lo_hi_59 , core_csr_decoded_decoded_andMatrixInput_5_60 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_0_60 , core_csr_decoded_decoded_andMatrixInput_1_60 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_60 ={ core_csr_decoded_decoded_hi_hi_hi_60 , core_csr_decoded_decoded_andMatrixInput_2_60 }; 
    wire[5:0] core_csr_decoded_decoded_hi_60 ={ core_csr_decoded_decoded_hi_hi_60 , core_csr_decoded_decoded_hi_lo_60 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_61 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_61 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_61 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_61 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_61 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_61 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_61 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_61 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_61 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_61 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_60 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_56 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_56 ={ core_csr_decoded_decoded_andMatrixInput_9_61 , core_csr_decoded_decoded_andMatrixInput_10_60 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_61 ={ core_csr_decoded_decoded_lo_lo_hi_56 , core_csr_decoded_decoded_andMatrixInput_11_56 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_6_61 , core_csr_decoded_decoded_andMatrixInput_7_61 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_61 ={ core_csr_decoded_decoded_lo_hi_hi_61 , core_csr_decoded_decoded_andMatrixInput_8_61 }; 
    wire[5:0] core_csr_decoded_decoded_lo_61 ={ core_csr_decoded_decoded_lo_hi_61 , core_csr_decoded_decoded_lo_lo_61 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_3_61 , core_csr_decoded_decoded_andMatrixInput_4_61 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_61 ={ core_csr_decoded_decoded_hi_lo_hi_60 , core_csr_decoded_decoded_andMatrixInput_5_61 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_0_61 , core_csr_decoded_decoded_andMatrixInput_1_61 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_61 ={ core_csr_decoded_decoded_hi_hi_hi_61 , core_csr_decoded_decoded_andMatrixInput_2_61 }; 
    wire[5:0] core_csr_decoded_decoded_hi_61 ={ core_csr_decoded_decoded_hi_hi_61 , core_csr_decoded_decoded_hi_lo_61 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_62 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_62 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_62 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_62 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_62 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_62 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_62 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_62 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_62 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_62 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_61 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_57 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_57 ={ core_csr_decoded_decoded_andMatrixInput_9_62 , core_csr_decoded_decoded_andMatrixInput_10_61 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_62 ={ core_csr_decoded_decoded_lo_lo_hi_57 , core_csr_decoded_decoded_andMatrixInput_11_57 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_6_62 , core_csr_decoded_decoded_andMatrixInput_7_62 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_62 ={ core_csr_decoded_decoded_lo_hi_hi_62 , core_csr_decoded_decoded_andMatrixInput_8_62 }; 
    wire[5:0] core_csr_decoded_decoded_lo_62 ={ core_csr_decoded_decoded_lo_hi_62 , core_csr_decoded_decoded_lo_lo_62 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_3_62 , core_csr_decoded_decoded_andMatrixInput_4_62 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_62 ={ core_csr_decoded_decoded_hi_lo_hi_61 , core_csr_decoded_decoded_andMatrixInput_5_62 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_0_62 , core_csr_decoded_decoded_andMatrixInput_1_62 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_62 ={ core_csr_decoded_decoded_hi_hi_hi_62 , core_csr_decoded_decoded_andMatrixInput_2_62 }; 
    wire[5:0] core_csr_decoded_decoded_hi_62 ={ core_csr_decoded_decoded_hi_hi_62 , core_csr_decoded_decoded_hi_lo_62 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_63 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_63 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_63 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_63 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_63 = core_csr_decoded_decoded_plaInput [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_63 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_63 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_63 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_63 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_63 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_62 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_63 ={ core_csr_decoded_decoded_andMatrixInput_9_63 , core_csr_decoded_decoded_andMatrixInput_10_62 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_6_63 , core_csr_decoded_decoded_andMatrixInput_7_63 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_63 ={ core_csr_decoded_decoded_lo_hi_hi_63 , core_csr_decoded_decoded_andMatrixInput_8_63 }; 
    wire[4:0] core_csr_decoded_decoded_lo_63 ={ core_csr_decoded_decoded_lo_hi_63 , core_csr_decoded_decoded_lo_lo_63 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_3_63 , core_csr_decoded_decoded_andMatrixInput_4_63 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_63 ={ core_csr_decoded_decoded_hi_lo_hi_62 , core_csr_decoded_decoded_andMatrixInput_5_63 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_0_63 , core_csr_decoded_decoded_andMatrixInput_1_63 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_63 ={ core_csr_decoded_decoded_hi_hi_hi_63 , core_csr_decoded_decoded_andMatrixInput_2_63 }; 
    wire[5:0] core_csr_decoded_decoded_hi_63 ={ core_csr_decoded_decoded_hi_hi_63 , core_csr_decoded_decoded_hi_lo_63 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_64 = core_csr_decoded_decoded_plaInput [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_64 = core_csr_decoded_decoded_plaInput [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_64 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_64 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_64 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_64 = core_csr_decoded_decoded_invInputs [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_3_64 , core_csr_decoded_decoded_andMatrixInput_4_64 }; 
    wire[2:0] core_csr_decoded_decoded_lo_64 ={ core_csr_decoded_decoded_lo_hi_64 , core_csr_decoded_decoded_andMatrixInput_5_64 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_0_64 , core_csr_decoded_decoded_andMatrixInput_1_64 }; 
    wire[2:0] core_csr_decoded_decoded_hi_64 ={ core_csr_decoded_decoded_hi_hi_64 , core_csr_decoded_decoded_andMatrixInput_2_64 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_65 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_65 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_65 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_65 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_65 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_65 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_64 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_64 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_64 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_64 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_63 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_64 ={ core_csr_decoded_decoded_andMatrixInput_9_64 , core_csr_decoded_decoded_andMatrixInput_10_63 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_6_64 , core_csr_decoded_decoded_andMatrixInput_7_64 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_65 ={ core_csr_decoded_decoded_lo_hi_hi_64 , core_csr_decoded_decoded_andMatrixInput_8_64 }; 
    wire[4:0] core_csr_decoded_decoded_lo_65 ={ core_csr_decoded_decoded_lo_hi_65 , core_csr_decoded_decoded_lo_lo_64 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_3_65 , core_csr_decoded_decoded_andMatrixInput_4_65 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_64 ={ core_csr_decoded_decoded_hi_lo_hi_63 , core_csr_decoded_decoded_andMatrixInput_5_65 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_0_65 , core_csr_decoded_decoded_andMatrixInput_1_65 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_65 ={ core_csr_decoded_decoded_hi_hi_hi_64 , core_csr_decoded_decoded_andMatrixInput_2_65 }; 
    wire[5:0] core_csr_decoded_decoded_hi_65 ={ core_csr_decoded_decoded_hi_hi_65 , core_csr_decoded_decoded_hi_lo_64 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_66 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_66 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_66 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_66 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_66 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_66 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_65 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_65 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_65 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_65 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_64 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_58 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_58 ={ core_csr_decoded_decoded_andMatrixInput_9_65 , core_csr_decoded_decoded_andMatrixInput_10_64 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_65 ={ core_csr_decoded_decoded_lo_lo_hi_58 , core_csr_decoded_decoded_andMatrixInput_11_58 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_6_65 , core_csr_decoded_decoded_andMatrixInput_7_65 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_66 ={ core_csr_decoded_decoded_lo_hi_hi_65 , core_csr_decoded_decoded_andMatrixInput_8_65 }; 
    wire[5:0] core_csr_decoded_decoded_lo_66 ={ core_csr_decoded_decoded_lo_hi_66 , core_csr_decoded_decoded_lo_lo_65 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_3_66 , core_csr_decoded_decoded_andMatrixInput_4_66 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_65 ={ core_csr_decoded_decoded_hi_lo_hi_64 , core_csr_decoded_decoded_andMatrixInput_5_66 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_0_66 , core_csr_decoded_decoded_andMatrixInput_1_66 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_66 ={ core_csr_decoded_decoded_hi_hi_hi_65 , core_csr_decoded_decoded_andMatrixInput_2_66 }; 
    wire[5:0] core_csr_decoded_decoded_hi_66 ={ core_csr_decoded_decoded_hi_hi_66 , core_csr_decoded_decoded_hi_lo_65 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_67 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_67 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_67 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_67 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_67 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_67 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_66 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_66 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_66 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_66 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_65 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_59 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_59 ={ core_csr_decoded_decoded_andMatrixInput_9_66 , core_csr_decoded_decoded_andMatrixInput_10_65 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_66 ={ core_csr_decoded_decoded_lo_lo_hi_59 , core_csr_decoded_decoded_andMatrixInput_11_59 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_6_66 , core_csr_decoded_decoded_andMatrixInput_7_66 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_67 ={ core_csr_decoded_decoded_lo_hi_hi_66 , core_csr_decoded_decoded_andMatrixInput_8_66 }; 
    wire[5:0] core_csr_decoded_decoded_lo_67 ={ core_csr_decoded_decoded_lo_hi_67 , core_csr_decoded_decoded_lo_lo_66 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_3_67 , core_csr_decoded_decoded_andMatrixInput_4_67 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_66 ={ core_csr_decoded_decoded_hi_lo_hi_65 , core_csr_decoded_decoded_andMatrixInput_5_67 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_0_67 , core_csr_decoded_decoded_andMatrixInput_1_67 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_67 ={ core_csr_decoded_decoded_hi_hi_hi_66 , core_csr_decoded_decoded_andMatrixInput_2_67 }; 
    wire[5:0] core_csr_decoded_decoded_hi_67 ={ core_csr_decoded_decoded_hi_hi_67 , core_csr_decoded_decoded_hi_lo_66 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_68 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_68 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_68 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_68 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_68 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_68 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_67 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_67 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_67 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_67 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_66 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_60 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_60 ={ core_csr_decoded_decoded_andMatrixInput_9_67 , core_csr_decoded_decoded_andMatrixInput_10_66 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_67 ={ core_csr_decoded_decoded_lo_lo_hi_60 , core_csr_decoded_decoded_andMatrixInput_11_60 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_6_67 , core_csr_decoded_decoded_andMatrixInput_7_67 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_68 ={ core_csr_decoded_decoded_lo_hi_hi_67 , core_csr_decoded_decoded_andMatrixInput_8_67 }; 
    wire[5:0] core_csr_decoded_decoded_lo_68 ={ core_csr_decoded_decoded_lo_hi_68 , core_csr_decoded_decoded_lo_lo_67 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_3_68 , core_csr_decoded_decoded_andMatrixInput_4_68 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_67 ={ core_csr_decoded_decoded_hi_lo_hi_66 , core_csr_decoded_decoded_andMatrixInput_5_68 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_0_68 , core_csr_decoded_decoded_andMatrixInput_1_68 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_68 ={ core_csr_decoded_decoded_hi_hi_hi_67 , core_csr_decoded_decoded_andMatrixInput_2_68 }; 
    wire[5:0] core_csr_decoded_decoded_hi_68 ={ core_csr_decoded_decoded_hi_hi_68 , core_csr_decoded_decoded_hi_lo_67 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_69 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_69 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_69 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_69 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_69 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_69 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_68 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_68 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_68 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_68 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_67 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_61 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_61 ={ core_csr_decoded_decoded_andMatrixInput_9_68 , core_csr_decoded_decoded_andMatrixInput_10_67 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_68 ={ core_csr_decoded_decoded_lo_lo_hi_61 , core_csr_decoded_decoded_andMatrixInput_11_61 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_6_68 , core_csr_decoded_decoded_andMatrixInput_7_68 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_69 ={ core_csr_decoded_decoded_lo_hi_hi_68 , core_csr_decoded_decoded_andMatrixInput_8_68 }; 
    wire[5:0] core_csr_decoded_decoded_lo_69 ={ core_csr_decoded_decoded_lo_hi_69 , core_csr_decoded_decoded_lo_lo_68 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_3_69 , core_csr_decoded_decoded_andMatrixInput_4_69 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_68 ={ core_csr_decoded_decoded_hi_lo_hi_67 , core_csr_decoded_decoded_andMatrixInput_5_69 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_0_69 , core_csr_decoded_decoded_andMatrixInput_1_69 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_69 ={ core_csr_decoded_decoded_hi_hi_hi_68 , core_csr_decoded_decoded_andMatrixInput_2_69 }; 
    wire[5:0] core_csr_decoded_decoded_hi_69 ={ core_csr_decoded_decoded_hi_hi_69 , core_csr_decoded_decoded_hi_lo_68 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_70 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_70 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_70 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_70 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_70 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_70 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_69 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_69 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_69 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_69 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_68 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_62 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_62 ={ core_csr_decoded_decoded_andMatrixInput_9_69 , core_csr_decoded_decoded_andMatrixInput_10_68 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_69 ={ core_csr_decoded_decoded_lo_lo_hi_62 , core_csr_decoded_decoded_andMatrixInput_11_62 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_6_69 , core_csr_decoded_decoded_andMatrixInput_7_69 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_70 ={ core_csr_decoded_decoded_lo_hi_hi_69 , core_csr_decoded_decoded_andMatrixInput_8_69 }; 
    wire[5:0] core_csr_decoded_decoded_lo_70 ={ core_csr_decoded_decoded_lo_hi_70 , core_csr_decoded_decoded_lo_lo_69 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_3_70 , core_csr_decoded_decoded_andMatrixInput_4_70 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_69 ={ core_csr_decoded_decoded_hi_lo_hi_68 , core_csr_decoded_decoded_andMatrixInput_5_70 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_0_70 , core_csr_decoded_decoded_andMatrixInput_1_70 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_70 ={ core_csr_decoded_decoded_hi_hi_hi_69 , core_csr_decoded_decoded_andMatrixInput_2_70 }; 
    wire[5:0] core_csr_decoded_decoded_hi_70 ={ core_csr_decoded_decoded_hi_hi_70 , core_csr_decoded_decoded_hi_lo_69 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_71 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_71 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_71 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_71 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_71 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_71 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_70 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_70 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_70 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_70 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_69 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_63 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_63 ={ core_csr_decoded_decoded_andMatrixInput_9_70 , core_csr_decoded_decoded_andMatrixInput_10_69 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_70 ={ core_csr_decoded_decoded_lo_lo_hi_63 , core_csr_decoded_decoded_andMatrixInput_11_63 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_6_70 , core_csr_decoded_decoded_andMatrixInput_7_70 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_71 ={ core_csr_decoded_decoded_lo_hi_hi_70 , core_csr_decoded_decoded_andMatrixInput_8_70 }; 
    wire[5:0] core_csr_decoded_decoded_lo_71 ={ core_csr_decoded_decoded_lo_hi_71 , core_csr_decoded_decoded_lo_lo_70 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_3_71 , core_csr_decoded_decoded_andMatrixInput_4_71 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_70 ={ core_csr_decoded_decoded_hi_lo_hi_69 , core_csr_decoded_decoded_andMatrixInput_5_71 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_0_71 , core_csr_decoded_decoded_andMatrixInput_1_71 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_71 ={ core_csr_decoded_decoded_hi_hi_hi_70 , core_csr_decoded_decoded_andMatrixInput_2_71 }; 
    wire[5:0] core_csr_decoded_decoded_hi_71 ={ core_csr_decoded_decoded_hi_hi_71 , core_csr_decoded_decoded_hi_lo_70 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_72 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_72 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_72 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_72 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_72 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_72 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_71 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_71 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_71 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_71 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_70 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_64 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_64 ={ core_csr_decoded_decoded_andMatrixInput_9_71 , core_csr_decoded_decoded_andMatrixInput_10_70 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_71 ={ core_csr_decoded_decoded_lo_lo_hi_64 , core_csr_decoded_decoded_andMatrixInput_11_64 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_6_71 , core_csr_decoded_decoded_andMatrixInput_7_71 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_72 ={ core_csr_decoded_decoded_lo_hi_hi_71 , core_csr_decoded_decoded_andMatrixInput_8_71 }; 
    wire[5:0] core_csr_decoded_decoded_lo_72 ={ core_csr_decoded_decoded_lo_hi_72 , core_csr_decoded_decoded_lo_lo_71 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_3_72 , core_csr_decoded_decoded_andMatrixInput_4_72 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_71 ={ core_csr_decoded_decoded_hi_lo_hi_70 , core_csr_decoded_decoded_andMatrixInput_5_72 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_0_72 , core_csr_decoded_decoded_andMatrixInput_1_72 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_72 ={ core_csr_decoded_decoded_hi_hi_hi_71 , core_csr_decoded_decoded_andMatrixInput_2_72 }; 
    wire[5:0] core_csr_decoded_decoded_hi_72 ={ core_csr_decoded_decoded_hi_hi_72 , core_csr_decoded_decoded_hi_lo_71 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_73 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_73 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_73 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_73 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_73 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_73 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_72 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_72 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_72 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_72 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_71 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_65 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_65 ={ core_csr_decoded_decoded_andMatrixInput_9_72 , core_csr_decoded_decoded_andMatrixInput_10_71 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_72 ={ core_csr_decoded_decoded_lo_lo_hi_65 , core_csr_decoded_decoded_andMatrixInput_11_65 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_6_72 , core_csr_decoded_decoded_andMatrixInput_7_72 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_73 ={ core_csr_decoded_decoded_lo_hi_hi_72 , core_csr_decoded_decoded_andMatrixInput_8_72 }; 
    wire[5:0] core_csr_decoded_decoded_lo_73 ={ core_csr_decoded_decoded_lo_hi_73 , core_csr_decoded_decoded_lo_lo_72 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_3_73 , core_csr_decoded_decoded_andMatrixInput_4_73 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_72 ={ core_csr_decoded_decoded_hi_lo_hi_71 , core_csr_decoded_decoded_andMatrixInput_5_73 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_0_73 , core_csr_decoded_decoded_andMatrixInput_1_73 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_73 ={ core_csr_decoded_decoded_hi_hi_hi_72 , core_csr_decoded_decoded_andMatrixInput_2_73 }; 
    wire[5:0] core_csr_decoded_decoded_hi_73 ={ core_csr_decoded_decoded_hi_hi_73 , core_csr_decoded_decoded_hi_lo_72 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_74 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_74 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_74 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_74 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_74 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_74 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_73 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_73 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_73 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_73 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_72 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_66 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_66 ={ core_csr_decoded_decoded_andMatrixInput_9_73 , core_csr_decoded_decoded_andMatrixInput_10_72 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_73 ={ core_csr_decoded_decoded_lo_lo_hi_66 , core_csr_decoded_decoded_andMatrixInput_11_66 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_6_73 , core_csr_decoded_decoded_andMatrixInput_7_73 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_74 ={ core_csr_decoded_decoded_lo_hi_hi_73 , core_csr_decoded_decoded_andMatrixInput_8_73 }; 
    wire[5:0] core_csr_decoded_decoded_lo_74 ={ core_csr_decoded_decoded_lo_hi_74 , core_csr_decoded_decoded_lo_lo_73 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_3_74 , core_csr_decoded_decoded_andMatrixInput_4_74 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_73 ={ core_csr_decoded_decoded_hi_lo_hi_72 , core_csr_decoded_decoded_andMatrixInput_5_74 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_0_74 , core_csr_decoded_decoded_andMatrixInput_1_74 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_74 ={ core_csr_decoded_decoded_hi_hi_hi_73 , core_csr_decoded_decoded_andMatrixInput_2_74 }; 
    wire[5:0] core_csr_decoded_decoded_hi_74 ={ core_csr_decoded_decoded_hi_hi_74 , core_csr_decoded_decoded_hi_lo_73 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_75 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_75 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_75 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_75 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_75 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_75 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_74 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_74 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_74 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_74 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_73 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_67 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_67 ={ core_csr_decoded_decoded_andMatrixInput_9_74 , core_csr_decoded_decoded_andMatrixInput_10_73 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_74 ={ core_csr_decoded_decoded_lo_lo_hi_67 , core_csr_decoded_decoded_andMatrixInput_11_67 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_6_74 , core_csr_decoded_decoded_andMatrixInput_7_74 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_75 ={ core_csr_decoded_decoded_lo_hi_hi_74 , core_csr_decoded_decoded_andMatrixInput_8_74 }; 
    wire[5:0] core_csr_decoded_decoded_lo_75 ={ core_csr_decoded_decoded_lo_hi_75 , core_csr_decoded_decoded_lo_lo_74 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_3_75 , core_csr_decoded_decoded_andMatrixInput_4_75 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_74 ={ core_csr_decoded_decoded_hi_lo_hi_73 , core_csr_decoded_decoded_andMatrixInput_5_75 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_0_75 , core_csr_decoded_decoded_andMatrixInput_1_75 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_75 ={ core_csr_decoded_decoded_hi_hi_hi_74 , core_csr_decoded_decoded_andMatrixInput_2_75 }; 
    wire[5:0] core_csr_decoded_decoded_hi_75 ={ core_csr_decoded_decoded_hi_hi_75 , core_csr_decoded_decoded_hi_lo_74 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_76 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_76 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_76 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_76 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_76 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_76 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_75 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_75 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_75 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_75 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_74 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_68 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_68 ={ core_csr_decoded_decoded_andMatrixInput_9_75 , core_csr_decoded_decoded_andMatrixInput_10_74 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_75 ={ core_csr_decoded_decoded_lo_lo_hi_68 , core_csr_decoded_decoded_andMatrixInput_11_68 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_6_75 , core_csr_decoded_decoded_andMatrixInput_7_75 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_76 ={ core_csr_decoded_decoded_lo_hi_hi_75 , core_csr_decoded_decoded_andMatrixInput_8_75 }; 
    wire[5:0] core_csr_decoded_decoded_lo_76 ={ core_csr_decoded_decoded_lo_hi_76 , core_csr_decoded_decoded_lo_lo_75 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_3_76 , core_csr_decoded_decoded_andMatrixInput_4_76 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_75 ={ core_csr_decoded_decoded_hi_lo_hi_74 , core_csr_decoded_decoded_andMatrixInput_5_76 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_0_76 , core_csr_decoded_decoded_andMatrixInput_1_76 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_76 ={ core_csr_decoded_decoded_hi_hi_hi_75 , core_csr_decoded_decoded_andMatrixInput_2_76 }; 
    wire[5:0] core_csr_decoded_decoded_hi_76 ={ core_csr_decoded_decoded_hi_hi_76 , core_csr_decoded_decoded_hi_lo_75 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_77 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_77 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_77 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_77 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_77 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_77 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_76 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_76 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_76 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_76 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_75 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_69 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_69 ={ core_csr_decoded_decoded_andMatrixInput_9_76 , core_csr_decoded_decoded_andMatrixInput_10_75 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_76 ={ core_csr_decoded_decoded_lo_lo_hi_69 , core_csr_decoded_decoded_andMatrixInput_11_69 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_6_76 , core_csr_decoded_decoded_andMatrixInput_7_76 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_77 ={ core_csr_decoded_decoded_lo_hi_hi_76 , core_csr_decoded_decoded_andMatrixInput_8_76 }; 
    wire[5:0] core_csr_decoded_decoded_lo_77 ={ core_csr_decoded_decoded_lo_hi_77 , core_csr_decoded_decoded_lo_lo_76 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_3_77 , core_csr_decoded_decoded_andMatrixInput_4_77 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_76 ={ core_csr_decoded_decoded_hi_lo_hi_75 , core_csr_decoded_decoded_andMatrixInput_5_77 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_0_77 , core_csr_decoded_decoded_andMatrixInput_1_77 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_77 ={ core_csr_decoded_decoded_hi_hi_hi_76 , core_csr_decoded_decoded_andMatrixInput_2_77 }; 
    wire[5:0] core_csr_decoded_decoded_hi_77 ={ core_csr_decoded_decoded_hi_hi_77 , core_csr_decoded_decoded_hi_lo_76 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_78 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_78 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_78 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_78 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_78 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_78 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_77 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_77 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_77 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_77 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_76 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_70 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_70 ={ core_csr_decoded_decoded_andMatrixInput_9_77 , core_csr_decoded_decoded_andMatrixInput_10_76 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_77 ={ core_csr_decoded_decoded_lo_lo_hi_70 , core_csr_decoded_decoded_andMatrixInput_11_70 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_6_77 , core_csr_decoded_decoded_andMatrixInput_7_77 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_78 ={ core_csr_decoded_decoded_lo_hi_hi_77 , core_csr_decoded_decoded_andMatrixInput_8_77 }; 
    wire[5:0] core_csr_decoded_decoded_lo_78 ={ core_csr_decoded_decoded_lo_hi_78 , core_csr_decoded_decoded_lo_lo_77 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_3_78 , core_csr_decoded_decoded_andMatrixInput_4_78 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_77 ={ core_csr_decoded_decoded_hi_lo_hi_76 , core_csr_decoded_decoded_andMatrixInput_5_78 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_0_78 , core_csr_decoded_decoded_andMatrixInput_1_78 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_78 ={ core_csr_decoded_decoded_hi_hi_hi_77 , core_csr_decoded_decoded_andMatrixInput_2_78 }; 
    wire[5:0] core_csr_decoded_decoded_hi_78 ={ core_csr_decoded_decoded_hi_hi_78 , core_csr_decoded_decoded_hi_lo_77 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_79 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_79 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_79 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_79 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_79 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_79 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_78 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_78 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_78 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_78 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_77 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_71 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_71 ={ core_csr_decoded_decoded_andMatrixInput_9_78 , core_csr_decoded_decoded_andMatrixInput_10_77 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_78 ={ core_csr_decoded_decoded_lo_lo_hi_71 , core_csr_decoded_decoded_andMatrixInput_11_71 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_6_78 , core_csr_decoded_decoded_andMatrixInput_7_78 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_79 ={ core_csr_decoded_decoded_lo_hi_hi_78 , core_csr_decoded_decoded_andMatrixInput_8_78 }; 
    wire[5:0] core_csr_decoded_decoded_lo_79 ={ core_csr_decoded_decoded_lo_hi_79 , core_csr_decoded_decoded_lo_lo_78 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_3_79 , core_csr_decoded_decoded_andMatrixInput_4_79 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_78 ={ core_csr_decoded_decoded_hi_lo_hi_77 , core_csr_decoded_decoded_andMatrixInput_5_79 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_0_79 , core_csr_decoded_decoded_andMatrixInput_1_79 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_79 ={ core_csr_decoded_decoded_hi_hi_hi_78 , core_csr_decoded_decoded_andMatrixInput_2_79 }; 
    wire[5:0] core_csr_decoded_decoded_hi_79 ={ core_csr_decoded_decoded_hi_hi_79 , core_csr_decoded_decoded_hi_lo_78 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_80 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_80 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_80 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_80 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_80 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_80 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_79 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_79 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_79 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_79 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_78 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_72 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_72 ={ core_csr_decoded_decoded_andMatrixInput_9_79 , core_csr_decoded_decoded_andMatrixInput_10_78 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_79 ={ core_csr_decoded_decoded_lo_lo_hi_72 , core_csr_decoded_decoded_andMatrixInput_11_72 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_6_79 , core_csr_decoded_decoded_andMatrixInput_7_79 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_80 ={ core_csr_decoded_decoded_lo_hi_hi_79 , core_csr_decoded_decoded_andMatrixInput_8_79 }; 
    wire[5:0] core_csr_decoded_decoded_lo_80 ={ core_csr_decoded_decoded_lo_hi_80 , core_csr_decoded_decoded_lo_lo_79 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_3_80 , core_csr_decoded_decoded_andMatrixInput_4_80 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_79 ={ core_csr_decoded_decoded_hi_lo_hi_78 , core_csr_decoded_decoded_andMatrixInput_5_80 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_0_80 , core_csr_decoded_decoded_andMatrixInput_1_80 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_80 ={ core_csr_decoded_decoded_hi_hi_hi_79 , core_csr_decoded_decoded_andMatrixInput_2_80 }; 
    wire[5:0] core_csr_decoded_decoded_hi_80 ={ core_csr_decoded_decoded_hi_hi_80 , core_csr_decoded_decoded_hi_lo_79 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_81 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_81 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_81 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_81 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_81 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_81 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_80 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_80 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_80 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_80 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_79 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_73 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_73 ={ core_csr_decoded_decoded_andMatrixInput_9_80 , core_csr_decoded_decoded_andMatrixInput_10_79 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_80 ={ core_csr_decoded_decoded_lo_lo_hi_73 , core_csr_decoded_decoded_andMatrixInput_11_73 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_6_80 , core_csr_decoded_decoded_andMatrixInput_7_80 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_81 ={ core_csr_decoded_decoded_lo_hi_hi_80 , core_csr_decoded_decoded_andMatrixInput_8_80 }; 
    wire[5:0] core_csr_decoded_decoded_lo_81 ={ core_csr_decoded_decoded_lo_hi_81 , core_csr_decoded_decoded_lo_lo_80 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_3_81 , core_csr_decoded_decoded_andMatrixInput_4_81 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_80 ={ core_csr_decoded_decoded_hi_lo_hi_79 , core_csr_decoded_decoded_andMatrixInput_5_81 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_0_81 , core_csr_decoded_decoded_andMatrixInput_1_81 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_81 ={ core_csr_decoded_decoded_hi_hi_hi_80 , core_csr_decoded_decoded_andMatrixInput_2_81 }; 
    wire[5:0] core_csr_decoded_decoded_hi_81 ={ core_csr_decoded_decoded_hi_hi_81 , core_csr_decoded_decoded_hi_lo_80 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_82 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_82 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_82 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_82 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_82 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_82 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_81 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_81 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_81 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_81 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_80 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_74 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_74 ={ core_csr_decoded_decoded_andMatrixInput_9_81 , core_csr_decoded_decoded_andMatrixInput_10_80 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_81 ={ core_csr_decoded_decoded_lo_lo_hi_74 , core_csr_decoded_decoded_andMatrixInput_11_74 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_6_81 , core_csr_decoded_decoded_andMatrixInput_7_81 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_82 ={ core_csr_decoded_decoded_lo_hi_hi_81 , core_csr_decoded_decoded_andMatrixInput_8_81 }; 
    wire[5:0] core_csr_decoded_decoded_lo_82 ={ core_csr_decoded_decoded_lo_hi_82 , core_csr_decoded_decoded_lo_lo_81 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_3_82 , core_csr_decoded_decoded_andMatrixInput_4_82 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_81 ={ core_csr_decoded_decoded_hi_lo_hi_80 , core_csr_decoded_decoded_andMatrixInput_5_82 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_0_82 , core_csr_decoded_decoded_andMatrixInput_1_82 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_82 ={ core_csr_decoded_decoded_hi_hi_hi_81 , core_csr_decoded_decoded_andMatrixInput_2_82 }; 
    wire[5:0] core_csr_decoded_decoded_hi_82 ={ core_csr_decoded_decoded_hi_hi_82 , core_csr_decoded_decoded_hi_lo_81 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_83 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_83 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_83 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_83 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_83 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_83 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_82 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_82 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_82 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_82 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_81 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_75 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_75 ={ core_csr_decoded_decoded_andMatrixInput_9_82 , core_csr_decoded_decoded_andMatrixInput_10_81 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_82 ={ core_csr_decoded_decoded_lo_lo_hi_75 , core_csr_decoded_decoded_andMatrixInput_11_75 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_6_82 , core_csr_decoded_decoded_andMatrixInput_7_82 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_83 ={ core_csr_decoded_decoded_lo_hi_hi_82 , core_csr_decoded_decoded_andMatrixInput_8_82 }; 
    wire[5:0] core_csr_decoded_decoded_lo_83 ={ core_csr_decoded_decoded_lo_hi_83 , core_csr_decoded_decoded_lo_lo_82 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_3_83 , core_csr_decoded_decoded_andMatrixInput_4_83 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_82 ={ core_csr_decoded_decoded_hi_lo_hi_81 , core_csr_decoded_decoded_andMatrixInput_5_83 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_0_83 , core_csr_decoded_decoded_andMatrixInput_1_83 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_83 ={ core_csr_decoded_decoded_hi_hi_hi_82 , core_csr_decoded_decoded_andMatrixInput_2_83 }; 
    wire[5:0] core_csr_decoded_decoded_hi_83 ={ core_csr_decoded_decoded_hi_hi_83 , core_csr_decoded_decoded_hi_lo_82 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_84 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_84 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_84 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_84 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_84 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_84 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_83 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_83 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_83 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_83 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_82 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_76 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_76 ={ core_csr_decoded_decoded_andMatrixInput_9_83 , core_csr_decoded_decoded_andMatrixInput_10_82 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_83 ={ core_csr_decoded_decoded_lo_lo_hi_76 , core_csr_decoded_decoded_andMatrixInput_11_76 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_6_83 , core_csr_decoded_decoded_andMatrixInput_7_83 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_84 ={ core_csr_decoded_decoded_lo_hi_hi_83 , core_csr_decoded_decoded_andMatrixInput_8_83 }; 
    wire[5:0] core_csr_decoded_decoded_lo_84 ={ core_csr_decoded_decoded_lo_hi_84 , core_csr_decoded_decoded_lo_lo_83 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_3_84 , core_csr_decoded_decoded_andMatrixInput_4_84 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_83 ={ core_csr_decoded_decoded_hi_lo_hi_82 , core_csr_decoded_decoded_andMatrixInput_5_84 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_0_84 , core_csr_decoded_decoded_andMatrixInput_1_84 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_84 ={ core_csr_decoded_decoded_hi_hi_hi_83 , core_csr_decoded_decoded_andMatrixInput_2_84 }; 
    wire[5:0] core_csr_decoded_decoded_hi_84 ={ core_csr_decoded_decoded_hi_hi_84 , core_csr_decoded_decoded_hi_lo_83 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_85 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_85 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_85 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_85 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_85 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_85 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_84 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_84 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_84 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_84 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_83 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_77 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_77 ={ core_csr_decoded_decoded_andMatrixInput_9_84 , core_csr_decoded_decoded_andMatrixInput_10_83 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_84 ={ core_csr_decoded_decoded_lo_lo_hi_77 , core_csr_decoded_decoded_andMatrixInput_11_77 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_6_84 , core_csr_decoded_decoded_andMatrixInput_7_84 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_85 ={ core_csr_decoded_decoded_lo_hi_hi_84 , core_csr_decoded_decoded_andMatrixInput_8_84 }; 
    wire[5:0] core_csr_decoded_decoded_lo_85 ={ core_csr_decoded_decoded_lo_hi_85 , core_csr_decoded_decoded_lo_lo_84 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_3_85 , core_csr_decoded_decoded_andMatrixInput_4_85 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_84 ={ core_csr_decoded_decoded_hi_lo_hi_83 , core_csr_decoded_decoded_andMatrixInput_5_85 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_0_85 , core_csr_decoded_decoded_andMatrixInput_1_85 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_85 ={ core_csr_decoded_decoded_hi_hi_hi_84 , core_csr_decoded_decoded_andMatrixInput_2_85 }; 
    wire[5:0] core_csr_decoded_decoded_hi_85 ={ core_csr_decoded_decoded_hi_hi_85 , core_csr_decoded_decoded_hi_lo_84 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_86 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_86 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_86 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_86 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_86 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_86 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_85 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_85 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_85 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_85 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_84 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_78 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_78 ={ core_csr_decoded_decoded_andMatrixInput_9_85 , core_csr_decoded_decoded_andMatrixInput_10_84 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_85 ={ core_csr_decoded_decoded_lo_lo_hi_78 , core_csr_decoded_decoded_andMatrixInput_11_78 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_6_85 , core_csr_decoded_decoded_andMatrixInput_7_85 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_86 ={ core_csr_decoded_decoded_lo_hi_hi_85 , core_csr_decoded_decoded_andMatrixInput_8_85 }; 
    wire[5:0] core_csr_decoded_decoded_lo_86 ={ core_csr_decoded_decoded_lo_hi_86 , core_csr_decoded_decoded_lo_lo_85 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_3_86 , core_csr_decoded_decoded_andMatrixInput_4_86 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_85 ={ core_csr_decoded_decoded_hi_lo_hi_84 , core_csr_decoded_decoded_andMatrixInput_5_86 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_0_86 , core_csr_decoded_decoded_andMatrixInput_1_86 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_86 ={ core_csr_decoded_decoded_hi_hi_hi_85 , core_csr_decoded_decoded_andMatrixInput_2_86 }; 
    wire[5:0] core_csr_decoded_decoded_hi_86 ={ core_csr_decoded_decoded_hi_hi_86 , core_csr_decoded_decoded_hi_lo_85 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_87 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_87 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_87 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_87 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_87 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_87 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_86 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_86 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_86 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_86 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_85 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_79 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_79 ={ core_csr_decoded_decoded_andMatrixInput_9_86 , core_csr_decoded_decoded_andMatrixInput_10_85 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_86 ={ core_csr_decoded_decoded_lo_lo_hi_79 , core_csr_decoded_decoded_andMatrixInput_11_79 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_6_86 , core_csr_decoded_decoded_andMatrixInput_7_86 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_87 ={ core_csr_decoded_decoded_lo_hi_hi_86 , core_csr_decoded_decoded_andMatrixInput_8_86 }; 
    wire[5:0] core_csr_decoded_decoded_lo_87 ={ core_csr_decoded_decoded_lo_hi_87 , core_csr_decoded_decoded_lo_lo_86 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_3_87 , core_csr_decoded_decoded_andMatrixInput_4_87 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_86 ={ core_csr_decoded_decoded_hi_lo_hi_85 , core_csr_decoded_decoded_andMatrixInput_5_87 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_0_87 , core_csr_decoded_decoded_andMatrixInput_1_87 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_87 ={ core_csr_decoded_decoded_hi_hi_hi_86 , core_csr_decoded_decoded_andMatrixInput_2_87 }; 
    wire[5:0] core_csr_decoded_decoded_hi_87 ={ core_csr_decoded_decoded_hi_hi_87 , core_csr_decoded_decoded_hi_lo_86 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_88 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_88 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_88 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_88 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_88 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_88 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_87 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_87 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_87 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_87 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_86 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_80 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_80 ={ core_csr_decoded_decoded_andMatrixInput_9_87 , core_csr_decoded_decoded_andMatrixInput_10_86 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_87 ={ core_csr_decoded_decoded_lo_lo_hi_80 , core_csr_decoded_decoded_andMatrixInput_11_80 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_6_87 , core_csr_decoded_decoded_andMatrixInput_7_87 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_88 ={ core_csr_decoded_decoded_lo_hi_hi_87 , core_csr_decoded_decoded_andMatrixInput_8_87 }; 
    wire[5:0] core_csr_decoded_decoded_lo_88 ={ core_csr_decoded_decoded_lo_hi_88 , core_csr_decoded_decoded_lo_lo_87 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_3_88 , core_csr_decoded_decoded_andMatrixInput_4_88 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_87 ={ core_csr_decoded_decoded_hi_lo_hi_86 , core_csr_decoded_decoded_andMatrixInput_5_88 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_0_88 , core_csr_decoded_decoded_andMatrixInput_1_88 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_88 ={ core_csr_decoded_decoded_hi_hi_hi_87 , core_csr_decoded_decoded_andMatrixInput_2_88 }; 
    wire[5:0] core_csr_decoded_decoded_hi_88 ={ core_csr_decoded_decoded_hi_hi_88 , core_csr_decoded_decoded_hi_lo_87 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_89 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_89 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_89 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_89 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_89 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_89 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_88 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_88 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_88 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_88 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_87 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_81 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_81 ={ core_csr_decoded_decoded_andMatrixInput_9_88 , core_csr_decoded_decoded_andMatrixInput_10_87 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_88 ={ core_csr_decoded_decoded_lo_lo_hi_81 , core_csr_decoded_decoded_andMatrixInput_11_81 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_6_88 , core_csr_decoded_decoded_andMatrixInput_7_88 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_89 ={ core_csr_decoded_decoded_lo_hi_hi_88 , core_csr_decoded_decoded_andMatrixInput_8_88 }; 
    wire[5:0] core_csr_decoded_decoded_lo_89 ={ core_csr_decoded_decoded_lo_hi_89 , core_csr_decoded_decoded_lo_lo_88 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_3_89 , core_csr_decoded_decoded_andMatrixInput_4_89 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_88 ={ core_csr_decoded_decoded_hi_lo_hi_87 , core_csr_decoded_decoded_andMatrixInput_5_89 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_0_89 , core_csr_decoded_decoded_andMatrixInput_1_89 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_89 ={ core_csr_decoded_decoded_hi_hi_hi_88 , core_csr_decoded_decoded_andMatrixInput_2_89 }; 
    wire[5:0] core_csr_decoded_decoded_hi_89 ={ core_csr_decoded_decoded_hi_hi_89 , core_csr_decoded_decoded_hi_lo_88 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_90 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_90 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_90 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_90 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_90 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_90 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_89 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_89 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_89 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_89 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_88 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_82 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_82 ={ core_csr_decoded_decoded_andMatrixInput_9_89 , core_csr_decoded_decoded_andMatrixInput_10_88 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_89 ={ core_csr_decoded_decoded_lo_lo_hi_82 , core_csr_decoded_decoded_andMatrixInput_11_82 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_6_89 , core_csr_decoded_decoded_andMatrixInput_7_89 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_90 ={ core_csr_decoded_decoded_lo_hi_hi_89 , core_csr_decoded_decoded_andMatrixInput_8_89 }; 
    wire[5:0] core_csr_decoded_decoded_lo_90 ={ core_csr_decoded_decoded_lo_hi_90 , core_csr_decoded_decoded_lo_lo_89 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_3_90 , core_csr_decoded_decoded_andMatrixInput_4_90 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_89 ={ core_csr_decoded_decoded_hi_lo_hi_88 , core_csr_decoded_decoded_andMatrixInput_5_90 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_0_90 , core_csr_decoded_decoded_andMatrixInput_1_90 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_90 ={ core_csr_decoded_decoded_hi_hi_hi_89 , core_csr_decoded_decoded_andMatrixInput_2_90 }; 
    wire[5:0] core_csr_decoded_decoded_hi_90 ={ core_csr_decoded_decoded_hi_hi_90 , core_csr_decoded_decoded_hi_lo_89 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_91 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_91 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_91 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_91 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_91 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_91 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_90 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_90 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_90 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_90 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_89 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_83 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_83 ={ core_csr_decoded_decoded_andMatrixInput_9_90 , core_csr_decoded_decoded_andMatrixInput_10_89 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_90 ={ core_csr_decoded_decoded_lo_lo_hi_83 , core_csr_decoded_decoded_andMatrixInput_11_83 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_6_90 , core_csr_decoded_decoded_andMatrixInput_7_90 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_91 ={ core_csr_decoded_decoded_lo_hi_hi_90 , core_csr_decoded_decoded_andMatrixInput_8_90 }; 
    wire[5:0] core_csr_decoded_decoded_lo_91 ={ core_csr_decoded_decoded_lo_hi_91 , core_csr_decoded_decoded_lo_lo_90 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_3_91 , core_csr_decoded_decoded_andMatrixInput_4_91 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_90 ={ core_csr_decoded_decoded_hi_lo_hi_89 , core_csr_decoded_decoded_andMatrixInput_5_91 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_0_91 , core_csr_decoded_decoded_andMatrixInput_1_91 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_91 ={ core_csr_decoded_decoded_hi_hi_hi_90 , core_csr_decoded_decoded_andMatrixInput_2_91 }; 
    wire[5:0] core_csr_decoded_decoded_hi_91 ={ core_csr_decoded_decoded_hi_hi_91 , core_csr_decoded_decoded_hi_lo_90 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_92 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_92 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_92 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_92 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_92 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_92 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_91 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_91 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_91 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_91 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_90 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_84 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_84 ={ core_csr_decoded_decoded_andMatrixInput_9_91 , core_csr_decoded_decoded_andMatrixInput_10_90 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_91 ={ core_csr_decoded_decoded_lo_lo_hi_84 , core_csr_decoded_decoded_andMatrixInput_11_84 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_6_91 , core_csr_decoded_decoded_andMatrixInput_7_91 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_92 ={ core_csr_decoded_decoded_lo_hi_hi_91 , core_csr_decoded_decoded_andMatrixInput_8_91 }; 
    wire[5:0] core_csr_decoded_decoded_lo_92 ={ core_csr_decoded_decoded_lo_hi_92 , core_csr_decoded_decoded_lo_lo_91 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_3_92 , core_csr_decoded_decoded_andMatrixInput_4_92 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_91 ={ core_csr_decoded_decoded_hi_lo_hi_90 , core_csr_decoded_decoded_andMatrixInput_5_92 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_0_92 , core_csr_decoded_decoded_andMatrixInput_1_92 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_92 ={ core_csr_decoded_decoded_hi_hi_hi_91 , core_csr_decoded_decoded_andMatrixInput_2_92 }; 
    wire[5:0] core_csr_decoded_decoded_hi_92 ={ core_csr_decoded_decoded_hi_hi_92 , core_csr_decoded_decoded_hi_lo_91 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_93 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_93 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_93 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_93 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_93 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_93 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_92 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_92 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_92 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_92 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_91 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_85 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_85 ={ core_csr_decoded_decoded_andMatrixInput_9_92 , core_csr_decoded_decoded_andMatrixInput_10_91 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_92 ={ core_csr_decoded_decoded_lo_lo_hi_85 , core_csr_decoded_decoded_andMatrixInput_11_85 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_6_92 , core_csr_decoded_decoded_andMatrixInput_7_92 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_93 ={ core_csr_decoded_decoded_lo_hi_hi_92 , core_csr_decoded_decoded_andMatrixInput_8_92 }; 
    wire[5:0] core_csr_decoded_decoded_lo_93 ={ core_csr_decoded_decoded_lo_hi_93 , core_csr_decoded_decoded_lo_lo_92 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_3_93 , core_csr_decoded_decoded_andMatrixInput_4_93 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_92 ={ core_csr_decoded_decoded_hi_lo_hi_91 , core_csr_decoded_decoded_andMatrixInput_5_93 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_0_93 , core_csr_decoded_decoded_andMatrixInput_1_93 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_93 ={ core_csr_decoded_decoded_hi_hi_hi_92 , core_csr_decoded_decoded_andMatrixInput_2_93 }; 
    wire[5:0] core_csr_decoded_decoded_hi_93 ={ core_csr_decoded_decoded_hi_hi_93 , core_csr_decoded_decoded_hi_lo_92 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_94 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_94 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_94 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_94 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_94 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_94 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_93 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_93 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_93 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_93 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_92 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_86 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_86 ={ core_csr_decoded_decoded_andMatrixInput_9_93 , core_csr_decoded_decoded_andMatrixInput_10_92 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_93 ={ core_csr_decoded_decoded_lo_lo_hi_86 , core_csr_decoded_decoded_andMatrixInput_11_86 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_6_93 , core_csr_decoded_decoded_andMatrixInput_7_93 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_94 ={ core_csr_decoded_decoded_lo_hi_hi_93 , core_csr_decoded_decoded_andMatrixInput_8_93 }; 
    wire[5:0] core_csr_decoded_decoded_lo_94 ={ core_csr_decoded_decoded_lo_hi_94 , core_csr_decoded_decoded_lo_lo_93 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_3_94 , core_csr_decoded_decoded_andMatrixInput_4_94 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_93 ={ core_csr_decoded_decoded_hi_lo_hi_92 , core_csr_decoded_decoded_andMatrixInput_5_94 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_0_94 , core_csr_decoded_decoded_andMatrixInput_1_94 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_94 ={ core_csr_decoded_decoded_hi_hi_hi_93 , core_csr_decoded_decoded_andMatrixInput_2_94 }; 
    wire[5:0] core_csr_decoded_decoded_hi_94 ={ core_csr_decoded_decoded_hi_hi_94 , core_csr_decoded_decoded_hi_lo_93 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_95 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_95 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_95 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_95 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_95 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_95 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_94 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_94 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_94 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_94 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_93 = core_csr_decoded_decoded_invInputs [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_87 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_87 ={ core_csr_decoded_decoded_andMatrixInput_9_94 , core_csr_decoded_decoded_andMatrixInput_10_93 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_94 ={ core_csr_decoded_decoded_lo_lo_hi_87 , core_csr_decoded_decoded_andMatrixInput_11_87 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_6_94 , core_csr_decoded_decoded_andMatrixInput_7_94 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_95 ={ core_csr_decoded_decoded_lo_hi_hi_94 , core_csr_decoded_decoded_andMatrixInput_8_94 }; 
    wire[5:0] core_csr_decoded_decoded_lo_95 ={ core_csr_decoded_decoded_lo_hi_95 , core_csr_decoded_decoded_lo_lo_94 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_3_95 , core_csr_decoded_decoded_andMatrixInput_4_95 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_94 ={ core_csr_decoded_decoded_hi_lo_hi_93 , core_csr_decoded_decoded_andMatrixInput_5_95 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_0_95 , core_csr_decoded_decoded_andMatrixInput_1_95 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_95 ={ core_csr_decoded_decoded_hi_hi_hi_94 , core_csr_decoded_decoded_andMatrixInput_2_95 }; 
    wire[5:0] core_csr_decoded_decoded_hi_95 ={ core_csr_decoded_decoded_hi_hi_95 , core_csr_decoded_decoded_hi_lo_94 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_96 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_96 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_96 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_96 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_96 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_96 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_95 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_95 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_95 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_95 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_94 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_95 ={ core_csr_decoded_decoded_andMatrixInput_9_95 , core_csr_decoded_decoded_andMatrixInput_10_94 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_6_95 , core_csr_decoded_decoded_andMatrixInput_7_95 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_96 ={ core_csr_decoded_decoded_lo_hi_hi_95 , core_csr_decoded_decoded_andMatrixInput_8_95 }; 
    wire[4:0] core_csr_decoded_decoded_lo_96 ={ core_csr_decoded_decoded_lo_hi_96 , core_csr_decoded_decoded_lo_lo_95 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_3_96 , core_csr_decoded_decoded_andMatrixInput_4_96 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_95 ={ core_csr_decoded_decoded_hi_lo_hi_94 , core_csr_decoded_decoded_andMatrixInput_5_96 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_0_96 , core_csr_decoded_decoded_andMatrixInput_1_96 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_96 ={ core_csr_decoded_decoded_hi_hi_hi_95 , core_csr_decoded_decoded_andMatrixInput_2_96 }; 
    wire[5:0] core_csr_decoded_decoded_hi_96 ={ core_csr_decoded_decoded_hi_hi_96 , core_csr_decoded_decoded_hi_lo_95 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_97 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_97 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_97 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_97 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_97 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_97 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_96 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_96 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_96 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_96 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_95 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_88 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_88 ={ core_csr_decoded_decoded_andMatrixInput_9_96 , core_csr_decoded_decoded_andMatrixInput_10_95 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_96 ={ core_csr_decoded_decoded_lo_lo_hi_88 , core_csr_decoded_decoded_andMatrixInput_11_88 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_6_96 , core_csr_decoded_decoded_andMatrixInput_7_96 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_97 ={ core_csr_decoded_decoded_lo_hi_hi_96 , core_csr_decoded_decoded_andMatrixInput_8_96 }; 
    wire[5:0] core_csr_decoded_decoded_lo_97 ={ core_csr_decoded_decoded_lo_hi_97 , core_csr_decoded_decoded_lo_lo_96 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_3_97 , core_csr_decoded_decoded_andMatrixInput_4_97 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_96 ={ core_csr_decoded_decoded_hi_lo_hi_95 , core_csr_decoded_decoded_andMatrixInput_5_97 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_0_97 , core_csr_decoded_decoded_andMatrixInput_1_97 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_97 ={ core_csr_decoded_decoded_hi_hi_hi_96 , core_csr_decoded_decoded_andMatrixInput_2_97 }; 
    wire[5:0] core_csr_decoded_decoded_hi_97 ={ core_csr_decoded_decoded_hi_hi_97 , core_csr_decoded_decoded_hi_lo_96 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_98 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_98 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_98 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_98 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_98 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_98 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_97 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_97 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_97 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_97 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_96 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_89 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_89 ={ core_csr_decoded_decoded_andMatrixInput_9_97 , core_csr_decoded_decoded_andMatrixInput_10_96 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_97 ={ core_csr_decoded_decoded_lo_lo_hi_89 , core_csr_decoded_decoded_andMatrixInput_11_89 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_6_97 , core_csr_decoded_decoded_andMatrixInput_7_97 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_98 ={ core_csr_decoded_decoded_lo_hi_hi_97 , core_csr_decoded_decoded_andMatrixInput_8_97 }; 
    wire[5:0] core_csr_decoded_decoded_lo_98 ={ core_csr_decoded_decoded_lo_hi_98 , core_csr_decoded_decoded_lo_lo_97 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_3_98 , core_csr_decoded_decoded_andMatrixInput_4_98 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_97 ={ core_csr_decoded_decoded_hi_lo_hi_96 , core_csr_decoded_decoded_andMatrixInput_5_98 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_0_98 , core_csr_decoded_decoded_andMatrixInput_1_98 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_98 ={ core_csr_decoded_decoded_hi_hi_hi_97 , core_csr_decoded_decoded_andMatrixInput_2_98 }; 
    wire[5:0] core_csr_decoded_decoded_hi_98 ={ core_csr_decoded_decoded_hi_hi_98 , core_csr_decoded_decoded_hi_lo_97 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_99 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_99 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_99 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_99 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_99 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_99 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_98 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_98 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_98 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_98 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_97 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_90 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_90 ={ core_csr_decoded_decoded_andMatrixInput_9_98 , core_csr_decoded_decoded_andMatrixInput_10_97 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_98 ={ core_csr_decoded_decoded_lo_lo_hi_90 , core_csr_decoded_decoded_andMatrixInput_11_90 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_6_98 , core_csr_decoded_decoded_andMatrixInput_7_98 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_99 ={ core_csr_decoded_decoded_lo_hi_hi_98 , core_csr_decoded_decoded_andMatrixInput_8_98 }; 
    wire[5:0] core_csr_decoded_decoded_lo_99 ={ core_csr_decoded_decoded_lo_hi_99 , core_csr_decoded_decoded_lo_lo_98 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_3_99 , core_csr_decoded_decoded_andMatrixInput_4_99 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_98 ={ core_csr_decoded_decoded_hi_lo_hi_97 , core_csr_decoded_decoded_andMatrixInput_5_99 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_0_99 , core_csr_decoded_decoded_andMatrixInput_1_99 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_99 ={ core_csr_decoded_decoded_hi_hi_hi_98 , core_csr_decoded_decoded_andMatrixInput_2_99 }; 
    wire[5:0] core_csr_decoded_decoded_hi_99 ={ core_csr_decoded_decoded_hi_hi_99 , core_csr_decoded_decoded_hi_lo_98 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_100 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_100 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_100 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_100 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_100 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_100 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_99 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_99 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_99 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_99 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_98 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_91 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_91 ={ core_csr_decoded_decoded_andMatrixInput_9_99 , core_csr_decoded_decoded_andMatrixInput_10_98 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_99 ={ core_csr_decoded_decoded_lo_lo_hi_91 , core_csr_decoded_decoded_andMatrixInput_11_91 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_6_99 , core_csr_decoded_decoded_andMatrixInput_7_99 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_100 ={ core_csr_decoded_decoded_lo_hi_hi_99 , core_csr_decoded_decoded_andMatrixInput_8_99 }; 
    wire[5:0] core_csr_decoded_decoded_lo_100 ={ core_csr_decoded_decoded_lo_hi_100 , core_csr_decoded_decoded_lo_lo_99 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_3_100 , core_csr_decoded_decoded_andMatrixInput_4_100 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_99 ={ core_csr_decoded_decoded_hi_lo_hi_98 , core_csr_decoded_decoded_andMatrixInput_5_100 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_0_100 , core_csr_decoded_decoded_andMatrixInput_1_100 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_100 ={ core_csr_decoded_decoded_hi_hi_hi_99 , core_csr_decoded_decoded_andMatrixInput_2_100 }; 
    wire[5:0] core_csr_decoded_decoded_hi_100 ={ core_csr_decoded_decoded_hi_hi_100 , core_csr_decoded_decoded_hi_lo_99 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_101 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_101 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_101 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_101 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_101 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_101 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_100 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_100 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_100 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_100 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_99 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_92 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_92 ={ core_csr_decoded_decoded_andMatrixInput_9_100 , core_csr_decoded_decoded_andMatrixInput_10_99 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_100 ={ core_csr_decoded_decoded_lo_lo_hi_92 , core_csr_decoded_decoded_andMatrixInput_11_92 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_6_100 , core_csr_decoded_decoded_andMatrixInput_7_100 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_101 ={ core_csr_decoded_decoded_lo_hi_hi_100 , core_csr_decoded_decoded_andMatrixInput_8_100 }; 
    wire[5:0] core_csr_decoded_decoded_lo_101 ={ core_csr_decoded_decoded_lo_hi_101 , core_csr_decoded_decoded_lo_lo_100 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_3_101 , core_csr_decoded_decoded_andMatrixInput_4_101 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_100 ={ core_csr_decoded_decoded_hi_lo_hi_99 , core_csr_decoded_decoded_andMatrixInput_5_101 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_0_101 , core_csr_decoded_decoded_andMatrixInput_1_101 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_101 ={ core_csr_decoded_decoded_hi_hi_hi_100 , core_csr_decoded_decoded_andMatrixInput_2_101 }; 
    wire[5:0] core_csr_decoded_decoded_hi_101 ={ core_csr_decoded_decoded_hi_hi_101 , core_csr_decoded_decoded_hi_lo_100 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_102 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_102 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_102 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_102 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_102 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_102 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_101 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_101 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_101 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_101 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_100 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_93 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_93 ={ core_csr_decoded_decoded_andMatrixInput_9_101 , core_csr_decoded_decoded_andMatrixInput_10_100 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_101 ={ core_csr_decoded_decoded_lo_lo_hi_93 , core_csr_decoded_decoded_andMatrixInput_11_93 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_6_101 , core_csr_decoded_decoded_andMatrixInput_7_101 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_102 ={ core_csr_decoded_decoded_lo_hi_hi_101 , core_csr_decoded_decoded_andMatrixInput_8_101 }; 
    wire[5:0] core_csr_decoded_decoded_lo_102 ={ core_csr_decoded_decoded_lo_hi_102 , core_csr_decoded_decoded_lo_lo_101 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_3_102 , core_csr_decoded_decoded_andMatrixInput_4_102 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_101 ={ core_csr_decoded_decoded_hi_lo_hi_100 , core_csr_decoded_decoded_andMatrixInput_5_102 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_0_102 , core_csr_decoded_decoded_andMatrixInput_1_102 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_102 ={ core_csr_decoded_decoded_hi_hi_hi_101 , core_csr_decoded_decoded_andMatrixInput_2_102 }; 
    wire[5:0] core_csr_decoded_decoded_hi_102 ={ core_csr_decoded_decoded_hi_hi_102 , core_csr_decoded_decoded_hi_lo_101 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_103 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_103 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_103 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_103 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_103 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_103 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_102 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_102 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_102 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_102 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_101 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_94 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_94 ={ core_csr_decoded_decoded_andMatrixInput_9_102 , core_csr_decoded_decoded_andMatrixInput_10_101 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_102 ={ core_csr_decoded_decoded_lo_lo_hi_94 , core_csr_decoded_decoded_andMatrixInput_11_94 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_6_102 , core_csr_decoded_decoded_andMatrixInput_7_102 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_103 ={ core_csr_decoded_decoded_lo_hi_hi_102 , core_csr_decoded_decoded_andMatrixInput_8_102 }; 
    wire[5:0] core_csr_decoded_decoded_lo_103 ={ core_csr_decoded_decoded_lo_hi_103 , core_csr_decoded_decoded_lo_lo_102 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_3_103 , core_csr_decoded_decoded_andMatrixInput_4_103 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_102 ={ core_csr_decoded_decoded_hi_lo_hi_101 , core_csr_decoded_decoded_andMatrixInput_5_103 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_0_103 , core_csr_decoded_decoded_andMatrixInput_1_103 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_103 ={ core_csr_decoded_decoded_hi_hi_hi_102 , core_csr_decoded_decoded_andMatrixInput_2_103 }; 
    wire[5:0] core_csr_decoded_decoded_hi_103 ={ core_csr_decoded_decoded_hi_hi_103 , core_csr_decoded_decoded_hi_lo_102 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_104 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_104 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_104 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_104 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_104 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_104 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_103 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_103 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_103 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_103 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_102 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_95 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_95 ={ core_csr_decoded_decoded_andMatrixInput_9_103 , core_csr_decoded_decoded_andMatrixInput_10_102 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_103 ={ core_csr_decoded_decoded_lo_lo_hi_95 , core_csr_decoded_decoded_andMatrixInput_11_95 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_6_103 , core_csr_decoded_decoded_andMatrixInput_7_103 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_104 ={ core_csr_decoded_decoded_lo_hi_hi_103 , core_csr_decoded_decoded_andMatrixInput_8_103 }; 
    wire[5:0] core_csr_decoded_decoded_lo_104 ={ core_csr_decoded_decoded_lo_hi_104 , core_csr_decoded_decoded_lo_lo_103 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_3_104 , core_csr_decoded_decoded_andMatrixInput_4_104 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_103 ={ core_csr_decoded_decoded_hi_lo_hi_102 , core_csr_decoded_decoded_andMatrixInput_5_104 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_0_104 , core_csr_decoded_decoded_andMatrixInput_1_104 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_104 ={ core_csr_decoded_decoded_hi_hi_hi_103 , core_csr_decoded_decoded_andMatrixInput_2_104 }; 
    wire[5:0] core_csr_decoded_decoded_hi_104 ={ core_csr_decoded_decoded_hi_hi_104 , core_csr_decoded_decoded_hi_lo_103 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_105 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_105 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_105 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_105 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_105 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_105 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_104 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_104 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_104 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_104 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_103 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_96 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_96 ={ core_csr_decoded_decoded_andMatrixInput_9_104 , core_csr_decoded_decoded_andMatrixInput_10_103 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_104 ={ core_csr_decoded_decoded_lo_lo_hi_96 , core_csr_decoded_decoded_andMatrixInput_11_96 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_6_104 , core_csr_decoded_decoded_andMatrixInput_7_104 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_105 ={ core_csr_decoded_decoded_lo_hi_hi_104 , core_csr_decoded_decoded_andMatrixInput_8_104 }; 
    wire[5:0] core_csr_decoded_decoded_lo_105 ={ core_csr_decoded_decoded_lo_hi_105 , core_csr_decoded_decoded_lo_lo_104 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_3_105 , core_csr_decoded_decoded_andMatrixInput_4_105 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_104 ={ core_csr_decoded_decoded_hi_lo_hi_103 , core_csr_decoded_decoded_andMatrixInput_5_105 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_0_105 , core_csr_decoded_decoded_andMatrixInput_1_105 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_105 ={ core_csr_decoded_decoded_hi_hi_hi_104 , core_csr_decoded_decoded_andMatrixInput_2_105 }; 
    wire[5:0] core_csr_decoded_decoded_hi_105 ={ core_csr_decoded_decoded_hi_hi_105 , core_csr_decoded_decoded_hi_lo_104 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_106 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_106 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_106 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_106 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_106 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_106 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_105 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_105 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_105 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_105 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_104 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_97 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_97 ={ core_csr_decoded_decoded_andMatrixInput_9_105 , core_csr_decoded_decoded_andMatrixInput_10_104 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_105 ={ core_csr_decoded_decoded_lo_lo_hi_97 , core_csr_decoded_decoded_andMatrixInput_11_97 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_6_105 , core_csr_decoded_decoded_andMatrixInput_7_105 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_106 ={ core_csr_decoded_decoded_lo_hi_hi_105 , core_csr_decoded_decoded_andMatrixInput_8_105 }; 
    wire[5:0] core_csr_decoded_decoded_lo_106 ={ core_csr_decoded_decoded_lo_hi_106 , core_csr_decoded_decoded_lo_lo_105 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_3_106 , core_csr_decoded_decoded_andMatrixInput_4_106 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_105 ={ core_csr_decoded_decoded_hi_lo_hi_104 , core_csr_decoded_decoded_andMatrixInput_5_106 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_0_106 , core_csr_decoded_decoded_andMatrixInput_1_106 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_106 ={ core_csr_decoded_decoded_hi_hi_hi_105 , core_csr_decoded_decoded_andMatrixInput_2_106 }; 
    wire[5:0] core_csr_decoded_decoded_hi_106 ={ core_csr_decoded_decoded_hi_hi_106 , core_csr_decoded_decoded_hi_lo_105 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_107 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_107 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_107 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_107 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_107 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_107 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_106 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_106 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_106 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_106 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_105 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_98 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_98 ={ core_csr_decoded_decoded_andMatrixInput_9_106 , core_csr_decoded_decoded_andMatrixInput_10_105 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_106 ={ core_csr_decoded_decoded_lo_lo_hi_98 , core_csr_decoded_decoded_andMatrixInput_11_98 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_6_106 , core_csr_decoded_decoded_andMatrixInput_7_106 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_107 ={ core_csr_decoded_decoded_lo_hi_hi_106 , core_csr_decoded_decoded_andMatrixInput_8_106 }; 
    wire[5:0] core_csr_decoded_decoded_lo_107 ={ core_csr_decoded_decoded_lo_hi_107 , core_csr_decoded_decoded_lo_lo_106 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_3_107 , core_csr_decoded_decoded_andMatrixInput_4_107 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_106 ={ core_csr_decoded_decoded_hi_lo_hi_105 , core_csr_decoded_decoded_andMatrixInput_5_107 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_0_107 , core_csr_decoded_decoded_andMatrixInput_1_107 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_107 ={ core_csr_decoded_decoded_hi_hi_hi_106 , core_csr_decoded_decoded_andMatrixInput_2_107 }; 
    wire[5:0] core_csr_decoded_decoded_hi_107 ={ core_csr_decoded_decoded_hi_hi_107 , core_csr_decoded_decoded_hi_lo_106 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_108 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_108 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_108 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_108 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_108 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_108 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_107 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_107 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_107 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_107 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_106 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_99 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_99 ={ core_csr_decoded_decoded_andMatrixInput_9_107 , core_csr_decoded_decoded_andMatrixInput_10_106 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_107 ={ core_csr_decoded_decoded_lo_lo_hi_99 , core_csr_decoded_decoded_andMatrixInput_11_99 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_6_107 , core_csr_decoded_decoded_andMatrixInput_7_107 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_108 ={ core_csr_decoded_decoded_lo_hi_hi_107 , core_csr_decoded_decoded_andMatrixInput_8_107 }; 
    wire[5:0] core_csr_decoded_decoded_lo_108 ={ core_csr_decoded_decoded_lo_hi_108 , core_csr_decoded_decoded_lo_lo_107 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_3_108 , core_csr_decoded_decoded_andMatrixInput_4_108 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_107 ={ core_csr_decoded_decoded_hi_lo_hi_106 , core_csr_decoded_decoded_andMatrixInput_5_108 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_0_108 , core_csr_decoded_decoded_andMatrixInput_1_108 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_108 ={ core_csr_decoded_decoded_hi_hi_hi_107 , core_csr_decoded_decoded_andMatrixInput_2_108 }; 
    wire[5:0] core_csr_decoded_decoded_hi_108 ={ core_csr_decoded_decoded_hi_hi_108 , core_csr_decoded_decoded_hi_lo_107 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_109 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_109 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_109 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_109 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_109 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_109 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_108 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_108 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_108 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_108 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_107 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_100 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_100 ={ core_csr_decoded_decoded_andMatrixInput_9_108 , core_csr_decoded_decoded_andMatrixInput_10_107 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_108 ={ core_csr_decoded_decoded_lo_lo_hi_100 , core_csr_decoded_decoded_andMatrixInput_11_100 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_6_108 , core_csr_decoded_decoded_andMatrixInput_7_108 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_109 ={ core_csr_decoded_decoded_lo_hi_hi_108 , core_csr_decoded_decoded_andMatrixInput_8_108 }; 
    wire[5:0] core_csr_decoded_decoded_lo_109 ={ core_csr_decoded_decoded_lo_hi_109 , core_csr_decoded_decoded_lo_lo_108 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_3_109 , core_csr_decoded_decoded_andMatrixInput_4_109 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_108 ={ core_csr_decoded_decoded_hi_lo_hi_107 , core_csr_decoded_decoded_andMatrixInput_5_109 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_0_109 , core_csr_decoded_decoded_andMatrixInput_1_109 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_109 ={ core_csr_decoded_decoded_hi_hi_hi_108 , core_csr_decoded_decoded_andMatrixInput_2_109 }; 
    wire[5:0] core_csr_decoded_decoded_hi_109 ={ core_csr_decoded_decoded_hi_hi_109 , core_csr_decoded_decoded_hi_lo_108 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_110 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_110 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_110 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_110 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_110 = core_csr_decoded_decoded_invInputs [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_110 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_109 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_109 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_109 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_109 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_108 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_101 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_101 ={ core_csr_decoded_decoded_andMatrixInput_9_109 , core_csr_decoded_decoded_andMatrixInput_10_108 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_109 ={ core_csr_decoded_decoded_lo_lo_hi_101 , core_csr_decoded_decoded_andMatrixInput_11_101 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_6_109 , core_csr_decoded_decoded_andMatrixInput_7_109 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_110 ={ core_csr_decoded_decoded_lo_hi_hi_109 , core_csr_decoded_decoded_andMatrixInput_8_109 }; 
    wire[5:0] core_csr_decoded_decoded_lo_110 ={ core_csr_decoded_decoded_lo_hi_110 , core_csr_decoded_decoded_lo_lo_109 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_3_110 , core_csr_decoded_decoded_andMatrixInput_4_110 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_109 ={ core_csr_decoded_decoded_hi_lo_hi_108 , core_csr_decoded_decoded_andMatrixInput_5_110 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_0_110 , core_csr_decoded_decoded_andMatrixInput_1_110 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_110 ={ core_csr_decoded_decoded_hi_hi_hi_109 , core_csr_decoded_decoded_andMatrixInput_2_110 }; 
    wire[5:0] core_csr_decoded_decoded_hi_110 ={ core_csr_decoded_decoded_hi_hi_110 , core_csr_decoded_decoded_hi_lo_109 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_111 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_111 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_111 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_111 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_111 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_111 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_110 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_110 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_110 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_110 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_109 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_102 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_102 ={ core_csr_decoded_decoded_andMatrixInput_9_110 , core_csr_decoded_decoded_andMatrixInput_10_109 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_110 ={ core_csr_decoded_decoded_lo_lo_hi_102 , core_csr_decoded_decoded_andMatrixInput_11_102 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_6_110 , core_csr_decoded_decoded_andMatrixInput_7_110 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_111 ={ core_csr_decoded_decoded_lo_hi_hi_110 , core_csr_decoded_decoded_andMatrixInput_8_110 }; 
    wire[5:0] core_csr_decoded_decoded_lo_111 ={ core_csr_decoded_decoded_lo_hi_111 , core_csr_decoded_decoded_lo_lo_110 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_3_111 , core_csr_decoded_decoded_andMatrixInput_4_111 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_110 ={ core_csr_decoded_decoded_hi_lo_hi_109 , core_csr_decoded_decoded_andMatrixInput_5_111 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_0_111 , core_csr_decoded_decoded_andMatrixInput_1_111 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_111 ={ core_csr_decoded_decoded_hi_hi_hi_110 , core_csr_decoded_decoded_andMatrixInput_2_111 }; 
    wire[5:0] core_csr_decoded_decoded_hi_111 ={ core_csr_decoded_decoded_hi_hi_111 , core_csr_decoded_decoded_hi_lo_110 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_112 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_112 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_112 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_112 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_112 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_112 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_111 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_111 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_111 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_111 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_110 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_103 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_103 ={ core_csr_decoded_decoded_andMatrixInput_9_111 , core_csr_decoded_decoded_andMatrixInput_10_110 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_111 ={ core_csr_decoded_decoded_lo_lo_hi_103 , core_csr_decoded_decoded_andMatrixInput_11_103 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_6_111 , core_csr_decoded_decoded_andMatrixInput_7_111 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_112 ={ core_csr_decoded_decoded_lo_hi_hi_111 , core_csr_decoded_decoded_andMatrixInput_8_111 }; 
    wire[5:0] core_csr_decoded_decoded_lo_112 ={ core_csr_decoded_decoded_lo_hi_112 , core_csr_decoded_decoded_lo_lo_111 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_3_112 , core_csr_decoded_decoded_andMatrixInput_4_112 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_111 ={ core_csr_decoded_decoded_hi_lo_hi_110 , core_csr_decoded_decoded_andMatrixInput_5_112 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_0_112 , core_csr_decoded_decoded_andMatrixInput_1_112 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_112 ={ core_csr_decoded_decoded_hi_hi_hi_111 , core_csr_decoded_decoded_andMatrixInput_2_112 }; 
    wire[5:0] core_csr_decoded_decoded_hi_112 ={ core_csr_decoded_decoded_hi_hi_112 , core_csr_decoded_decoded_hi_lo_111 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_113 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_113 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_113 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_113 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_113 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_113 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_112 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_112 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_112 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_112 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_111 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_104 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_104 ={ core_csr_decoded_decoded_andMatrixInput_9_112 , core_csr_decoded_decoded_andMatrixInput_10_111 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_112 ={ core_csr_decoded_decoded_lo_lo_hi_104 , core_csr_decoded_decoded_andMatrixInput_11_104 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_6_112 , core_csr_decoded_decoded_andMatrixInput_7_112 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_113 ={ core_csr_decoded_decoded_lo_hi_hi_112 , core_csr_decoded_decoded_andMatrixInput_8_112 }; 
    wire[5:0] core_csr_decoded_decoded_lo_113 ={ core_csr_decoded_decoded_lo_hi_113 , core_csr_decoded_decoded_lo_lo_112 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_3_113 , core_csr_decoded_decoded_andMatrixInput_4_113 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_112 ={ core_csr_decoded_decoded_hi_lo_hi_111 , core_csr_decoded_decoded_andMatrixInput_5_113 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_0_113 , core_csr_decoded_decoded_andMatrixInput_1_113 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_113 ={ core_csr_decoded_decoded_hi_hi_hi_112 , core_csr_decoded_decoded_andMatrixInput_2_113 }; 
    wire[5:0] core_csr_decoded_decoded_hi_113 ={ core_csr_decoded_decoded_hi_hi_113 , core_csr_decoded_decoded_hi_lo_112 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_114 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_114 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_114 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_114 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_114 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_114 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_113 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_113 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_113 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_113 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_112 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_105 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_105 ={ core_csr_decoded_decoded_andMatrixInput_9_113 , core_csr_decoded_decoded_andMatrixInput_10_112 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_113 ={ core_csr_decoded_decoded_lo_lo_hi_105 , core_csr_decoded_decoded_andMatrixInput_11_105 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_6_113 , core_csr_decoded_decoded_andMatrixInput_7_113 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_114 ={ core_csr_decoded_decoded_lo_hi_hi_113 , core_csr_decoded_decoded_andMatrixInput_8_113 }; 
    wire[5:0] core_csr_decoded_decoded_lo_114 ={ core_csr_decoded_decoded_lo_hi_114 , core_csr_decoded_decoded_lo_lo_113 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_3_114 , core_csr_decoded_decoded_andMatrixInput_4_114 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_113 ={ core_csr_decoded_decoded_hi_lo_hi_112 , core_csr_decoded_decoded_andMatrixInput_5_114 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_0_114 , core_csr_decoded_decoded_andMatrixInput_1_114 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_114 ={ core_csr_decoded_decoded_hi_hi_hi_113 , core_csr_decoded_decoded_andMatrixInput_2_114 }; 
    wire[5:0] core_csr_decoded_decoded_hi_114 ={ core_csr_decoded_decoded_hi_hi_114 , core_csr_decoded_decoded_hi_lo_113 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_115 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_115 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_115 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_115 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_115 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_115 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_114 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_114 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_114 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_114 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_113 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_106 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_106 ={ core_csr_decoded_decoded_andMatrixInput_9_114 , core_csr_decoded_decoded_andMatrixInput_10_113 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_114 ={ core_csr_decoded_decoded_lo_lo_hi_106 , core_csr_decoded_decoded_andMatrixInput_11_106 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_6_114 , core_csr_decoded_decoded_andMatrixInput_7_114 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_115 ={ core_csr_decoded_decoded_lo_hi_hi_114 , core_csr_decoded_decoded_andMatrixInput_8_114 }; 
    wire[5:0] core_csr_decoded_decoded_lo_115 ={ core_csr_decoded_decoded_lo_hi_115 , core_csr_decoded_decoded_lo_lo_114 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_3_115 , core_csr_decoded_decoded_andMatrixInput_4_115 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_114 ={ core_csr_decoded_decoded_hi_lo_hi_113 , core_csr_decoded_decoded_andMatrixInput_5_115 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_0_115 , core_csr_decoded_decoded_andMatrixInput_1_115 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_115 ={ core_csr_decoded_decoded_hi_hi_hi_114 , core_csr_decoded_decoded_andMatrixInput_2_115 }; 
    wire[5:0] core_csr_decoded_decoded_hi_115 ={ core_csr_decoded_decoded_hi_hi_115 , core_csr_decoded_decoded_hi_lo_114 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_116 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_116 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_116 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_116 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_116 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_116 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_115 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_115 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_115 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_115 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_114 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_107 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_107 ={ core_csr_decoded_decoded_andMatrixInput_9_115 , core_csr_decoded_decoded_andMatrixInput_10_114 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_115 ={ core_csr_decoded_decoded_lo_lo_hi_107 , core_csr_decoded_decoded_andMatrixInput_11_107 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_6_115 , core_csr_decoded_decoded_andMatrixInput_7_115 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_116 ={ core_csr_decoded_decoded_lo_hi_hi_115 , core_csr_decoded_decoded_andMatrixInput_8_115 }; 
    wire[5:0] core_csr_decoded_decoded_lo_116 ={ core_csr_decoded_decoded_lo_hi_116 , core_csr_decoded_decoded_lo_lo_115 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_3_116 , core_csr_decoded_decoded_andMatrixInput_4_116 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_115 ={ core_csr_decoded_decoded_hi_lo_hi_114 , core_csr_decoded_decoded_andMatrixInput_5_116 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_0_116 , core_csr_decoded_decoded_andMatrixInput_1_116 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_116 ={ core_csr_decoded_decoded_hi_hi_hi_115 , core_csr_decoded_decoded_andMatrixInput_2_116 }; 
    wire[5:0] core_csr_decoded_decoded_hi_116 ={ core_csr_decoded_decoded_hi_hi_116 , core_csr_decoded_decoded_hi_lo_115 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_117 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_117 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_117 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_117 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_117 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_117 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_116 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_116 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_116 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_116 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_115 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_108 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_108 ={ core_csr_decoded_decoded_andMatrixInput_9_116 , core_csr_decoded_decoded_andMatrixInput_10_115 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_116 ={ core_csr_decoded_decoded_lo_lo_hi_108 , core_csr_decoded_decoded_andMatrixInput_11_108 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_6_116 , core_csr_decoded_decoded_andMatrixInput_7_116 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_117 ={ core_csr_decoded_decoded_lo_hi_hi_116 , core_csr_decoded_decoded_andMatrixInput_8_116 }; 
    wire[5:0] core_csr_decoded_decoded_lo_117 ={ core_csr_decoded_decoded_lo_hi_117 , core_csr_decoded_decoded_lo_lo_116 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_3_117 , core_csr_decoded_decoded_andMatrixInput_4_117 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_116 ={ core_csr_decoded_decoded_hi_lo_hi_115 , core_csr_decoded_decoded_andMatrixInput_5_117 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_0_117 , core_csr_decoded_decoded_andMatrixInput_1_117 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_117 ={ core_csr_decoded_decoded_hi_hi_hi_116 , core_csr_decoded_decoded_andMatrixInput_2_117 }; 
    wire[5:0] core_csr_decoded_decoded_hi_117 ={ core_csr_decoded_decoded_hi_hi_117 , core_csr_decoded_decoded_hi_lo_116 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_118 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_118 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_118 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_118 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_118 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_118 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_117 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_117 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_117 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_117 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_116 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_109 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_109 ={ core_csr_decoded_decoded_andMatrixInput_9_117 , core_csr_decoded_decoded_andMatrixInput_10_116 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_117 ={ core_csr_decoded_decoded_lo_lo_hi_109 , core_csr_decoded_decoded_andMatrixInput_11_109 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_6_117 , core_csr_decoded_decoded_andMatrixInput_7_117 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_118 ={ core_csr_decoded_decoded_lo_hi_hi_117 , core_csr_decoded_decoded_andMatrixInput_8_117 }; 
    wire[5:0] core_csr_decoded_decoded_lo_118 ={ core_csr_decoded_decoded_lo_hi_118 , core_csr_decoded_decoded_lo_lo_117 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_3_118 , core_csr_decoded_decoded_andMatrixInput_4_118 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_117 ={ core_csr_decoded_decoded_hi_lo_hi_116 , core_csr_decoded_decoded_andMatrixInput_5_118 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_0_118 , core_csr_decoded_decoded_andMatrixInput_1_118 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_118 ={ core_csr_decoded_decoded_hi_hi_hi_117 , core_csr_decoded_decoded_andMatrixInput_2_118 }; 
    wire[5:0] core_csr_decoded_decoded_hi_118 ={ core_csr_decoded_decoded_hi_hi_118 , core_csr_decoded_decoded_hi_lo_117 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_119 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_119 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_119 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_119 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_119 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_119 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_118 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_118 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_118 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_118 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_117 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_110 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_110 ={ core_csr_decoded_decoded_andMatrixInput_9_118 , core_csr_decoded_decoded_andMatrixInput_10_117 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_118 ={ core_csr_decoded_decoded_lo_lo_hi_110 , core_csr_decoded_decoded_andMatrixInput_11_110 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_6_118 , core_csr_decoded_decoded_andMatrixInput_7_118 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_119 ={ core_csr_decoded_decoded_lo_hi_hi_118 , core_csr_decoded_decoded_andMatrixInput_8_118 }; 
    wire[5:0] core_csr_decoded_decoded_lo_119 ={ core_csr_decoded_decoded_lo_hi_119 , core_csr_decoded_decoded_lo_lo_118 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_3_119 , core_csr_decoded_decoded_andMatrixInput_4_119 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_118 ={ core_csr_decoded_decoded_hi_lo_hi_117 , core_csr_decoded_decoded_andMatrixInput_5_119 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_0_119 , core_csr_decoded_decoded_andMatrixInput_1_119 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_119 ={ core_csr_decoded_decoded_hi_hi_hi_118 , core_csr_decoded_decoded_andMatrixInput_2_119 }; 
    wire[5:0] core_csr_decoded_decoded_hi_119 ={ core_csr_decoded_decoded_hi_hi_119 , core_csr_decoded_decoded_hi_lo_118 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_120 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_120 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_120 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_120 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_120 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_120 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_119 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_119 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_119 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_119 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_118 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_111 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_111 ={ core_csr_decoded_decoded_andMatrixInput_9_119 , core_csr_decoded_decoded_andMatrixInput_10_118 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_119 ={ core_csr_decoded_decoded_lo_lo_hi_111 , core_csr_decoded_decoded_andMatrixInput_11_111 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_6_119 , core_csr_decoded_decoded_andMatrixInput_7_119 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_120 ={ core_csr_decoded_decoded_lo_hi_hi_119 , core_csr_decoded_decoded_andMatrixInput_8_119 }; 
    wire[5:0] core_csr_decoded_decoded_lo_120 ={ core_csr_decoded_decoded_lo_hi_120 , core_csr_decoded_decoded_lo_lo_119 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_3_120 , core_csr_decoded_decoded_andMatrixInput_4_120 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_119 ={ core_csr_decoded_decoded_hi_lo_hi_118 , core_csr_decoded_decoded_andMatrixInput_5_120 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_0_120 , core_csr_decoded_decoded_andMatrixInput_1_120 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_120 ={ core_csr_decoded_decoded_hi_hi_hi_119 , core_csr_decoded_decoded_andMatrixInput_2_120 }; 
    wire[5:0] core_csr_decoded_decoded_hi_120 ={ core_csr_decoded_decoded_hi_hi_120 , core_csr_decoded_decoded_hi_lo_119 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_121 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_121 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_121 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_121 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_121 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_121 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_120 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_120 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_120 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_120 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_119 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_112 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_112 ={ core_csr_decoded_decoded_andMatrixInput_9_120 , core_csr_decoded_decoded_andMatrixInput_10_119 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_120 ={ core_csr_decoded_decoded_lo_lo_hi_112 , core_csr_decoded_decoded_andMatrixInput_11_112 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_6_120 , core_csr_decoded_decoded_andMatrixInput_7_120 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_121 ={ core_csr_decoded_decoded_lo_hi_hi_120 , core_csr_decoded_decoded_andMatrixInput_8_120 }; 
    wire[5:0] core_csr_decoded_decoded_lo_121 ={ core_csr_decoded_decoded_lo_hi_121 , core_csr_decoded_decoded_lo_lo_120 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_3_121 , core_csr_decoded_decoded_andMatrixInput_4_121 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_120 ={ core_csr_decoded_decoded_hi_lo_hi_119 , core_csr_decoded_decoded_andMatrixInput_5_121 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_0_121 , core_csr_decoded_decoded_andMatrixInput_1_121 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_121 ={ core_csr_decoded_decoded_hi_hi_hi_120 , core_csr_decoded_decoded_andMatrixInput_2_121 }; 
    wire[5:0] core_csr_decoded_decoded_hi_121 ={ core_csr_decoded_decoded_hi_hi_121 , core_csr_decoded_decoded_hi_lo_120 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_122 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_122 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_122 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_122 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_122 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_122 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_121 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_121 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_121 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_121 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_120 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_113 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_113 ={ core_csr_decoded_decoded_andMatrixInput_9_121 , core_csr_decoded_decoded_andMatrixInput_10_120 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_121 ={ core_csr_decoded_decoded_lo_lo_hi_113 , core_csr_decoded_decoded_andMatrixInput_11_113 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_6_121 , core_csr_decoded_decoded_andMatrixInput_7_121 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_122 ={ core_csr_decoded_decoded_lo_hi_hi_121 , core_csr_decoded_decoded_andMatrixInput_8_121 }; 
    wire[5:0] core_csr_decoded_decoded_lo_122 ={ core_csr_decoded_decoded_lo_hi_122 , core_csr_decoded_decoded_lo_lo_121 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_3_122 , core_csr_decoded_decoded_andMatrixInput_4_122 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_121 ={ core_csr_decoded_decoded_hi_lo_hi_120 , core_csr_decoded_decoded_andMatrixInput_5_122 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_0_122 , core_csr_decoded_decoded_andMatrixInput_1_122 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_122 ={ core_csr_decoded_decoded_hi_hi_hi_121 , core_csr_decoded_decoded_andMatrixInput_2_122 }; 
    wire[5:0] core_csr_decoded_decoded_hi_122 ={ core_csr_decoded_decoded_hi_hi_122 , core_csr_decoded_decoded_hi_lo_121 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_123 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_123 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_123 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_123 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_123 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_123 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_122 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_122 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_122 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_122 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_121 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_114 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_114 ={ core_csr_decoded_decoded_andMatrixInput_9_122 , core_csr_decoded_decoded_andMatrixInput_10_121 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_122 ={ core_csr_decoded_decoded_lo_lo_hi_114 , core_csr_decoded_decoded_andMatrixInput_11_114 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_6_122 , core_csr_decoded_decoded_andMatrixInput_7_122 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_123 ={ core_csr_decoded_decoded_lo_hi_hi_122 , core_csr_decoded_decoded_andMatrixInput_8_122 }; 
    wire[5:0] core_csr_decoded_decoded_lo_123 ={ core_csr_decoded_decoded_lo_hi_123 , core_csr_decoded_decoded_lo_lo_122 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_3_123 , core_csr_decoded_decoded_andMatrixInput_4_123 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_122 ={ core_csr_decoded_decoded_hi_lo_hi_121 , core_csr_decoded_decoded_andMatrixInput_5_123 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_0_123 , core_csr_decoded_decoded_andMatrixInput_1_123 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_123 ={ core_csr_decoded_decoded_hi_hi_hi_122 , core_csr_decoded_decoded_andMatrixInput_2_123 }; 
    wire[5:0] core_csr_decoded_decoded_hi_123 ={ core_csr_decoded_decoded_hi_hi_123 , core_csr_decoded_decoded_hi_lo_122 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_124 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_124 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_124 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_124 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_124 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_124 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_123 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_123 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_123 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_123 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_122 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_115 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_115 ={ core_csr_decoded_decoded_andMatrixInput_9_123 , core_csr_decoded_decoded_andMatrixInput_10_122 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_123 ={ core_csr_decoded_decoded_lo_lo_hi_115 , core_csr_decoded_decoded_andMatrixInput_11_115 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_6_123 , core_csr_decoded_decoded_andMatrixInput_7_123 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_124 ={ core_csr_decoded_decoded_lo_hi_hi_123 , core_csr_decoded_decoded_andMatrixInput_8_123 }; 
    wire[5:0] core_csr_decoded_decoded_lo_124 ={ core_csr_decoded_decoded_lo_hi_124 , core_csr_decoded_decoded_lo_lo_123 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_122 ={ core_csr_decoded_decoded_andMatrixInput_3_124 , core_csr_decoded_decoded_andMatrixInput_4_124 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_123 ={ core_csr_decoded_decoded_hi_lo_hi_122 , core_csr_decoded_decoded_andMatrixInput_5_124 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_0_124 , core_csr_decoded_decoded_andMatrixInput_1_124 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_124 ={ core_csr_decoded_decoded_hi_hi_hi_123 , core_csr_decoded_decoded_andMatrixInput_2_124 }; 
    wire[5:0] core_csr_decoded_decoded_hi_124 ={ core_csr_decoded_decoded_hi_hi_124 , core_csr_decoded_decoded_hi_lo_123 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_125 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_125 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_125 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_125 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_125 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_125 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_124 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_124 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_124 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_124 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_123 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_116 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_116 ={ core_csr_decoded_decoded_andMatrixInput_9_124 , core_csr_decoded_decoded_andMatrixInput_10_123 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_124 ={ core_csr_decoded_decoded_lo_lo_hi_116 , core_csr_decoded_decoded_andMatrixInput_11_116 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_6_124 , core_csr_decoded_decoded_andMatrixInput_7_124 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_125 ={ core_csr_decoded_decoded_lo_hi_hi_124 , core_csr_decoded_decoded_andMatrixInput_8_124 }; 
    wire[5:0] core_csr_decoded_decoded_lo_125 ={ core_csr_decoded_decoded_lo_hi_125 , core_csr_decoded_decoded_lo_lo_124 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_123 ={ core_csr_decoded_decoded_andMatrixInput_3_125 , core_csr_decoded_decoded_andMatrixInput_4_125 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_124 ={ core_csr_decoded_decoded_hi_lo_hi_123 , core_csr_decoded_decoded_andMatrixInput_5_125 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_0_125 , core_csr_decoded_decoded_andMatrixInput_1_125 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_125 ={ core_csr_decoded_decoded_hi_hi_hi_124 , core_csr_decoded_decoded_andMatrixInput_2_125 }; 
    wire[5:0] core_csr_decoded_decoded_hi_125 ={ core_csr_decoded_decoded_hi_hi_125 , core_csr_decoded_decoded_hi_lo_124 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_126 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_126 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_126 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_126 = core_csr_decoded_decoded_plaInput [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_126 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_126 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_125 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_125 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_125 = core_csr_decoded_decoded_invInputs [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_125 = core_csr_decoded_decoded_invInputs [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_124 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_117 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_117 ={ core_csr_decoded_decoded_andMatrixInput_9_125 , core_csr_decoded_decoded_andMatrixInput_10_124 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_125 ={ core_csr_decoded_decoded_lo_lo_hi_117 , core_csr_decoded_decoded_andMatrixInput_11_117 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_6_125 , core_csr_decoded_decoded_andMatrixInput_7_125 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_126 ={ core_csr_decoded_decoded_lo_hi_hi_125 , core_csr_decoded_decoded_andMatrixInput_8_125 }; 
    wire[5:0] core_csr_decoded_decoded_lo_126 ={ core_csr_decoded_decoded_lo_hi_126 , core_csr_decoded_decoded_lo_lo_125 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_124 ={ core_csr_decoded_decoded_andMatrixInput_3_126 , core_csr_decoded_decoded_andMatrixInput_4_126 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_125 ={ core_csr_decoded_decoded_hi_lo_hi_124 , core_csr_decoded_decoded_andMatrixInput_5_126 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_0_126 , core_csr_decoded_decoded_andMatrixInput_1_126 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_126 ={ core_csr_decoded_decoded_hi_hi_hi_125 , core_csr_decoded_decoded_andMatrixInput_2_126 }; 
    wire[5:0] core_csr_decoded_decoded_hi_126 ={ core_csr_decoded_decoded_hi_hi_126 , core_csr_decoded_decoded_hi_lo_125 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_127 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_127 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_127 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_127 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_127 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_127 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_126 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_126 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_126 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_126 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_125 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_126 ={ core_csr_decoded_decoded_andMatrixInput_9_126 , core_csr_decoded_decoded_andMatrixInput_10_125 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_6_126 , core_csr_decoded_decoded_andMatrixInput_7_126 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_127 ={ core_csr_decoded_decoded_lo_hi_hi_126 , core_csr_decoded_decoded_andMatrixInput_8_126 }; 
    wire[4:0] core_csr_decoded_decoded_lo_127 ={ core_csr_decoded_decoded_lo_hi_127 , core_csr_decoded_decoded_lo_lo_126 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_125 ={ core_csr_decoded_decoded_andMatrixInput_3_127 , core_csr_decoded_decoded_andMatrixInput_4_127 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_126 ={ core_csr_decoded_decoded_hi_lo_hi_125 , core_csr_decoded_decoded_andMatrixInput_5_127 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_0_127 , core_csr_decoded_decoded_andMatrixInput_1_127 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_127 ={ core_csr_decoded_decoded_hi_hi_hi_126 , core_csr_decoded_decoded_andMatrixInput_2_127 }; 
    wire[5:0] core_csr_decoded_decoded_hi_127 ={ core_csr_decoded_decoded_hi_hi_127 , core_csr_decoded_decoded_hi_lo_126 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_128 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_128 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_128 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_128 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_128 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_128 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_127 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_127 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_127 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_127 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_126 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_118 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_118 ={ core_csr_decoded_decoded_andMatrixInput_9_127 , core_csr_decoded_decoded_andMatrixInput_10_126 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_127 ={ core_csr_decoded_decoded_lo_lo_hi_118 , core_csr_decoded_decoded_andMatrixInput_11_118 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_6_127 , core_csr_decoded_decoded_andMatrixInput_7_127 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_128 ={ core_csr_decoded_decoded_lo_hi_hi_127 , core_csr_decoded_decoded_andMatrixInput_8_127 }; 
    wire[5:0] core_csr_decoded_decoded_lo_128 ={ core_csr_decoded_decoded_lo_hi_128 , core_csr_decoded_decoded_lo_lo_127 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_126 ={ core_csr_decoded_decoded_andMatrixInput_3_128 , core_csr_decoded_decoded_andMatrixInput_4_128 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_127 ={ core_csr_decoded_decoded_hi_lo_hi_126 , core_csr_decoded_decoded_andMatrixInput_5_128 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_0_128 , core_csr_decoded_decoded_andMatrixInput_1_128 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_128 ={ core_csr_decoded_decoded_hi_hi_hi_127 , core_csr_decoded_decoded_andMatrixInput_2_128 }; 
    wire[5:0] core_csr_decoded_decoded_hi_128 ={ core_csr_decoded_decoded_hi_hi_128 , core_csr_decoded_decoded_hi_lo_127 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_129 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_129 = core_csr_decoded_decoded_plaInput [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_129 = core_csr_decoded_decoded_invInputs [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_129 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_129 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_129 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_128 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_128 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_128 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_128 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_127 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_119 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_119 ={ core_csr_decoded_decoded_andMatrixInput_9_128 , core_csr_decoded_decoded_andMatrixInput_10_127 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_128 ={ core_csr_decoded_decoded_lo_lo_hi_119 , core_csr_decoded_decoded_andMatrixInput_11_119 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_6_128 , core_csr_decoded_decoded_andMatrixInput_7_128 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_129 ={ core_csr_decoded_decoded_lo_hi_hi_128 , core_csr_decoded_decoded_andMatrixInput_8_128 }; 
    wire[5:0] core_csr_decoded_decoded_lo_129 ={ core_csr_decoded_decoded_lo_hi_129 , core_csr_decoded_decoded_lo_lo_128 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_127 ={ core_csr_decoded_decoded_andMatrixInput_3_129 , core_csr_decoded_decoded_andMatrixInput_4_129 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_128 ={ core_csr_decoded_decoded_hi_lo_hi_127 , core_csr_decoded_decoded_andMatrixInput_5_129 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_0_129 , core_csr_decoded_decoded_andMatrixInput_1_129 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_129 ={ core_csr_decoded_decoded_hi_hi_hi_128 , core_csr_decoded_decoded_andMatrixInput_2_129 }; 
    wire[5:0] core_csr_decoded_decoded_hi_129 ={ core_csr_decoded_decoded_hi_hi_129 , core_csr_decoded_decoded_hi_lo_128 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_130 = core_csr_decoded_decoded_invInputs [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_130 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_130 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_130 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_130 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_130 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_129 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_129 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_129 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_129 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_128 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_120 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_120 ={ core_csr_decoded_decoded_andMatrixInput_9_129 , core_csr_decoded_decoded_andMatrixInput_10_128 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_129 ={ core_csr_decoded_decoded_lo_lo_hi_120 , core_csr_decoded_decoded_andMatrixInput_11_120 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_6_129 , core_csr_decoded_decoded_andMatrixInput_7_129 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_130 ={ core_csr_decoded_decoded_lo_hi_hi_129 , core_csr_decoded_decoded_andMatrixInput_8_129 }; 
    wire[5:0] core_csr_decoded_decoded_lo_130 ={ core_csr_decoded_decoded_lo_hi_130 , core_csr_decoded_decoded_lo_lo_129 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_128 ={ core_csr_decoded_decoded_andMatrixInput_3_130 , core_csr_decoded_decoded_andMatrixInput_4_130 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_129 ={ core_csr_decoded_decoded_hi_lo_hi_128 , core_csr_decoded_decoded_andMatrixInput_5_130 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_0_130 , core_csr_decoded_decoded_andMatrixInput_1_130 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_130 ={ core_csr_decoded_decoded_hi_hi_hi_129 , core_csr_decoded_decoded_andMatrixInput_2_130 }; 
    wire[5:0] core_csr_decoded_decoded_hi_130 ={ core_csr_decoded_decoded_hi_hi_130 , core_csr_decoded_decoded_hi_lo_129 }; 
    wire core_csr_decoded_decoded_andMatrixInput_0_131 = core_csr_decoded_decoded_plaInput [0]; 
    wire core_csr_decoded_decoded_andMatrixInput_1_131 = core_csr_decoded_decoded_invInputs [1]; 
    wire core_csr_decoded_decoded_andMatrixInput_2_131 = core_csr_decoded_decoded_plaInput [2]; 
    wire core_csr_decoded_decoded_andMatrixInput_3_131 = core_csr_decoded_decoded_invInputs [3]; 
    wire core_csr_decoded_decoded_andMatrixInput_4_131 = core_csr_decoded_decoded_plaInput [4]; 
    wire core_csr_decoded_decoded_andMatrixInput_5_131 = core_csr_decoded_decoded_invInputs [5]; 
    wire core_csr_decoded_decoded_andMatrixInput_6_130 = core_csr_decoded_decoded_invInputs [6]; 
    wire core_csr_decoded_decoded_andMatrixInput_7_130 = core_csr_decoded_decoded_invInputs [7]; 
    wire core_csr_decoded_decoded_andMatrixInput_8_130 = core_csr_decoded_decoded_plaInput [8]; 
    wire core_csr_decoded_decoded_andMatrixInput_9_130 = core_csr_decoded_decoded_plaInput [9]; 
    wire core_csr_decoded_decoded_andMatrixInput_10_129 = core_csr_decoded_decoded_plaInput [10]; 
    wire core_csr_decoded_decoded_andMatrixInput_11_121 = core_csr_decoded_decoded_plaInput [11]; 
    wire[1:0] core_csr_decoded_decoded_lo_lo_hi_121 ={ core_csr_decoded_decoded_andMatrixInput_9_130 , core_csr_decoded_decoded_andMatrixInput_10_129 }; 
    wire[2:0] core_csr_decoded_decoded_lo_lo_130 ={ core_csr_decoded_decoded_lo_lo_hi_121 , core_csr_decoded_decoded_andMatrixInput_11_121 }; 
    wire[1:0] core_csr_decoded_decoded_lo_hi_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_6_130 , core_csr_decoded_decoded_andMatrixInput_7_130 }; 
    wire[2:0] core_csr_decoded_decoded_lo_hi_131 ={ core_csr_decoded_decoded_lo_hi_hi_130 , core_csr_decoded_decoded_andMatrixInput_8_130 }; 
    wire[5:0] core_csr_decoded_decoded_lo_131 ={ core_csr_decoded_decoded_lo_hi_131 , core_csr_decoded_decoded_lo_lo_130 }; 
    wire[1:0] core_csr_decoded_decoded_hi_lo_hi_129 ={ core_csr_decoded_decoded_andMatrixInput_3_131 , core_csr_decoded_decoded_andMatrixInput_4_131 }; 
    wire[2:0] core_csr_decoded_decoded_hi_lo_130 ={ core_csr_decoded_decoded_hi_lo_hi_129 , core_csr_decoded_decoded_andMatrixInput_5_131 }; 
    wire[1:0] core_csr_decoded_decoded_hi_hi_hi_130 ={ core_csr_decoded_decoded_andMatrixInput_0_131 , core_csr_decoded_decoded_andMatrixInput_1_131 }; 
    wire[2:0] core_csr_decoded_decoded_hi_hi_131 ={ core_csr_decoded_decoded_hi_hi_hi_130 , core_csr_decoded_decoded_andMatrixInput_2_131 }; 
    wire[5:0] core_csr_decoded_decoded_hi_131 ={ core_csr_decoded_decoded_hi_hi_131 , core_csr_decoded_decoded_hi_lo_130 }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_129 , core_csr_decoded_decoded_lo_129 }),|(&{ core_csr_decoded_decoded_hi_131 , core_csr_decoded_decoded_lo_131 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_128 , core_csr_decoded_decoded_lo_128 }),|(&{ core_csr_decoded_decoded_hi_127 , core_csr_decoded_decoded_lo_127 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_56 , core_csr_decoded_decoded_lo_56 }),|(&{ core_csr_decoded_decoded_hi_64 , core_csr_decoded_decoded_lo_64 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_54 , core_csr_decoded_decoded_lo_54 }),|(&{ core_csr_decoded_decoded_hi_55 , core_csr_decoded_decoded_lo_55 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_52 , core_csr_decoded_decoded_lo_52 }),|(&{ core_csr_decoded_decoded_hi_53 , core_csr_decoded_decoded_lo_53 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_50 , core_csr_decoded_decoded_lo_50 }),|(&{ core_csr_decoded_decoded_hi_51 , core_csr_decoded_decoded_lo_51 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_48 , core_csr_decoded_decoded_lo_48 }),|(&{ core_csr_decoded_decoded_hi_49 , core_csr_decoded_decoded_lo_49 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_46 , core_csr_decoded_decoded_lo_46 }),|(&{ core_csr_decoded_decoded_hi_47 , core_csr_decoded_decoded_lo_47 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_44 , core_csr_decoded_decoded_lo_44 }),|(&{ core_csr_decoded_decoded_hi_45 , core_csr_decoded_decoded_lo_45 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_42 , core_csr_decoded_decoded_lo_42 }),|(&{ core_csr_decoded_decoded_hi_43 , core_csr_decoded_decoded_lo_43 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_40 , core_csr_decoded_decoded_lo_40 }),|(&{ core_csr_decoded_decoded_hi_41 , core_csr_decoded_decoded_lo_41 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_97 , core_csr_decoded_decoded_lo_97 }),|(&{ core_csr_decoded_decoded_hi_39 , core_csr_decoded_decoded_lo_39 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_126 , core_csr_decoded_decoded_lo_126 }),|(&{ core_csr_decoded_decoded_hi_96 , core_csr_decoded_decoded_lo_96 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_33 , core_csr_decoded_decoded_lo_33 }),|(&{ core_csr_decoded_decoded_hi_95 , core_csr_decoded_decoded_lo_95 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_94 , core_csr_decoded_decoded_lo_94 }),|(&{ core_csr_decoded_decoded_hi_125 , core_csr_decoded_decoded_lo_125 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_93 , core_csr_decoded_decoded_lo_93 }),|(&{ core_csr_decoded_decoded_hi_124 , core_csr_decoded_decoded_lo_124 })}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi_hi ,|(&{ core_csr_decoded_decoded_hi_32 , core_csr_decoded_decoded_lo_32 })}; 
    wire[4:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_orMatrixOutputs_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_123 , core_csr_decoded_decoded_lo_123 }),|(&{ core_csr_decoded_decoded_hi_31 , core_csr_decoded_decoded_lo_31 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_30 , core_csr_decoded_decoded_lo_30 }),|(&{ core_csr_decoded_decoded_hi_92 , core_csr_decoded_decoded_lo_92 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_91 , core_csr_decoded_decoded_lo_91 }),|(&{ core_csr_decoded_decoded_hi_122 , core_csr_decoded_decoded_lo_122 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_121 , core_csr_decoded_decoded_lo_121 }),|(&{ core_csr_decoded_decoded_hi_29 , core_csr_decoded_decoded_lo_29 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_28 , core_csr_decoded_decoded_lo_28 }),|(&{ core_csr_decoded_decoded_hi_90 , core_csr_decoded_decoded_lo_90 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_89 , core_csr_decoded_decoded_lo_89 }),|(&{ core_csr_decoded_decoded_hi_120 , core_csr_decoded_decoded_lo_120 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_119 , core_csr_decoded_decoded_lo_119 }),|(&{ core_csr_decoded_decoded_hi_27 , core_csr_decoded_decoded_lo_27 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_26 , core_csr_decoded_decoded_lo_26 }),|(&{ core_csr_decoded_decoded_hi_88 , core_csr_decoded_decoded_lo_88 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_87 , core_csr_decoded_decoded_lo_87 }),|(&{ core_csr_decoded_decoded_hi_118 , core_csr_decoded_decoded_lo_118 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_117 , core_csr_decoded_decoded_lo_117 }),|(&{ core_csr_decoded_decoded_hi_25 , core_csr_decoded_decoded_lo_25 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_24 , core_csr_decoded_decoded_lo_24 }),|(&{ core_csr_decoded_decoded_hi_86 , core_csr_decoded_decoded_lo_86 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_85 , core_csr_decoded_decoded_lo_85 }),|(&{ core_csr_decoded_decoded_hi_116 , core_csr_decoded_decoded_lo_116 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_115 , core_csr_decoded_decoded_lo_115 }),|(&{ core_csr_decoded_decoded_hi_23 , core_csr_decoded_decoded_lo_23 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_22 , core_csr_decoded_decoded_lo_22 }),|(&{ core_csr_decoded_decoded_hi_84 , core_csr_decoded_decoded_lo_84 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_83 , core_csr_decoded_decoded_lo_83 }),|(&{ core_csr_decoded_decoded_hi_114 , core_csr_decoded_decoded_lo_114 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_82 , core_csr_decoded_decoded_lo_82 }),|(&{ core_csr_decoded_decoded_hi_113 , core_csr_decoded_decoded_lo_113 })}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi_hi ,|(&{ core_csr_decoded_decoded_hi_21 , core_csr_decoded_decoded_lo_21 })}; 
    wire[4:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_orMatrixOutputs_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_hi_lo }; 
    wire[65:0] core_csr_decoded_decoded_orMatrixOutputs_lo ={ core_csr_decoded_decoded_orMatrixOutputs_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_112 , core_csr_decoded_decoded_lo_112 }),|(&{ core_csr_decoded_decoded_hi_20 , core_csr_decoded_decoded_lo_20 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_19 , core_csr_decoded_decoded_lo_19 }),|(&{ core_csr_decoded_decoded_hi_81 , core_csr_decoded_decoded_lo_81 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_80 , core_csr_decoded_decoded_lo_80 }),|(&{ core_csr_decoded_decoded_hi_111 , core_csr_decoded_decoded_lo_111 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_110 , core_csr_decoded_decoded_lo_110 }),|(&{ core_csr_decoded_decoded_hi_18 , core_csr_decoded_decoded_lo_18 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_17 , core_csr_decoded_decoded_lo_17 }),|(&{ core_csr_decoded_decoded_hi_79 , core_csr_decoded_decoded_lo_79 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_78 , core_csr_decoded_decoded_lo_78 }),|(&{ core_csr_decoded_decoded_hi_109 , core_csr_decoded_decoded_lo_109 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_108 , core_csr_decoded_decoded_lo_108 }),|(&{ core_csr_decoded_decoded_hi_16 , core_csr_decoded_decoded_lo_16 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_15 , core_csr_decoded_decoded_lo_15 }),|(&{ core_csr_decoded_decoded_hi_77 , core_csr_decoded_decoded_lo_77 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_76 , core_csr_decoded_decoded_lo_76 }),|(&{ core_csr_decoded_decoded_hi_107 , core_csr_decoded_decoded_lo_107 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_106 , core_csr_decoded_decoded_lo_106 }),|(&{ core_csr_decoded_decoded_hi_14 , core_csr_decoded_decoded_lo_14 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_13 , core_csr_decoded_decoded_lo_13 }),|(&{ core_csr_decoded_decoded_hi_75 , core_csr_decoded_decoded_lo_75 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_74 , core_csr_decoded_decoded_lo_74 }),|(&{ core_csr_decoded_decoded_hi_105 , core_csr_decoded_decoded_lo_105 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_104 , core_csr_decoded_decoded_lo_104 }),|(&{ core_csr_decoded_decoded_hi_12 , core_csr_decoded_decoded_lo_12 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_11 , core_csr_decoded_decoded_lo_11 }),|(&{ core_csr_decoded_decoded_hi_73 , core_csr_decoded_decoded_lo_73 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_72 , core_csr_decoded_decoded_lo_72 }),|(&{ core_csr_decoded_decoded_hi_103 , core_csr_decoded_decoded_lo_103 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_71 , core_csr_decoded_decoded_lo_71 }),|(&{ core_csr_decoded_decoded_hi_102 , core_csr_decoded_decoded_lo_102 })}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi_hi ,|(&{ core_csr_decoded_decoded_hi_10 , core_csr_decoded_decoded_lo_10 })}; 
    wire[4:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_orMatrixOutputs_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_101 , core_csr_decoded_decoded_lo_101 }),|(&{ core_csr_decoded_decoded_hi_9 , core_csr_decoded_decoded_lo_9 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_8 , core_csr_decoded_decoded_lo_8 }),|(&{ core_csr_decoded_decoded_hi_70 , core_csr_decoded_decoded_lo_70 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_69 , core_csr_decoded_decoded_lo_69 }),|(&{ core_csr_decoded_decoded_hi_100 , core_csr_decoded_decoded_lo_100 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_99 , core_csr_decoded_decoded_lo_99 }),|(&{ core_csr_decoded_decoded_hi_7 , core_csr_decoded_decoded_lo_7 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_6 , core_csr_decoded_decoded_lo_6 }),|(&{ core_csr_decoded_decoded_hi_68 , core_csr_decoded_decoded_lo_68 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi_67 , core_csr_decoded_decoded_lo_67 }),|(&{ core_csr_decoded_decoded_hi_98 , core_csr_decoded_decoded_lo_98 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_66 , core_csr_decoded_decoded_lo_66 }),|(&{ core_csr_decoded_decoded_hi_5 , core_csr_decoded_decoded_lo_5 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_4 , core_csr_decoded_decoded_lo_4 }),|(&{ core_csr_decoded_decoded_hi_65 , core_csr_decoded_decoded_lo_65 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo ={|(&{ core_csr_decoded_decoded_hi_62 , core_csr_decoded_decoded_lo_62 }),|(&{ core_csr_decoded_decoded_hi_63 , core_csr_decoded_decoded_lo_63 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi ={|(&{ core_csr_decoded_decoded_hi_130 , core_csr_decoded_decoded_lo_130 }),|(&{ core_csr_decoded_decoded_hi_61 , core_csr_decoded_decoded_lo_61 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo ={|(&{ core_csr_decoded_decoded_hi_37 , core_csr_decoded_decoded_lo_37 }),|(&{ core_csr_decoded_decoded_hi_36 , core_csr_decoded_decoded_lo_36 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi ={|(&{ core_csr_decoded_decoded_hi_34 , core_csr_decoded_decoded_lo_34 }),|(&{ core_csr_decoded_decoded_hi_35 , core_csr_decoded_decoded_lo_35 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo ={|(&{ core_csr_decoded_decoded_hi_38 , core_csr_decoded_decoded_lo_38 }),|(&{ core_csr_decoded_decoded_hi_2 , core_csr_decoded_decoded_lo_2 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi ={|(&{ core_csr_decoded_decoded_hi , core_csr_decoded_decoded_lo }),|(&{ core_csr_decoded_decoded_hi_3 , core_csr_decoded_decoded_lo_3 })}; 
    wire[3:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo ={|(&{ core_csr_decoded_decoded_hi_60 , core_csr_decoded_decoded_lo_60 }),|(&{ core_csr_decoded_decoded_hi_1 , core_csr_decoded_decoded_lo_1 })}; 
    wire[1:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_hi ={|(&{ core_csr_decoded_decoded_hi_57 , core_csr_decoded_decoded_lo_57 }),|(&{ core_csr_decoded_decoded_hi_58 , core_csr_decoded_decoded_lo_58 })}; 
    wire[2:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi_hi ,|(&{ core_csr_decoded_decoded_hi_59 , core_csr_decoded_decoded_lo_59 })}; 
    wire[4:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_orMatrixOutputs_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_hi_lo }; 
    wire[65:0] core_csr_decoded_decoded_orMatrixOutputs_hi ={ core_csr_decoded_decoded_orMatrixOutputs_hi_hi , core_csr_decoded_decoded_orMatrixOutputs_hi_lo }; 
    wire[131:0] core_csr_decoded_decoded_orMatrixOutputs ={ core_csr_decoded_decoded_orMatrixOutputs_hi , core_csr_decoded_decoded_orMatrixOutputs_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [1], core_csr_decoded_decoded_orMatrixOutputs [0]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [3], core_csr_decoded_decoded_orMatrixOutputs [2]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [5], core_csr_decoded_decoded_orMatrixOutputs [4]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [7], core_csr_decoded_decoded_orMatrixOutputs [6]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [9], core_csr_decoded_decoded_orMatrixOutputs [8]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [11], core_csr_decoded_decoded_orMatrixOutputs [10]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [13], core_csr_decoded_decoded_orMatrixOutputs [12]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [15], core_csr_decoded_decoded_orMatrixOutputs [14]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [17], core_csr_decoded_decoded_orMatrixOutputs [16]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [19], core_csr_decoded_decoded_orMatrixOutputs [18]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [21], core_csr_decoded_decoded_orMatrixOutputs [20]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [23], core_csr_decoded_decoded_orMatrixOutputs [22]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [25], core_csr_decoded_decoded_orMatrixOutputs [24]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [27], core_csr_decoded_decoded_orMatrixOutputs [26]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [29], core_csr_decoded_decoded_orMatrixOutputs [28]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [32], core_csr_decoded_decoded_orMatrixOutputs [31]}; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [30]}; 
    wire[4:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_invMatrixOutputs_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [34], core_csr_decoded_decoded_orMatrixOutputs [33]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [36], core_csr_decoded_decoded_orMatrixOutputs [35]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [38], core_csr_decoded_decoded_orMatrixOutputs [37]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [40], core_csr_decoded_decoded_orMatrixOutputs [39]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [42], core_csr_decoded_decoded_orMatrixOutputs [41]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [44], core_csr_decoded_decoded_orMatrixOutputs [43]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [46], core_csr_decoded_decoded_orMatrixOutputs [45]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [48], core_csr_decoded_decoded_orMatrixOutputs [47]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [50], core_csr_decoded_decoded_orMatrixOutputs [49]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [52], core_csr_decoded_decoded_orMatrixOutputs [51]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [54], core_csr_decoded_decoded_orMatrixOutputs [53]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [56], core_csr_decoded_decoded_orMatrixOutputs [55]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [58], core_csr_decoded_decoded_orMatrixOutputs [57]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [60], core_csr_decoded_decoded_orMatrixOutputs [59]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [62], core_csr_decoded_decoded_orMatrixOutputs [61]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [65], core_csr_decoded_decoded_orMatrixOutputs [64]}; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [63]}; 
    wire[4:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_invMatrixOutputs_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_hi_lo }; 
    wire[65:0] core_csr_decoded_decoded_invMatrixOutputs_lo ={ core_csr_decoded_decoded_invMatrixOutputs_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [67], core_csr_decoded_decoded_orMatrixOutputs [66]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [69], core_csr_decoded_decoded_orMatrixOutputs [68]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [71], core_csr_decoded_decoded_orMatrixOutputs [70]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [73], core_csr_decoded_decoded_orMatrixOutputs [72]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [75], core_csr_decoded_decoded_orMatrixOutputs [74]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [77], core_csr_decoded_decoded_orMatrixOutputs [76]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [79], core_csr_decoded_decoded_orMatrixOutputs [78]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [81], core_csr_decoded_decoded_orMatrixOutputs [80]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [83], core_csr_decoded_decoded_orMatrixOutputs [82]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [85], core_csr_decoded_decoded_orMatrixOutputs [84]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [87], core_csr_decoded_decoded_orMatrixOutputs [86]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [89], core_csr_decoded_decoded_orMatrixOutputs [88]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [91], core_csr_decoded_decoded_orMatrixOutputs [90]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [93], core_csr_decoded_decoded_orMatrixOutputs [92]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [95], core_csr_decoded_decoded_orMatrixOutputs [94]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [98], core_csr_decoded_decoded_orMatrixOutputs [97]}; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [96]}; 
    wire[4:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_invMatrixOutputs_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [100], core_csr_decoded_decoded_orMatrixOutputs [99]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [102], core_csr_decoded_decoded_orMatrixOutputs [101]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [104], core_csr_decoded_decoded_orMatrixOutputs [103]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [106], core_csr_decoded_decoded_orMatrixOutputs [105]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [108], core_csr_decoded_decoded_orMatrixOutputs [107]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [110], core_csr_decoded_decoded_orMatrixOutputs [109]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [112], core_csr_decoded_decoded_orMatrixOutputs [111]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [114], core_csr_decoded_decoded_orMatrixOutputs [113]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi_lo }; 
    wire[15:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [116], core_csr_decoded_decoded_orMatrixOutputs [115]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [118], core_csr_decoded_decoded_orMatrixOutputs [117]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [120], core_csr_decoded_decoded_orMatrixOutputs [119]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [122], core_csr_decoded_decoded_orMatrixOutputs [121]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi_lo }; 
    wire[7:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo ={ core_csr_decoded_decoded_orMatrixOutputs [124], core_csr_decoded_decoded_orMatrixOutputs [123]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi ={ core_csr_decoded_decoded_orMatrixOutputs [126], core_csr_decoded_decoded_orMatrixOutputs [125]}; 
    wire[3:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo_lo }; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo ={ core_csr_decoded_decoded_orMatrixOutputs [128], core_csr_decoded_decoded_orMatrixOutputs [127]}; 
    wire[1:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_orMatrixOutputs [131], core_csr_decoded_decoded_orMatrixOutputs [130]}; 
    wire[2:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_orMatrixOutputs [129]}; 
    wire[4:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi_lo }; 
    wire[8:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi_lo }; 
    wire[16:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi_lo }; 
    wire[32:0] core_csr_decoded_decoded_invMatrixOutputs_hi_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_hi_lo }; 
    wire[65:0] core_csr_decoded_decoded_invMatrixOutputs_hi ={ core_csr_decoded_decoded_invMatrixOutputs_hi_hi , core_csr_decoded_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_csr_decoded_decoded_invMatrixOutputs ={ core_csr_decoded_decoded_invMatrixOutputs_hi , core_csr_decoded_decoded_invMatrixOutputs_lo }; 
    wire[131:0] core_csr_decoded_decoded = core_csr_decoded_decoded_invMatrixOutputs ; 
  assign  core_csr_decoded_decoded_plaInput = core_csr_addr [11:0]; 
    wire core_csr_decoded_0 = core_csr_decoded_decoded [131]; 
    wire core_csr_decoded_1 = core_csr_decoded_decoded [130]; 
    wire core_csr_decoded_2 = core_csr_decoded_decoded [129]; 
    wire core_csr_decoded_3 = core_csr_decoded_decoded [128]; 
    wire core_csr_decoded_4 = core_csr_decoded_decoded [127]; 
    wire core_csr_decoded_5 = core_csr_decoded_decoded [126]; 
    wire core_csr_decoded_6 = core_csr_decoded_decoded [125]; 
    wire core_csr_decoded_7 = core_csr_decoded_decoded [124]; 
    wire core_csr_decoded_8 = core_csr_decoded_decoded [123]; 
    wire core_csr_decoded_9 = core_csr_decoded_decoded [122]; 
    wire core_csr_decoded_10 = core_csr_decoded_decoded [121]; 
    wire core_csr_decoded_11 = core_csr_decoded_decoded [120]; 
    wire core_csr_decoded_12 = core_csr_decoded_decoded [119]; 
    wire core_csr_decoded_13 = core_csr_decoded_decoded [118]; 
    wire core_csr_decoded_14 = core_csr_decoded_decoded [117]; 
    wire core_csr_decoded_15 = core_csr_decoded_decoded [116]; 
    wire core_csr_decoded_16 = core_csr_decoded_decoded [115]; 
    wire core_csr_decoded_17 = core_csr_decoded_decoded [114]; 
    wire core_csr_decoded_18 = core_csr_decoded_decoded [113]; 
    wire core_csr_decoded_19 = core_csr_decoded_decoded [112]; 
    wire core_csr_decoded_20 = core_csr_decoded_decoded [111]; 
    wire core_csr_decoded_21 = core_csr_decoded_decoded [110]; 
    wire core_csr_decoded_22 = core_csr_decoded_decoded [109]; 
    wire core_csr_decoded_23 = core_csr_decoded_decoded [108]; 
    wire core_csr_decoded_24 = core_csr_decoded_decoded [107]; 
    wire core_csr_decoded_25 = core_csr_decoded_decoded [106]; 
    wire core_csr_decoded_26 = core_csr_decoded_decoded [105]; 
    wire core_csr_decoded_27 = core_csr_decoded_decoded [104]; 
    wire core_csr_decoded_28 = core_csr_decoded_decoded [103]; 
    wire core_csr_decoded_29 = core_csr_decoded_decoded [102]; 
    wire core_csr_decoded_30 = core_csr_decoded_decoded [101]; 
    wire core_csr_decoded_31 = core_csr_decoded_decoded [100]; 
    wire core_csr_decoded_32 = core_csr_decoded_decoded [99]; 
    wire core_csr_decoded_33 = core_csr_decoded_decoded [98]; 
    wire core_csr_decoded_34 = core_csr_decoded_decoded [97]; 
    wire core_csr_decoded_35 = core_csr_decoded_decoded [96]; 
    wire core_csr_decoded_36 = core_csr_decoded_decoded [95]; 
    wire core_csr_decoded_37 = core_csr_decoded_decoded [94]; 
    wire core_csr_decoded_38 = core_csr_decoded_decoded [93]; 
    wire core_csr_decoded_39 = core_csr_decoded_decoded [92]; 
    wire core_csr_decoded_40 = core_csr_decoded_decoded [91]; 
    wire core_csr_decoded_41 = core_csr_decoded_decoded [90]; 
    wire core_csr_decoded_42 = core_csr_decoded_decoded [89]; 
    wire core_csr_decoded_43 = core_csr_decoded_decoded [88]; 
    wire core_csr_decoded_44 = core_csr_decoded_decoded [87]; 
    wire core_csr_decoded_45 = core_csr_decoded_decoded [86]; 
    wire core_csr_decoded_46 = core_csr_decoded_decoded [85]; 
    wire core_csr_decoded_47 = core_csr_decoded_decoded [84]; 
    wire core_csr_decoded_48 = core_csr_decoded_decoded [83]; 
    wire core_csr_decoded_49 = core_csr_decoded_decoded [82]; 
    wire core_csr_decoded_50 = core_csr_decoded_decoded [81]; 
    wire core_csr_decoded_51 = core_csr_decoded_decoded [80]; 
    wire core_csr_decoded_52 = core_csr_decoded_decoded [79]; 
    wire core_csr_decoded_53 = core_csr_decoded_decoded [78]; 
    wire core_csr_decoded_54 = core_csr_decoded_decoded [77]; 
    wire core_csr_decoded_55 = core_csr_decoded_decoded [76]; 
    wire core_csr_decoded_56 = core_csr_decoded_decoded [75]; 
    wire core_csr_decoded_57 = core_csr_decoded_decoded [74]; 
    wire core_csr_decoded_58 = core_csr_decoded_decoded [73]; 
    wire core_csr_decoded_59 = core_csr_decoded_decoded [72]; 
    wire core_csr_decoded_60 = core_csr_decoded_decoded [71]; 
    wire core_csr_decoded_61 = core_csr_decoded_decoded [70]; 
    wire core_csr_decoded_62 = core_csr_decoded_decoded [69]; 
    wire core_csr_decoded_63 = core_csr_decoded_decoded [68]; 
    wire core_csr_decoded_64 = core_csr_decoded_decoded [67]; 
    wire core_csr_decoded_65 = core_csr_decoded_decoded [66]; 
    wire core_csr_decoded_66 = core_csr_decoded_decoded [65]; 
    wire core_csr_decoded_67 = core_csr_decoded_decoded [64]; 
    wire core_csr_decoded_68 = core_csr_decoded_decoded [63]; 
    wire core_csr_decoded_69 = core_csr_decoded_decoded [62]; 
    wire core_csr_decoded_70 = core_csr_decoded_decoded [61]; 
    wire core_csr_decoded_71 = core_csr_decoded_decoded [60]; 
    wire core_csr_decoded_72 = core_csr_decoded_decoded [59]; 
    wire core_csr_decoded_73 = core_csr_decoded_decoded [58]; 
    wire core_csr_decoded_74 = core_csr_decoded_decoded [57]; 
    wire core_csr_decoded_75 = core_csr_decoded_decoded [56]; 
    wire core_csr_decoded_76 = core_csr_decoded_decoded [55]; 
    wire core_csr_decoded_77 = core_csr_decoded_decoded [54]; 
    wire core_csr_decoded_78 = core_csr_decoded_decoded [53]; 
    wire core_csr_decoded_79 = core_csr_decoded_decoded [52]; 
    wire core_csr_decoded_80 = core_csr_decoded_decoded [51]; 
    wire core_csr_decoded_81 = core_csr_decoded_decoded [50]; 
    wire core_csr_decoded_82 = core_csr_decoded_decoded [49]; 
    wire core_csr_decoded_83 = core_csr_decoded_decoded [48]; 
    wire core_csr_decoded_84 = core_csr_decoded_decoded [47]; 
    wire core_csr_decoded_85 = core_csr_decoded_decoded [46]; 
    wire core_csr_decoded_86 = core_csr_decoded_decoded [45]; 
    wire core_csr_decoded_87 = core_csr_decoded_decoded [44]; 
    wire core_csr_decoded_88 = core_csr_decoded_decoded [43]; 
    wire core_csr_decoded_89 = core_csr_decoded_decoded [42]; 
    wire core_csr_decoded_90 = core_csr_decoded_decoded [41]; 
    wire core_csr_decoded_91 = core_csr_decoded_decoded [40]; 
    wire core_csr_decoded_92 = core_csr_decoded_decoded [39]; 
    wire core_csr_decoded_93 = core_csr_decoded_decoded [38]; 
    wire core_csr_decoded_94 = core_csr_decoded_decoded [37]; 
    wire core_csr_decoded_95 = core_csr_decoded_decoded [36]; 
    wire core_csr_decoded_96 = core_csr_decoded_decoded [35]; 
    wire core_csr_decoded_97 = core_csr_decoded_decoded [34]; 
    wire core_csr_decoded_98 = core_csr_decoded_decoded [33]; 
    wire core_csr_decoded_99 = core_csr_decoded_decoded [32]; 
    wire core_csr_decoded_100 = core_csr_decoded_decoded [31]; 
    wire core_csr_decoded_101 = core_csr_decoded_decoded [30]; 
    wire core_csr_decoded_102 = core_csr_decoded_decoded [29]; 
    wire core_csr_decoded_103 = core_csr_decoded_decoded [28]; 
    wire core_csr_decoded_104 = core_csr_decoded_decoded [27]; 
    wire core_csr_decoded_105 = core_csr_decoded_decoded [26]; 
    wire core_csr_decoded_106 = core_csr_decoded_decoded [25]; 
    wire core_csr_decoded_107 = core_csr_decoded_decoded [24]; 
    wire core_csr_decoded_108 = core_csr_decoded_decoded [23]; 
    wire core_csr_decoded_109 = core_csr_decoded_decoded [22]; 
    wire core_csr_decoded_110 = core_csr_decoded_decoded [21]; 
    wire core_csr_decoded_111 = core_csr_decoded_decoded [20]; 
    wire core_csr_decoded_112 = core_csr_decoded_decoded [19]; 
    wire core_csr_decoded_113 = core_csr_decoded_decoded [18]; 
    wire core_csr_decoded_114 = core_csr_decoded_decoded [17]; 
    wire core_csr_decoded_115 = core_csr_decoded_decoded [16]; 
    wire core_csr_decoded_116 = core_csr_decoded_decoded [15]; 
    wire core_csr_decoded_117 = core_csr_decoded_decoded [14]; 
    wire core_csr_decoded_118 = core_csr_decoded_decoded [13]; 
    wire core_csr_decoded_119 = core_csr_decoded_decoded [12]; 
    wire core_csr_decoded_120 = core_csr_decoded_decoded [11]; 
    wire core_csr_decoded_121 = core_csr_decoded_decoded [10]; 
    wire core_csr_decoded_122 = core_csr_decoded_decoded [9]; 
    wire core_csr_decoded_123 = core_csr_decoded_decoded [8]; 
    wire core_csr_decoded_124 = core_csr_decoded_decoded [7]; 
    wire core_csr_decoded_125 = core_csr_decoded_decoded [6]; 
    wire core_csr_decoded_126 = core_csr_decoded_decoded [5]; 
    wire core_csr_decoded_127 = core_csr_decoded_decoded [4]; 
    wire core_csr_decoded_128 = core_csr_decoded_decoded [3]; 
    wire core_csr_decoded_129 = core_csr_decoded_decoded [2]; 
    wire core_csr_decoded_130 = core_csr_decoded_decoded [1]; 
    wire core_csr_decoded_131 = core_csr_decoded_decoded [0]; 
    wire[63:0] core_csr__io_rw_rdata_output ; 
    wire[63:0] core_csr_wdata =(( core_csr_io_rw_cmd [1] ?  core_csr__io_rw_rdata_output :64'h0)| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :64'h0); 
    wire[63:0] core_csr__reg_bp_0_control_WIRE_1 = core_csr_wdata ; 
    wire[63:0] core_csr__reg_bp_1_control_WIRE_1 = core_csr_wdata ; 
    wire core_csr_system_insn = core_csr_io_rw_cmd ==3'h4; 
    wire[31:0] core_csr_insn ={ core_csr_io_rw_addr ,20'h0}|32'h73; 
    wire[31:0] core_csr_decoded_plaInput = core_csr_insn ; 
    wire[31:0] core_csr_decoded_invInputs =~ core_csr_decoded_plaInput ; 
    wire[8:0] core_csr_decoded_invMatrixOutputs ; 
    wire core_csr_decoded_andMatrixInput_0 = core_csr_decoded_invInputs [20]; 
    wire core_csr_decoded_andMatrixInput_1 = core_csr_decoded_invInputs [21]; 
    wire core_csr_decoded_andMatrixInput_2 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_3 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_4 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_5 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_6 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_7 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_8 = core_csr_decoded_invInputs [28]; 
    wire core_csr_decoded_andMatrixInput_9 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_10 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_11 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi ={ core_csr_decoded_andMatrixInput_9 , core_csr_decoded_andMatrixInput_10 }; 
    wire[2:0] core_csr_decoded_lo_lo ={ core_csr_decoded_lo_lo_hi , core_csr_decoded_andMatrixInput_11 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi ={ core_csr_decoded_andMatrixInput_6 , core_csr_decoded_andMatrixInput_7 }; 
    wire[2:0] core_csr_decoded_lo_hi ={ core_csr_decoded_lo_hi_hi , core_csr_decoded_andMatrixInput_8 }; 
    wire[5:0] core_csr_decoded_lo ={ core_csr_decoded_lo_hi , core_csr_decoded_lo_lo }; 
    wire[1:0] core_csr_decoded_hi_lo_hi ={ core_csr_decoded_andMatrixInput_3 , core_csr_decoded_andMatrixInput_4 }; 
    wire[2:0] core_csr_decoded_hi_lo ={ core_csr_decoded_hi_lo_hi , core_csr_decoded_andMatrixInput_5 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi ={ core_csr_decoded_andMatrixInput_0 , core_csr_decoded_andMatrixInput_1 }; 
    wire[2:0] core_csr_decoded_hi_hi ={ core_csr_decoded_hi_hi_hi , core_csr_decoded_andMatrixInput_2 }; 
    wire[5:0] core_csr_decoded_hi ={ core_csr_decoded_hi_hi , core_csr_decoded_hi_lo }; 
    wire core_csr_decoded_andMatrixInput_0_1 = core_csr_decoded_plaInput [20]; 
    wire core_csr_decoded_andMatrixInput_1_1 = core_csr_decoded_invInputs [21]; 
    wire core_csr_decoded_andMatrixInput_2_1 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_3_1 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_4_1 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_5_1 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_6_1 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_7_1 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_8_1 = core_csr_decoded_invInputs [28]; 
    wire core_csr_decoded_andMatrixInput_9_1 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_10_1 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_11_1 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_1 ={ core_csr_decoded_andMatrixInput_9_1 , core_csr_decoded_andMatrixInput_10_1 }; 
    wire[2:0] core_csr_decoded_lo_lo_1 ={ core_csr_decoded_lo_lo_hi_1 , core_csr_decoded_andMatrixInput_11_1 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_1 ={ core_csr_decoded_andMatrixInput_6_1 , core_csr_decoded_andMatrixInput_7_1 }; 
    wire[2:0] core_csr_decoded_lo_hi_1 ={ core_csr_decoded_lo_hi_hi_1 , core_csr_decoded_andMatrixInput_8_1 }; 
    wire[5:0] core_csr_decoded_lo_1 ={ core_csr_decoded_lo_hi_1 , core_csr_decoded_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_1 ={ core_csr_decoded_andMatrixInput_3_1 , core_csr_decoded_andMatrixInput_4_1 }; 
    wire[2:0] core_csr_decoded_hi_lo_1 ={ core_csr_decoded_hi_lo_hi_1 , core_csr_decoded_andMatrixInput_5_1 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_1 ={ core_csr_decoded_andMatrixInput_0_1 , core_csr_decoded_andMatrixInput_1_1 }; 
    wire[2:0] core_csr_decoded_hi_hi_1 ={ core_csr_decoded_hi_hi_hi_1 , core_csr_decoded_andMatrixInput_2_1 }; 
    wire[5:0] core_csr_decoded_hi_1 ={ core_csr_decoded_hi_hi_1 , core_csr_decoded_hi_lo_1 }; 
    wire core_csr_decoded_andMatrixInput_0_2 = core_csr_decoded_plaInput [28]; 
    wire core_csr_decoded_andMatrixInput_1_2 = core_csr_decoded_invInputs [29]; 
    wire core_csr_decoded_andMatrixInput_2_2 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_3_2 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_2 ={ core_csr_decoded_andMatrixInput_2_2 , core_csr_decoded_andMatrixInput_3_2 }; 
    wire[1:0] core_csr_decoded_hi_2 ={ core_csr_decoded_andMatrixInput_0_2 , core_csr_decoded_andMatrixInput_1_2 }; 
    wire core_csr_decoded_andMatrixInput_0_3 = core_csr_decoded_invInputs [22]; 
    wire core_csr_decoded_andMatrixInput_1_3 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_2_3 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_3_3 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_4_2 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_5_2 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_6_2 = core_csr_decoded_plaInput [28]; 
    wire core_csr_decoded_andMatrixInput_7_2 = core_csr_decoded_plaInput [29]; 
    wire core_csr_decoded_andMatrixInput_8_2 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_9_2 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_lo_2 ={ core_csr_decoded_andMatrixInput_8_2 , core_csr_decoded_andMatrixInput_9_2 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_2 ={ core_csr_decoded_andMatrixInput_5_2 , core_csr_decoded_andMatrixInput_6_2 }; 
    wire[2:0] core_csr_decoded_lo_hi_2 ={ core_csr_decoded_lo_hi_hi_2 , core_csr_decoded_andMatrixInput_7_2 }; 
    wire[4:0] core_csr_decoded_lo_3 ={ core_csr_decoded_lo_hi_2 , core_csr_decoded_lo_lo_2 }; 
    wire[1:0] core_csr_decoded_hi_lo_2 ={ core_csr_decoded_andMatrixInput_3_3 , core_csr_decoded_andMatrixInput_4_2 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_2 ={ core_csr_decoded_andMatrixInput_0_3 , core_csr_decoded_andMatrixInput_1_3 }; 
    wire[2:0] core_csr_decoded_hi_hi_2 ={ core_csr_decoded_hi_hi_hi_2 , core_csr_decoded_andMatrixInput_2_3 }; 
    wire[4:0] core_csr_decoded_hi_3 ={ core_csr_decoded_hi_hi_2 , core_csr_decoded_hi_lo_2 }; 
    wire core_csr_decoded_andMatrixInput_0_4 = core_csr_decoded_plaInput [22]; 
    wire core_csr_decoded_andMatrixInput_1_4 = core_csr_decoded_invInputs [23]; 
    wire core_csr_decoded_andMatrixInput_2_4 = core_csr_decoded_invInputs [24]; 
    wire core_csr_decoded_andMatrixInput_3_4 = core_csr_decoded_invInputs [25]; 
    wire core_csr_decoded_andMatrixInput_4_3 = core_csr_decoded_invInputs [26]; 
    wire core_csr_decoded_andMatrixInput_5_3 = core_csr_decoded_invInputs [27]; 
    wire core_csr_decoded_andMatrixInput_6_3 = core_csr_decoded_plaInput [28]; 
    wire core_csr_decoded_andMatrixInput_7_3 = core_csr_decoded_plaInput [29]; 
    wire core_csr_decoded_andMatrixInput_8_3 = core_csr_decoded_invInputs [30]; 
    wire core_csr_decoded_andMatrixInput_9_3 = core_csr_decoded_invInputs [31]; 
    wire[1:0] core_csr_decoded_lo_lo_3 ={ core_csr_decoded_andMatrixInput_8_3 , core_csr_decoded_andMatrixInput_9_3 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_3 ={ core_csr_decoded_andMatrixInput_5_3 , core_csr_decoded_andMatrixInput_6_3 }; 
    wire[2:0] core_csr_decoded_lo_hi_3 ={ core_csr_decoded_lo_hi_hi_3 , core_csr_decoded_andMatrixInput_7_3 }; 
    wire[4:0] core_csr_decoded_lo_4 ={ core_csr_decoded_lo_hi_3 , core_csr_decoded_lo_lo_3 }; 
    wire[1:0] core_csr_decoded_hi_lo_3 ={ core_csr_decoded_andMatrixInput_3_4 , core_csr_decoded_andMatrixInput_4_3 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_3 ={ core_csr_decoded_andMatrixInput_0_4 , core_csr_decoded_andMatrixInput_1_4 }; 
    wire[2:0] core_csr_decoded_hi_hi_3 ={ core_csr_decoded_hi_hi_hi_3 , core_csr_decoded_andMatrixInput_2_4 }; 
    wire[4:0] core_csr_decoded_hi_4 ={ core_csr_decoded_hi_hi_3 , core_csr_decoded_hi_lo_3 }; 
    wire core_csr_decoded_andMatrixInput_0_5 = core_csr_decoded_plaInput [30]; 
    wire core_csr_decoded_andMatrixInput_1_5 = core_csr_decoded_invInputs [31]; 
    wire[3:0] core_csr_decoded_orMatrixOutputs_lo ={ core_csr_decoded_orMatrixOutputs_lo_hi , core_csr_decoded_orMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_lo ={|(&{ core_csr_decoded_hi_4 , core_csr_decoded_lo_4 }),|(&{ core_csr_decoded_hi_2 , core_csr_decoded_lo_2 })}; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_hi_hi ={|(&{ core_csr_decoded_hi , core_csr_decoded_lo }),|(&{ core_csr_decoded_hi_1 , core_csr_decoded_lo_1 })}; 
    wire[2:0] core_csr_decoded_orMatrixOutputs_hi_hi ={ core_csr_decoded_orMatrixOutputs_hi_hi_hi ,|{&{ core_csr_decoded_hi_3 , core_csr_decoded_lo_3 },&{ core_csr_decoded_andMatrixInput_0_5 , core_csr_decoded_andMatrixInput_1_5 }}}; 
    wire[4:0] core_csr_decoded_orMatrixOutputs_hi ={ core_csr_decoded_orMatrixOutputs_hi_hi , core_csr_decoded_orMatrixOutputs_hi_lo }; 
    wire[8:0] core_csr_decoded_orMatrixOutputs ={ core_csr_decoded_orMatrixOutputs_hi , core_csr_decoded_orMatrixOutputs_lo }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_lo ={ core_csr_decoded_orMatrixOutputs [1], core_csr_decoded_orMatrixOutputs [0]}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_hi ={ core_csr_decoded_orMatrixOutputs [3], core_csr_decoded_orMatrixOutputs [2]}; 
    wire[3:0] core_csr_decoded_invMatrixOutputs_lo ={ core_csr_decoded_invMatrixOutputs_lo_hi , core_csr_decoded_invMatrixOutputs_lo_lo }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_lo ={ core_csr_decoded_orMatrixOutputs [5], core_csr_decoded_orMatrixOutputs [4]}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_hi_hi ={ core_csr_decoded_orMatrixOutputs [8], core_csr_decoded_orMatrixOutputs [7]}; 
    wire[2:0] core_csr_decoded_invMatrixOutputs_hi_hi ={ core_csr_decoded_invMatrixOutputs_hi_hi_hi , core_csr_decoded_orMatrixOutputs [6]}; 
    wire[4:0] core_csr_decoded_invMatrixOutputs_hi ={ core_csr_decoded_invMatrixOutputs_hi_hi , core_csr_decoded_invMatrixOutputs_hi_lo }; 
  assign  core_csr_decoded_invMatrixOutputs ={ core_csr_decoded_invMatrixOutputs_hi , core_csr_decoded_invMatrixOutputs_lo }; 
    wire[8:0] core_csr_decoded = core_csr_decoded_invMatrixOutputs ; 
    wire core_csr_insn_call = core_csr_system_insn & core_csr_decoded [8]; 
    wire core_csr_insn_break = core_csr_system_insn & core_csr_decoded [7]; 
    wire core_csr_insn_ret = core_csr_system_insn & core_csr_decoded [6]; 
    wire core_csr_insn_cease = core_csr_system_insn & core_csr_decoded [5]; 
    wire core_csr_insn_wfi = core_csr_system_insn & core_csr_decoded [4]; 
    wire[11:0] core_csr_addr_1 = core_csr_io_decode_0_inst [31:20]; 
    wire[11:0] core_csr_io_decode_0_fp_csr_plaInput = core_csr_addr_1 ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_plaInput = core_csr_addr_1 ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_plaInput_1 = core_csr_addr_1 ; 
    wire[31:0] core_csr_decoded_invInputs_1 =~ core_csr_decoded_plaInput_1 ; 
    wire[8:0] core_csr_decoded_invMatrixOutputs_1 ; 
    wire core_csr_decoded_andMatrixInput_0_6 = core_csr_decoded_invInputs_1 [20]; 
    wire core_csr_decoded_andMatrixInput_1_6 = core_csr_decoded_invInputs_1 [21]; 
    wire core_csr_decoded_andMatrixInput_2_5 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_3_5 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_4_4 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_5_4 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_6_4 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_7_4 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_8_4 = core_csr_decoded_invInputs_1 [28]; 
    wire core_csr_decoded_andMatrixInput_9_4 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_10_2 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_11_2 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_2 ={ core_csr_decoded_andMatrixInput_9_4 , core_csr_decoded_andMatrixInput_10_2 }; 
    wire[2:0] core_csr_decoded_lo_lo_4 ={ core_csr_decoded_lo_lo_hi_2 , core_csr_decoded_andMatrixInput_11_2 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_4 ={ core_csr_decoded_andMatrixInput_6_4 , core_csr_decoded_andMatrixInput_7_4 }; 
    wire[2:0] core_csr_decoded_lo_hi_4 ={ core_csr_decoded_lo_hi_hi_4 , core_csr_decoded_andMatrixInput_8_4 }; 
    wire[5:0] core_csr_decoded_lo_5 ={ core_csr_decoded_lo_hi_4 , core_csr_decoded_lo_lo_4 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_2 ={ core_csr_decoded_andMatrixInput_3_5 , core_csr_decoded_andMatrixInput_4_4 }; 
    wire[2:0] core_csr_decoded_hi_lo_4 ={ core_csr_decoded_hi_lo_hi_2 , core_csr_decoded_andMatrixInput_5_4 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_4 ={ core_csr_decoded_andMatrixInput_0_6 , core_csr_decoded_andMatrixInput_1_6 }; 
    wire[2:0] core_csr_decoded_hi_hi_4 ={ core_csr_decoded_hi_hi_hi_4 , core_csr_decoded_andMatrixInput_2_5 }; 
    wire[5:0] core_csr_decoded_hi_5 ={ core_csr_decoded_hi_hi_4 , core_csr_decoded_hi_lo_4 }; 
    wire core_csr_decoded_andMatrixInput_0_7 = core_csr_decoded_plaInput_1 [20]; 
    wire core_csr_decoded_andMatrixInput_1_7 = core_csr_decoded_invInputs_1 [21]; 
    wire core_csr_decoded_andMatrixInput_2_6 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_3_6 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_4_5 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_5_5 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_6_5 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_7_5 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_8_5 = core_csr_decoded_invInputs_1 [28]; 
    wire core_csr_decoded_andMatrixInput_9_5 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_10_3 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_11_3 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_lo_hi_3 ={ core_csr_decoded_andMatrixInput_9_5 , core_csr_decoded_andMatrixInput_10_3 }; 
    wire[2:0] core_csr_decoded_lo_lo_5 ={ core_csr_decoded_lo_lo_hi_3 , core_csr_decoded_andMatrixInput_11_3 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_5 ={ core_csr_decoded_andMatrixInput_6_5 , core_csr_decoded_andMatrixInput_7_5 }; 
    wire[2:0] core_csr_decoded_lo_hi_5 ={ core_csr_decoded_lo_hi_hi_5 , core_csr_decoded_andMatrixInput_8_5 }; 
    wire[5:0] core_csr_decoded_lo_6 ={ core_csr_decoded_lo_hi_5 , core_csr_decoded_lo_lo_5 }; 
    wire[1:0] core_csr_decoded_hi_lo_hi_3 ={ core_csr_decoded_andMatrixInput_3_6 , core_csr_decoded_andMatrixInput_4_5 }; 
    wire[2:0] core_csr_decoded_hi_lo_5 ={ core_csr_decoded_hi_lo_hi_3 , core_csr_decoded_andMatrixInput_5_5 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_5 ={ core_csr_decoded_andMatrixInput_0_7 , core_csr_decoded_andMatrixInput_1_7 }; 
    wire[2:0] core_csr_decoded_hi_hi_5 ={ core_csr_decoded_hi_hi_hi_5 , core_csr_decoded_andMatrixInput_2_6 }; 
    wire[5:0] core_csr_decoded_hi_6 ={ core_csr_decoded_hi_hi_5 , core_csr_decoded_hi_lo_5 }; 
    wire core_csr_decoded_andMatrixInput_0_8 = core_csr_decoded_plaInput_1 [28]; 
    wire core_csr_decoded_andMatrixInput_1_8 = core_csr_decoded_invInputs_1 [29]; 
    wire core_csr_decoded_andMatrixInput_2_7 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_3_7 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_7 ={ core_csr_decoded_andMatrixInput_2_7 , core_csr_decoded_andMatrixInput_3_7 }; 
    wire[1:0] core_csr_decoded_hi_7 ={ core_csr_decoded_andMatrixInput_0_8 , core_csr_decoded_andMatrixInput_1_8 }; 
    wire core_csr_decoded_andMatrixInput_0_9 = core_csr_decoded_invInputs_1 [22]; 
    wire core_csr_decoded_andMatrixInput_1_9 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_2_8 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_3_8 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_4_6 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_5_6 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_6_6 = core_csr_decoded_plaInput_1 [28]; 
    wire core_csr_decoded_andMatrixInput_7_6 = core_csr_decoded_plaInput_1 [29]; 
    wire core_csr_decoded_andMatrixInput_8_6 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_9_6 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_lo_6 ={ core_csr_decoded_andMatrixInput_8_6 , core_csr_decoded_andMatrixInput_9_6 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_6 ={ core_csr_decoded_andMatrixInput_5_6 , core_csr_decoded_andMatrixInput_6_6 }; 
    wire[2:0] core_csr_decoded_lo_hi_6 ={ core_csr_decoded_lo_hi_hi_6 , core_csr_decoded_andMatrixInput_7_6 }; 
    wire[4:0] core_csr_decoded_lo_8 ={ core_csr_decoded_lo_hi_6 , core_csr_decoded_lo_lo_6 }; 
    wire[1:0] core_csr_decoded_hi_lo_6 ={ core_csr_decoded_andMatrixInput_3_8 , core_csr_decoded_andMatrixInput_4_6 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_6 ={ core_csr_decoded_andMatrixInput_0_9 , core_csr_decoded_andMatrixInput_1_9 }; 
    wire[2:0] core_csr_decoded_hi_hi_6 ={ core_csr_decoded_hi_hi_hi_6 , core_csr_decoded_andMatrixInput_2_8 }; 
    wire[4:0] core_csr_decoded_hi_8 ={ core_csr_decoded_hi_hi_6 , core_csr_decoded_hi_lo_6 }; 
    wire core_csr_decoded_andMatrixInput_0_10 = core_csr_decoded_plaInput_1 [22]; 
    wire core_csr_decoded_andMatrixInput_1_10 = core_csr_decoded_invInputs_1 [23]; 
    wire core_csr_decoded_andMatrixInput_2_9 = core_csr_decoded_invInputs_1 [24]; 
    wire core_csr_decoded_andMatrixInput_3_9 = core_csr_decoded_invInputs_1 [25]; 
    wire core_csr_decoded_andMatrixInput_4_7 = core_csr_decoded_invInputs_1 [26]; 
    wire core_csr_decoded_andMatrixInput_5_7 = core_csr_decoded_invInputs_1 [27]; 
    wire core_csr_decoded_andMatrixInput_6_7 = core_csr_decoded_plaInput_1 [28]; 
    wire core_csr_decoded_andMatrixInput_7_7 = core_csr_decoded_plaInput_1 [29]; 
    wire core_csr_decoded_andMatrixInput_8_7 = core_csr_decoded_invInputs_1 [30]; 
    wire core_csr_decoded_andMatrixInput_9_7 = core_csr_decoded_invInputs_1 [31]; 
    wire[1:0] core_csr_decoded_lo_lo_7 ={ core_csr_decoded_andMatrixInput_8_7 , core_csr_decoded_andMatrixInput_9_7 }; 
    wire[1:0] core_csr_decoded_lo_hi_hi_7 ={ core_csr_decoded_andMatrixInput_5_7 , core_csr_decoded_andMatrixInput_6_7 }; 
    wire[2:0] core_csr_decoded_lo_hi_7 ={ core_csr_decoded_lo_hi_hi_7 , core_csr_decoded_andMatrixInput_7_7 }; 
    wire[4:0] core_csr_decoded_lo_9 ={ core_csr_decoded_lo_hi_7 , core_csr_decoded_lo_lo_7 }; 
    wire[1:0] core_csr_decoded_hi_lo_7 ={ core_csr_decoded_andMatrixInput_3_9 , core_csr_decoded_andMatrixInput_4_7 }; 
    wire[1:0] core_csr_decoded_hi_hi_hi_7 ={ core_csr_decoded_andMatrixInput_0_10 , core_csr_decoded_andMatrixInput_1_10 }; 
    wire[2:0] core_csr_decoded_hi_hi_7 ={ core_csr_decoded_hi_hi_hi_7 , core_csr_decoded_andMatrixInput_2_9 }; 
    wire[4:0] core_csr_decoded_hi_9 ={ core_csr_decoded_hi_hi_7 , core_csr_decoded_hi_lo_7 }; 
    wire core_csr_decoded_andMatrixInput_0_11 = core_csr_decoded_plaInput_1 [30]; 
    wire core_csr_decoded_andMatrixInput_1_11 = core_csr_decoded_invInputs_1 [31]; 
    wire[3:0] core_csr_decoded_orMatrixOutputs_lo_1 ={ core_csr_decoded_orMatrixOutputs_lo_hi_1 , core_csr_decoded_orMatrixOutputs_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_lo_1 ={|(&{ core_csr_decoded_hi_9 , core_csr_decoded_lo_9 }),|(&{ core_csr_decoded_hi_7 , core_csr_decoded_lo_7 })}; 
    wire[1:0] core_csr_decoded_orMatrixOutputs_hi_hi_hi_1 ={|(&{ core_csr_decoded_hi_5 , core_csr_decoded_lo_5 }),|(&{ core_csr_decoded_hi_6 , core_csr_decoded_lo_6 })}; 
    wire[2:0] core_csr_decoded_orMatrixOutputs_hi_hi_1 ={ core_csr_decoded_orMatrixOutputs_hi_hi_hi_1 ,|{&{ core_csr_decoded_hi_8 , core_csr_decoded_lo_8 },&{ core_csr_decoded_andMatrixInput_0_11 , core_csr_decoded_andMatrixInput_1_11 }}}; 
    wire[4:0] core_csr_decoded_orMatrixOutputs_hi_1 ={ core_csr_decoded_orMatrixOutputs_hi_hi_1 , core_csr_decoded_orMatrixOutputs_hi_lo_1 }; 
    wire[8:0] core_csr_decoded_orMatrixOutputs_1 ={ core_csr_decoded_orMatrixOutputs_hi_1 , core_csr_decoded_orMatrixOutputs_lo_1 }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_lo_1 ={ core_csr_decoded_orMatrixOutputs_1 [1], core_csr_decoded_orMatrixOutputs_1 [0]}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_lo_hi_1 ={ core_csr_decoded_orMatrixOutputs_1 [3], core_csr_decoded_orMatrixOutputs_1 [2]}; 
    wire[3:0] core_csr_decoded_invMatrixOutputs_lo_1 ={ core_csr_decoded_invMatrixOutputs_lo_hi_1 , core_csr_decoded_invMatrixOutputs_lo_lo_1 }; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_lo_1 ={ core_csr_decoded_orMatrixOutputs_1 [5], core_csr_decoded_orMatrixOutputs_1 [4]}; 
    wire[1:0] core_csr_decoded_invMatrixOutputs_hi_hi_hi_1 ={ core_csr_decoded_orMatrixOutputs_1 [8], core_csr_decoded_orMatrixOutputs_1 [7]}; 
    wire[2:0] core_csr_decoded_invMatrixOutputs_hi_hi_1 ={ core_csr_decoded_invMatrixOutputs_hi_hi_hi_1 , core_csr_decoded_orMatrixOutputs_1 [6]}; 
    wire[4:0] core_csr_decoded_invMatrixOutputs_hi_1 ={ core_csr_decoded_invMatrixOutputs_hi_hi_1 , core_csr_decoded_invMatrixOutputs_hi_lo_1 }; 
  assign  core_csr_decoded_invMatrixOutputs_1 ={ core_csr_decoded_invMatrixOutputs_hi_1 , core_csr_decoded_invMatrixOutputs_lo_1 }; 
    wire[8:0] core_csr_decoded_132 = core_csr_decoded_invMatrixOutputs_1 ; 
    wire core_csr_is_break = core_csr_decoded_132 [7]; 
    wire core_csr_is_ret = core_csr_decoded_132 [6]; 
    wire core_csr_is_wfi = core_csr_decoded_132 [4]; 
    wire core_csr_is_sfence = core_csr_decoded_132 [3]; 
    wire core_csr_is_hfence_vvma = core_csr_decoded_132 [2]; 
    wire core_csr_is_hfence_gvma = core_csr_decoded_132 [1]; 
    wire core_csr_is_hlsv = core_csr_decoded_132 [0]; 
    wire core_csr_is_counter = core_csr_addr_1 >=12'hC00& core_csr_addr_1 <12'hC20| core_csr_addr_1 >=12'hC80& core_csr_addr_1 <12'hCA0; 
    wire[4:0] core_csr_counter_addr = core_csr_addr_1 [4:0]; 
    wire[31:0] core_csr__GEN_31 = core_csr_read_mcounteren >> core_csr_counter_addr ; 
    wire core_csr_allow_counter = core_csr_reg_mstatus_prv >2'h1| core_csr__GEN_31 [0]; 
    wire[31:0] core_csr__GEN_32 = core_csr_read_scounteren >> core_csr_counter_addr ; 
    wire[31:0] core_csr__GEN_33 = core_csr_read_hcounteren >> core_csr_counter_addr ; 
    wire core_csr__io_decode_0_fp_illegal_output = core_csr__io_status_fs_output ==2'h0| core_csr_reg_mstatus_v & core_csr_reg_vsstatus_fs ==2'h0| core_csr_reg_misa [5]==1'h0; 
    wire core_csr__io_decode_0_vector_illegal_output = core_csr__io_status_vs_output ==2'h0| core_csr_reg_mstatus_v & core_csr_reg_vsstatus_vs ==2'h0| core_csr_reg_misa [21]==1'h0; 
    wire[11:0] core_csr_io_decode_0_fp_csr_invInputs =~ core_csr_io_decode_0_fp_csr_plaInput ; 
    wire core_csr__io_decode_0_fp_csr_output = core_csr_io_decode_0_fp_csr_plaOutput ; 
    wire core_csr_csr_addr_legal = core_csr_reg_mstatus_prv >= core_csr_addr_1 [9:8]; 
    wire core_csr__GEN_34 = core_csr_addr_1 ==12'h7A0| core_csr_addr_1 ==12'h7A1| core_csr_addr_1 ==12'h7A2| core_csr_addr_1 ==12'h7A3| core_csr_addr_1 ==12'h301| core_csr_addr_1 ==12'h300| core_csr_addr_1 ==12'h305| core_csr_addr_1 ==12'h344| core_csr_addr_1 ==12'h304| core_csr_addr_1 ==12'h340| core_csr_addr_1 ==12'h341| core_csr_addr_1 ==12'h343| core_csr_addr_1 ==12'h342| core_csr_addr_1 ==12'hF14| core_csr_addr_1 ==12'h7B0| core_csr_addr_1 ==12'h7B1| core_csr_addr_1 ==12'h7B2| core_csr_addr_1 ==12'h320| core_csr_addr_1 ==12'hB00| core_csr_addr_1 ==12'hB02| core_csr_addr_1 ==12'h323| core_csr_addr_1 ==12'hB03| core_csr_addr_1 ==12'hC03| core_csr_addr_1 ==12'h324| core_csr_addr_1 ==12'hB04| core_csr_addr_1 ==12'hC04| core_csr_addr_1 ==12'h325| core_csr_addr_1 ==12'hB05| core_csr_addr_1 ==12'hC05| core_csr_addr_1 ==12'h326| core_csr_addr_1 ==12'hB06| core_csr_addr_1 ==12'hC06| core_csr_addr_1 ==12'h327| core_csr_addr_1 ==12'hB07| core_csr_addr_1 ==12'hC07| core_csr_addr_1 ==12'h328| core_csr_addr_1 ==12'hB08| core_csr_addr_1 ==12'hC08| core_csr_addr_1 ==12'h329| core_csr_addr_1 ==12'hB09| core_csr_addr_1 ==12'hC09| core_csr_addr_1 ==12'h32A| core_csr_addr_1 ==12'hB0A| core_csr_addr_1 ==12'hC0A| core_csr_addr_1 ==12'h32B| core_csr_addr_1 ==12'hB0B| core_csr_addr_1 ==12'hC0B| core_csr_addr_1 ==12'h32C| core_csr_addr_1 ==12'hB0C| core_csr_addr_1 ==12'hC0C| core_csr_addr_1 ==12'h32D| core_csr_addr_1 ==12'hB0D| core_csr_addr_1 ==12'hC0D| core_csr_addr_1 ==12'h32E| core_csr_addr_1 ==12'hB0E| core_csr_addr_1 ==12'hC0E| core_csr_addr_1 ==12'h32F| core_csr_addr_1 ==12'hB0F| core_csr_addr_1 ==12'hC0F| core_csr_addr_1 ==12'h330| core_csr_addr_1 ==12'hB10| core_csr_addr_1 ==12'hC10| core_csr_addr_1 ==12'h331| core_csr_addr_1 ==12'hB11| core_csr_addr_1 ==12'hC11| core_csr_addr_1 ==12'h332| core_csr_addr_1 ==12'hB12| core_csr_addr_1 ==12'hC12| core_csr_addr_1 ==12'h333| core_csr_addr_1 ==12'hB13| core_csr_addr_1 ==12'hC13| core_csr_addr_1 ==12'h334| core_csr_addr_1 ==12'hB14| core_csr_addr_1 ==12'hC14| core_csr_addr_1 ==12'h335| core_csr_addr_1 ==12'hB15| core_csr_addr_1 ==12'hC15| core_csr_addr_1 ==12'h336| core_csr_addr_1 ==12'hB16| core_csr_addr_1 ==12'hC16| core_csr_addr_1 ==12'h337| core_csr_addr_1 ==12'hB17| core_csr_addr_1 ==12'hC17| core_csr_addr_1 ==12'h338| core_csr_addr_1 ==12'hB18| core_csr_addr_1 ==12'hC18| core_csr_addr_1 ==12'h339| core_csr_addr_1 ==12'hB19| core_csr_addr_1 ==12'hC19| core_csr_addr_1 ==12'h33A| core_csr_addr_1 ==12'hB1A| core_csr_addr_1 ==12'hC1A| core_csr_addr_1 ==12'h33B| core_csr_addr_1 ==12'hB1B| core_csr_addr_1 ==12'hC1B| core_csr_addr_1 ==12'h33C| core_csr_addr_1 ==12'hB1C| core_csr_addr_1 ==12'hC1C| core_csr_addr_1 ==12'h33D| core_csr_addr_1 ==12'hB1D| core_csr_addr_1 ==12'hC1D| core_csr_addr_1 ==12'h33E| core_csr_addr_1 ==12'hB1E| core_csr_addr_1 ==12'hC1E| core_csr_addr_1 ==12'h33F| core_csr_addr_1 ==12'hB1F| core_csr_addr_1 ==12'hC1F| core_csr_addr_1 ==12'hC00| core_csr_addr_1 ==12'hC02| core_csr_addr_1 ==12'h3A0| core_csr_addr_1 ==12'h3A2| core_csr_addr_1 ==12'h3B0| core_csr_addr_1 ==12'h3B1| core_csr_addr_1 ==12'h3B2| core_csr_addr_1 ==12'h3B3| core_csr_addr_1 ==12'h3B4| core_csr_addr_1 ==12'h3B5| core_csr_addr_1 ==12'h3B6| core_csr_addr_1 ==12'h3B7| core_csr_addr_1 ==12'h3B8| core_csr_addr_1 ==12'h3B9| core_csr_addr_1 ==12'h3BA| core_csr_addr_1 ==12'h3BB| core_csr_addr_1 ==12'h3BC| core_csr_addr_1 ==12'h3BD| core_csr_addr_1 ==12'h3BE| core_csr_addr_1 ==12'h3BF| core_csr_addr_1 ==12'h7C1| core_csr_addr_1 ==12'hF12; 
    wire core_csr_csr_exists = core_csr__GEN_34 | core_csr_addr_1 ==12'hF11| core_csr_addr_1 ==12'hF13| core_csr_addr_1 ==12'hF15; 
    wire[11:0] core_csr_io_decode_0_read_illegal_invInputs =~ core_csr_io_decode_0_read_illegal_plaInput ; 
    wire core_csr_io_decode_0_read_illegal_invMatrixOutputs ; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_0 = core_csr_io_decode_0_read_illegal_plaInput [4]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_1 = core_csr_io_decode_0_read_illegal_plaInput [5]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_2 = core_csr_io_decode_0_read_illegal_invInputs [6]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_3 = core_csr_io_decode_0_read_illegal_plaInput [7]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_4 = core_csr_io_decode_0_read_illegal_plaInput [8]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_5 = core_csr_io_decode_0_read_illegal_plaInput [9]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_6 = core_csr_io_decode_0_read_illegal_plaInput [10]; 
    wire core_csr_io_decode_0_read_illegal_andMatrixInput_7 = core_csr_io_decode_0_read_illegal_invInputs [11]; 
    wire[1:0] core_csr_io_decode_0_read_illegal_lo_lo ={ core_csr_io_decode_0_read_illegal_andMatrixInput_6 , core_csr_io_decode_0_read_illegal_andMatrixInput_7 }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_lo_hi ={ core_csr_io_decode_0_read_illegal_andMatrixInput_4 , core_csr_io_decode_0_read_illegal_andMatrixInput_5 }; 
    wire[3:0] core_csr_io_decode_0_read_illegal_lo ={ core_csr_io_decode_0_read_illegal_lo_hi , core_csr_io_decode_0_read_illegal_lo_lo }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_hi_lo ={ core_csr_io_decode_0_read_illegal_andMatrixInput_2 , core_csr_io_decode_0_read_illegal_andMatrixInput_3 }; 
    wire[1:0] core_csr_io_decode_0_read_illegal_hi_hi ={ core_csr_io_decode_0_read_illegal_andMatrixInput_0 , core_csr_io_decode_0_read_illegal_andMatrixInput_1 }; 
    wire[3:0] core_csr_io_decode_0_read_illegal_hi ={ core_csr_io_decode_0_read_illegal_hi_hi , core_csr_io_decode_0_read_illegal_hi_lo }; 
    wire core_csr_io_decode_0_read_illegal_orMatrixOutputs =|(&{ core_csr_io_decode_0_read_illegal_hi , core_csr_io_decode_0_read_illegal_lo }); 
  assign  core_csr_io_decode_0_read_illegal_invMatrixOutputs = core_csr_io_decode_0_read_illegal_orMatrixOutputs ; 
    wire core_csr_io_decode_0_read_illegal_plaOutput = core_csr_io_decode_0_read_illegal_invMatrixOutputs ; 
    wire[11:0] core_csr_io_decode_0_read_illegal_invInputs_1 =~ core_csr_io_decode_0_read_illegal_plaInput_1 ; 
    wire[11:0] core_csr_io_decode_0_write_flush_addr_m = core_csr_addr_1 |12'h300; 
    wire[31:0] core_csr__GEN_35 = core_csr_read_mcounteren >> core_csr_counter_addr ; 
    wire[31:0] core_csr__GEN_36 = core_csr_read_hcounteren >> core_csr_counter_addr ; 
    wire[31:0] core_csr__GEN_37 = core_csr_read_scounteren >> core_csr_counter_addr ; 
    wire[4:0] core_csr__GEN_38 ={3'h0, core_csr_reg_mstatus_prv [0]& core_csr_reg_mstatus_v  ? 2'h2: core_csr_reg_mstatus_prv }+5'h8; 
    wire[63:0] core_csr_cause = core_csr_insn_call  ? {60'h0, core_csr__GEN_38 [3:0]}: core_csr_insn_break  ? 64'h3: core_csr_io_cause ; 
    wire[7:0] core_csr_cause_lsbs = core_csr_cause [7:0]; 
    wire core_csr_causeIsDebugInt = core_csr_cause [63]& core_csr_cause_lsbs ==8'hE; 
    wire core_csr_causeIsDebugTrigger = core_csr_cause [63]==1'h0& core_csr_cause_lsbs ==8'hE; 
    wire[1:0] core_csr_causeIsDebugBreak_lo ={ core_csr_reg_dcsr_ebreaks , core_csr_reg_dcsr_ebreaku }; 
    wire[1:0] core_csr_causeIsDebugBreak_hi ={ core_csr_reg_dcsr_ebreakm , core_csr_reg_dcsr_ebreakh }; 
    wire[3:0] core_csr__GEN_39 ={ core_csr_causeIsDebugBreak_hi , core_csr_causeIsDebugBreak_lo }>> core_csr_reg_mstatus_prv ; 
    wire core_csr_causeIsDebugBreak = core_csr_cause [63]==1'h0& core_csr_insn_break & core_csr__GEN_39 [0]; 
    wire core_csr_trapToDebug =( core_csr_reg_singleStepped | core_csr_causeIsDebugInt | core_csr_causeIsDebugTrigger | core_csr_causeIsDebugBreak | core_csr_reg_debug )&1'h1; 
    wire[11:0] core_csr_debugTVec = core_csr_reg_debug  ? ( core_csr_insn_break  ? 12'h800:12'h808):12'h800; 
    wire[63:0] core_csr__GEN_40 = core_csr_read_mideleg >> core_csr_cause_lsbs ; 
    wire[63:0] core_csr__GEN_41 = core_csr_read_medeleg >> core_csr_cause_lsbs ; 
    wire[63:0] core_csr__GEN_42 = core_csr_read_hideleg >> core_csr_cause_lsbs ; 
    wire[63:0] core_csr__GEN_43 = core_csr_read_hedeleg >> core_csr_cause_lsbs ; 
    wire core_csr_delegateVS = core_csr_reg_mstatus_v & core_csr_delegate &( core_csr_cause [63] ?  core_csr__GEN_42 [0]: core_csr__GEN_43 [0]); 
    wire[63:0] core_csr_notDebugTVec_base = core_csr_delegate  ? ( core_csr_delegateVS  ?  core_csr_read_vstvec : core_csr_read_stvec ): core_csr_read_mtvec ; 
    wire[7:0] core_csr_notDebugTVec_interruptOffset ={ core_csr_cause [5:0],2'h0}; 
    wire[63:0] core_csr_notDebugTVec_interruptVec ={ core_csr_notDebugTVec_base [63:8], core_csr_notDebugTVec_interruptOffset }; 
    wire core_csr_notDebugTVec_doVector = core_csr_notDebugTVec_base [0]& core_csr_cause [63]& core_csr_cause_lsbs [7:6]==2'h0; 
    wire[63:0] core_csr_notDebugTVec = core_csr_notDebugTVec_doVector  ?  core_csr_notDebugTVec_interruptVec :{ core_csr_notDebugTVec_base [63:2],2'h0}; 
    wire core_csr_causeIsRnmiInt = core_csr_cause [63]& core_csr_cause [62]&( core_csr_cause_lsbs ==8'hD| core_csr_cause_lsbs ==8'hC); 
    wire core_csr_causeIsRnmiBEU = core_csr_cause [63]& core_csr_cause [62]& core_csr_cause_lsbs ==8'hC; 
    wire core_csr_trapToNmi = core_csr_trapToNmiInt | core_csr_trapToNmiXcpt ; 
    wire[63:0] core_csr_tvec = core_csr_trapToDebug  ? {52'h0, core_csr_debugTVec }: core_csr_trapToNmi  ? {62'h0, core_csr_nmiTVec }: core_csr_notDebugTVec ; 
  assign  core_csr__io_singleStep_output = core_csr_reg_dcsr_step & core_csr_reg_debug ==1'h0; 
  assign  core_csr__io_status_sd_output =(& core_csr__io_status_fs_output )|(& core_csr__io_status_xs_output )|(& core_csr__io_status_vs_output ); 
  assign  core_csr__io_status_isa_output = core_csr_reg_misa [31:0]; 
  assign  core_csr__io_status_dprv_output = core_csr_reg_mstatus_mprv & core_csr_reg_debug ==1'h0 ?  core_csr_reg_mstatus_mpp : core_csr_reg_mstatus_prv ; 
  assign  core_csr__io_status_dv_output = core_csr_reg_mstatus_v |( core_csr_reg_mstatus_mprv & core_csr_reg_debug ==1'h0 ?  core_csr_reg_mstatus_mpv :1'h0); 
    wire core_csr__io_gstatus_sd_output =(& core_csr__io_gstatus_fs_output )|(& core_csr__io_gstatus_xs_output )|(& core_csr__io_gstatus_vs_output ); 
    wire core_csr_exception = core_csr_insn_call | core_csr_insn_break | core_csr_io_exception ; 
    wire core_csr__GEN_44 ={1'h0,{1'h0, core_csr_insn_ret }+{1'h0, core_csr_insn_call }}+{1'h0,{1'h0, core_csr_insn_break }+{1'h0, core_csr_io_exception }}<=3'h1==1'h0; 
    wire core_csr__GEN_45 = core_csr_insn_wfi & core_csr__io_singleStep_output ==1'h0& core_csr_reg_debug ==1'h0; 
    wire core_csr__GEN_46 =(| core_csr_pending_interrupts )| core_csr_io_interrupts_debug | core_csr_exception ; 
    wire core_csr__GEN_47 = core_csr_io_retire | core_csr_exception ; 
    wire core_csr__GEN_48 = core_csr__io_singleStep_output ==1'h0; 
    wire core_csr__GEN_49 =( core_csr__io_singleStep_output ==1'h0| core_csr_io_retire <=1'h1)==1'h0; 
    wire core_csr__GEN_50 =( core_csr_reg_singleStepped ==1'h0| core_csr_io_retire ==1'h0)==1'h0; 
  always @( posedge  core_csr_clock )
         begin 
             if ( core_csr_reset ==1'h0& core_csr__GEN_44 )
                 begin 
                     if (1)$error("Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:1010 assert(PopCount(insn_ret :: insn_call :: insn_break :: io.exception :: Nil) <= 1.U, \"these conditions must be mutually exclusive\")\n");
                     if (1)$fatal;
                 end 
             if ( core_csr_reset ==1'h0& core_csr__GEN_49 )
                 begin 
                     if (1)$error("Assertion failed\n    at CSR.scala:1018 assert(!io.singleStep || io.retire <= 1.U)\n");
                     if (1)$fatal;
                 end 
             if ( core_csr_reset ==1'h0& core_csr__GEN_50 )
                 begin 
                     if (1)$error("Assertion failed\n    at CSR.scala:1019 assert(!reg_singleStepped || io.retire === 0.U)\n");
                     if (1)$fatal;
                 end 
         end
    wire[33:0] core_csr_epc =~(~ core_csr_io_pc |34'h1); 
    wire[33:0] core_csr_tval = core_csr_insn_break  ?  core_csr_epc : core_csr_io_tval ; 
    wire core_csr__GEN_51 = core_csr_reg_debug ==1'h0; 
    wire core_csr__GEN_52 = core_csr_exception  ? ( core_csr_trapToDebug  ? ( core_csr__GEN_51  ? 1'h1: core_csr_reg_debug ): core_csr_reg_debug ): core_csr_reg_debug ; 
    wire[33:0] core_csr__GEN_53 = core_csr_exception  ? ( core_csr_trapToDebug  ? ( core_csr__GEN_51  ?  core_csr_epc : core_csr_reg_dpc ): core_csr_reg_dpc ): core_csr_reg_dpc ; 
    wire[2:0] core_csr__GEN_54 = core_csr_reg_singleStepped  ? 3'h4:{1'h0, core_csr_causeIsDebugInt  ? 2'h3: core_csr_causeIsDebugTrigger  ? 2'h2:2'h1}; 
    wire core_csr__GEN_55 = core_csr_exception &~ core_csr_trapToDebug ; 
    wire[63:0] core_csr__GEN_56 ={62'h0, core_csr_causeIsRnmiBEU  ? 2'h3:2'h2}|64'h8000000000000000; 
    wire core_csr__GEN_57 = core_csr__GEN_55 &~ core_csr_trapToNmiInt ; 
    wire core_csr__GEN_58 = core_csr_delegateVS & core_csr_reg_rnmie ; 
    wire[63:0] core_csr__GEN_59 = core_csr_cause [63] ? { core_csr_cause [63:2],2'h1}: core_csr_cause ; 
    wire core_csr__GEN_60 = core_csr__GEN_57 &~ core_csr__GEN_58 ; 
    wire core_csr__GEN_61 = core_csr_delegate & core_csr_reg_rnmie ; 
    wire core_csr__GEN_62 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mstatus_mpv : core_csr_trapToNmiInt  ?  core_csr_reg_mstatus_mpv : core_csr__GEN_58  ?  core_csr_reg_mstatus_mpv : core_csr__GEN_61  ?  core_csr_reg_mstatus_mpv : core_csr_reg_mstatus_v ): core_csr_reg_mstatus_mpv ; 
    wire[33:0] core_csr__GEN_63 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mepc : core_csr_trapToNmiInt  ?  core_csr_reg_mepc : core_csr__GEN_58  ?  core_csr_reg_mepc : core_csr__GEN_61  ?  core_csr_reg_mepc : core_csr_epc ): core_csr_reg_mepc ; 
    wire[63:0] core_csr__GEN_64 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mcause : core_csr_trapToNmiInt  ?  core_csr_reg_mcause : core_csr__GEN_58  ?  core_csr_reg_mcause : core_csr__GEN_61  ?  core_csr_reg_mcause : core_csr_cause ): core_csr_reg_mcause ; 
    wire[33:0] core_csr__GEN_65 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mtval : core_csr_trapToNmiInt  ?  core_csr_reg_mtval : core_csr__GEN_58  ?  core_csr_reg_mtval : core_csr__GEN_61  ?  core_csr_reg_mtval : core_csr_tval ): core_csr_reg_mtval ; 
    wire core_csr__GEN_66 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mstatus_mpie : core_csr_trapToNmiInt  ?  core_csr_reg_mstatus_mpie : core_csr__GEN_58  ?  core_csr_reg_mstatus_mpie : core_csr__GEN_61  ?  core_csr_reg_mstatus_mpie : core_csr_reg_mstatus_mie ): core_csr_reg_mstatus_mpie ; 
    wire[1:0] core_csr__GEN_67 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mstatus_mpp : core_csr_trapToNmiInt  ?  core_csr_reg_mstatus_mpp : core_csr__GEN_58  ?  core_csr_reg_mstatus_mpp : core_csr__GEN_61  ?  core_csr_reg_mstatus_mpp :2'h3): core_csr_reg_mstatus_mpp ; 
    wire core_csr__GEN_68 = core_csr_exception  ? ( core_csr_trapToDebug  ?  core_csr_reg_mstatus_mie : core_csr_trapToNmiInt  ?  core_csr_reg_mstatus_mie : core_csr__GEN_58  ?  core_csr_reg_mstatus_mie : core_csr__GEN_61  ?  core_csr_reg_mstatus_mie :1'h0): core_csr_reg_mstatus_mie ; 
    wire core_csr_en = core_csr_exception &(|( core_csr_supported_interrupts &16'h1))& core_csr_cause ==64'h8000000000000000; 
    wire core_csr_delegable =|( core_csr_delegable_interrupts &16'h1); 
    wire core_csr_en_1 = core_csr_exception &(|( core_csr_supported_interrupts &16'h2))& core_csr_cause ==64'h8000000000000001; 
    wire core_csr_delegable_1 =|( core_csr_delegable_interrupts &16'h2); 
    wire core_csr_en_2 = core_csr_exception &(|( core_csr_supported_interrupts &16'h4))& core_csr_cause ==64'h8000000000000002; 
    wire core_csr_delegable_2 =|( core_csr_delegable_interrupts &16'h4); 
    wire core_csr_en_3 = core_csr_exception &(|( core_csr_supported_interrupts &16'h8))& core_csr_cause ==64'h8000000000000003; 
    wire core_csr_delegable_3 =|( core_csr_delegable_interrupts &16'h8); 
    wire core_csr_en_4 = core_csr_exception &(|( core_csr_supported_interrupts &16'h10))& core_csr_cause ==64'h8000000000000004; 
    wire core_csr_delegable_4 =|( core_csr_delegable_interrupts &16'h10); 
    wire core_csr_en_5 = core_csr_exception &(|( core_csr_supported_interrupts &16'h20))& core_csr_cause ==64'h8000000000000005; 
    wire core_csr_delegable_5 =|( core_csr_delegable_interrupts &16'h20); 
    wire core_csr_en_6 = core_csr_exception &(|( core_csr_supported_interrupts &16'h40))& core_csr_cause ==64'h8000000000000006; 
    wire core_csr_delegable_6 =|( core_csr_delegable_interrupts &16'h40); 
    wire core_csr_en_7 = core_csr_exception &(|( core_csr_supported_interrupts &16'h80))& core_csr_cause ==64'h8000000000000007; 
    wire core_csr_delegable_7 =|( core_csr_delegable_interrupts &16'h80); 
    wire core_csr_en_8 = core_csr_exception &(|( core_csr_supported_interrupts &16'h100))& core_csr_cause ==64'h8000000000000008; 
    wire core_csr_delegable_8 =|( core_csr_delegable_interrupts &16'h100); 
    wire core_csr_en_9 = core_csr_exception &(|( core_csr_supported_interrupts &16'h200))& core_csr_cause ==64'h8000000000000009; 
    wire core_csr_delegable_9 =|( core_csr_delegable_interrupts &16'h200); 
    wire core_csr_en_10 = core_csr_exception &(|( core_csr_supported_interrupts &16'h400))& core_csr_cause ==64'h800000000000000A; 
    wire core_csr_delegable_10 =|( core_csr_delegable_interrupts &16'h400); 
    wire core_csr_en_11 = core_csr_exception &(|( core_csr_supported_interrupts &16'h800))& core_csr_cause ==64'h800000000000000B; 
    wire core_csr_delegable_11 =|( core_csr_delegable_interrupts &16'h800); 
    wire core_csr_en_12 = core_csr_exception &(|( core_csr_supported_interrupts &16'h1000))& core_csr_cause ==64'h800000000000000C; 
    wire core_csr_delegable_12 =|( core_csr_delegable_interrupts &16'h1000); 
    wire core_csr_en_13 = core_csr_exception &(|( core_csr_supported_interrupts &16'h2000))& core_csr_cause ==64'h800000000000000D; 
    wire core_csr_delegable_13 =|( core_csr_delegable_interrupts &16'h2000); 
    wire core_csr_en_14 = core_csr_exception &(|( core_csr_supported_interrupts &16'h4000))& core_csr_cause ==64'h800000000000000E; 
    wire core_csr_delegable_14 =|( core_csr_delegable_interrupts &16'h4000); 
    wire core_csr_en_15 = core_csr_exception &(|( core_csr_supported_interrupts &16'h8000))& core_csr_cause ==64'h800000000000000F; 
    wire core_csr_delegable_15 =|( core_csr_delegable_interrupts &16'h8000); 
    wire core_csr_en_16 = core_csr_exception & core_csr_cause ==64'h0; 
    wire core_csr_en_17 = core_csr_exception & core_csr_cause ==64'h1; 
    wire core_csr_en_18 = core_csr_exception & core_csr_cause ==64'h2; 
    wire core_csr_en_19 = core_csr_exception & core_csr_cause ==64'h3; 
    wire core_csr_en_20 = core_csr_exception & core_csr_cause ==64'h4; 
    wire core_csr_en_21 = core_csr_exception & core_csr_cause ==64'h5; 
    wire core_csr_en_22 = core_csr_exception & core_csr_cause ==64'h6; 
    wire core_csr_en_23 = core_csr_exception & core_csr_cause ==64'h7; 
    wire core_csr_en_24 = core_csr_exception & core_csr_cause ==64'hB; 
    wire core_csr__GEN_69 = core_csr_reg_mstatus_v ==1'h0; 
    wire core_csr__GEN_70 = core_csr_io_rw_addr [10]&1'h1& core_csr_io_rw_addr [7]; 
    wire core_csr__GEN_71 = core_csr_insn_ret  ? ( core_csr__GEN_70  ?  core_csr__GEN_68 : core_csr_reg_mstatus_mpie ): core_csr__GEN_68 ; 
    wire core_csr__GEN_72 = core_csr_insn_ret  ? ( core_csr__GEN_70  ?  core_csr__GEN_66 :1'h1): core_csr__GEN_66 ; 
    wire[1:0] core_csr_ret_prv = core_csr__GEN_70  ?  core_csr_reg_dcsr_prv : core_csr_reg_mstatus_mpp ; 
    wire[1:0] core_csr_new_prv = core_csr_insn_ret  ?  core_csr_ret_prv : core_csr_exception  ? ( core_csr_trapToDebug  ? ( core_csr__GEN_51  ? 2'h3: core_csr_reg_mstatus_prv ): core_csr_trapToNmiInt  ? ( core_csr_reg_rnmie  ? 2'h3: core_csr_reg_mstatus_prv ): core_csr__GEN_58  ? 2'h1: core_csr__GEN_61  ? 2'h1:2'h3): core_csr_reg_mstatus_prv ; 
  assign  core_csr__io_csr_stall_output = core_csr_reg_wfi | core_csr__io_status_cease_output ; 
    reg core_csr_io_status_cease_r ; 
  assign  core_csr__io_status_cease_output = core_csr_io_status_cease_r ; 
  assign  core_csr__io_rw_rdata_WIRE ={63'h0, core_csr_decoded_0  ?  core_csr_reg_tselect :1'h0}|( core_csr_decoded_1  ? { core_csr_hi_4 , core_csr_lo_4 }:64'h0)|( core_csr_decoded_2  ? { core_csr_casez_tmp_314 [32] ? 31'h7FFFFFFF:31'h0, core_csr_casez_tmp_334 }:64'h0)|{13'h0, core_csr_decoded_3  ? { core_csr_hi_5 , core_csr_lo_5 }:51'h0}|( core_csr_decoded_4  ?  core_csr_reg_misa :64'h0)|( core_csr_decoded_5  ?  core_csr_read_mstatus :64'h0)|( core_csr_decoded_6  ?  core_csr_read_mtvec :64'h0)|{48'h0, core_csr_decoded_7  ?  core_csr_read_mip :16'h0}|( core_csr_decoded_8  ?  core_csr_reg_mie :64'h0)|( core_csr_decoded_9  ?  core_csr_reg_mscratch :64'h0)|( core_csr_decoded_10  ? { core_csr__GEN_29 [33] ? 30'h3FFFFFFF:30'h0, core_csr__GEN_29 }:64'h0)|( core_csr_decoded_11  ? { core_csr_reg_mtval [33] ? 30'h3FFFFFFF:30'h0, core_csr_reg_mtval }:64'h0)|( core_csr_decoded_12  ?  core_csr_reg_mcause :64'h0)|{63'h0, core_csr_decoded_13  ?  core_csr_io_hartid :1'h0}|{32'h0, core_csr_decoded_14  ? { core_csr_hi_6 , core_csr_lo_6 }:32'h0}|( core_csr_decoded_15  ? { core_csr__GEN_30 [33] ? 30'h3FFFFFFF:30'h0, core_csr__GEN_30 }:64'h0)|( core_csr_decoded_16  ?  core_csr_reg_dscratch0 :64'h0)|{61'h0, core_csr_decoded_17  ?  core_csr_reg_mcountinhibit :3'h0}|( core_csr_decoded_18  ?  core_csr_value_1 :64'h0)|( core_csr_decoded_19  ?  core_csr_value :64'h0)|( core_csr_decoded_107  ?  core_csr_value_1 :64'h0)|( core_csr_decoded_108  ?  core_csr_value :64'h0)|( core_csr_decoded_109  ? { core_csr_hi_15 , core_csr_lo_15 }:64'h0)|( core_csr_decoded_110  ? { core_csr_hi_24 , core_csr_lo_24 }:64'h0)|{34'h0, core_csr_decoded_111  ?  core_csr_reg_pmp_0_addr :30'h0}|{34'h0, core_csr_decoded_112  ?  core_csr_reg_pmp_1_addr :30'h0}|{34'h0, core_csr_decoded_113  ?  core_csr_reg_pmp_2_addr :30'h0}|{34'h0, core_csr_decoded_114  ?  core_csr_reg_pmp_3_addr :30'h0}|{34'h0, core_csr_decoded_115  ?  core_csr_reg_pmp_4_addr :30'h0}|{34'h0, core_csr_decoded_116  ?  core_csr_reg_pmp_5_addr :30'h0}|{34'h0, core_csr_decoded_117  ?  core_csr_reg_pmp_6_addr :30'h0}|{34'h0, core_csr_decoded_118  ?  core_csr_reg_pmp_7_addr :30'h0}|{34'h0, core_csr_decoded_119  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_120  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_121  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_122  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_123  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_124  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_125  ?  core_csr_read_pmp_15_addr :30'h0}|{34'h0, core_csr_decoded_126  ?  core_csr_read_pmp_15_addr :30'h0}|( core_csr_decoded_127  ?  core_csr_reg_custom_0 :64'h0)|( core_csr_decoded_128  ?  core_csr_reg_custom_1 :64'h0)|( core_csr_decoded_129  ?  core_csr_reg_custom_2 :64'h0)|( core_csr_decoded_130  ?  core_csr_reg_custom_3 :64'h0); 
  assign  core_csr__io_rw_rdata_output = core_csr__io_rw_rdata_WIRE ; 
    wire[4:0] core_csr__GEN_73 = core_csr_reg_fflags | core_csr_io_fcsr_flags_bits ; 
    wire core_csr_csr_wen =( core_csr_io_rw_cmd ==3'h6|(& core_csr_io_rw_cmd )| core_csr_io_rw_cmd ==3'h5)& core_csr__io_rw_stall_output ==1'h0; 
    wire[104:0] core_csr__new_mstatus_WIRE ={41'h0, core_csr_wdata }; 
    wire core_csr_new_mstatus_uie = core_csr__new_mstatus_WIRE [0]; 
    wire core_csr_new_mstatus_sie = core_csr__new_mstatus_WIRE [1]; 
    wire core_csr_new_mstatus_hie = core_csr__new_mstatus_WIRE [2]; 
    wire core_csr_new_mstatus_mie = core_csr__new_mstatus_WIRE [3]; 
    wire core_csr_new_mstatus_upie = core_csr__new_mstatus_WIRE [4]; 
    wire core_csr_new_mstatus_spie = core_csr__new_mstatus_WIRE [5]; 
    wire core_csr_new_mstatus_ube = core_csr__new_mstatus_WIRE [6]; 
    wire core_csr_new_mstatus_mpie = core_csr__new_mstatus_WIRE [7]; 
    wire core_csr_new_mstatus_spp = core_csr__new_mstatus_WIRE [8]; 
    wire[1:0] core_csr_new_mstatus_vs = core_csr__new_mstatus_WIRE [10:9]; 
    wire[1:0] core_csr_new_mstatus_mpp = core_csr__new_mstatus_WIRE [12:11]; 
    wire[1:0] core_csr_new_mstatus_fs = core_csr__new_mstatus_WIRE [14:13]; 
    wire[1:0] core_csr_new_mstatus_xs = core_csr__new_mstatus_WIRE [16:15]; 
    wire core_csr_new_mstatus_mprv = core_csr__new_mstatus_WIRE [17]; 
    wire core_csr_new_mstatus_sum = core_csr__new_mstatus_WIRE [18]; 
    wire core_csr_new_mstatus_mxr = core_csr__new_mstatus_WIRE [19]; 
    wire core_csr_new_mstatus_tvm = core_csr__new_mstatus_WIRE [20]; 
    wire core_csr_new_mstatus_tw = core_csr__new_mstatus_WIRE [21]; 
    wire core_csr_new_mstatus_tsr = core_csr__new_mstatus_WIRE [22]; 
    wire[7:0] core_csr_new_mstatus_zero1 = core_csr__new_mstatus_WIRE [30:23]; 
    wire core_csr_new_mstatus_sd_rv32 = core_csr__new_mstatus_WIRE [31]; 
    wire[1:0] core_csr_new_mstatus_uxl = core_csr__new_mstatus_WIRE [33:32]; 
    wire[1:0] core_csr_new_mstatus_sxl = core_csr__new_mstatus_WIRE [35:34]; 
    wire core_csr_new_mstatus_sbe = core_csr__new_mstatus_WIRE [36]; 
    wire core_csr_new_mstatus_mbe = core_csr__new_mstatus_WIRE [37]; 
    wire core_csr_new_mstatus_gva = core_csr__new_mstatus_WIRE [38]; 
    wire core_csr_new_mstatus_mpv = core_csr__new_mstatus_WIRE [39]; 
    wire[22:0] core_csr_new_mstatus_zero2 = core_csr__new_mstatus_WIRE [62:40]; 
    wire core_csr_new_mstatus_sd = core_csr__new_mstatus_WIRE [63]; 
    wire core_csr_new_mstatus_v = core_csr__new_mstatus_WIRE [64]; 
    wire[1:0] core_csr_new_mstatus_prv = core_csr__new_mstatus_WIRE [66:65]; 
    wire core_csr_new_mstatus_dv = core_csr__new_mstatus_WIRE [67]; 
    wire[1:0] core_csr_new_mstatus_dprv = core_csr__new_mstatus_WIRE [69:68]; 
    wire[31:0] core_csr_new_mstatus_isa = core_csr__new_mstatus_WIRE [101:70]; 
    wire core_csr_new_mstatus_wfi = core_csr__new_mstatus_WIRE [102]; 
    wire core_csr_new_mstatus_cease = core_csr__new_mstatus_WIRE [103]; 
    wire core_csr_new_mstatus_debug = core_csr__new_mstatus_WIRE [104]; 
    wire core_csr_f = core_csr_wdata [5]; 
    wire core_csr__GEN_74 = core_csr_io_pc [1]==1'h0|1'h0| core_csr_wdata [2]; 
    wire[63:0] core_csr__GEN_75 =~(~ core_csr_wdata |{60'h0,{ core_csr_f ==1'h0,3'h0}})&64'h1005| core_csr_reg_misa &64'hFFFFFFFFFFFFEFFA; 
    wire[1:0] core_csr_new_mip_lo_lo_lo ={ core_csr_reg_mip_ssip , core_csr_reg_mip_usip }; 
    wire[1:0] core_csr_new_mip_lo_lo_hi ={ core_csr_reg_mip_msip , core_csr_reg_mip_vssip }; 
    wire[3:0] core_csr_new_mip_lo_lo ={ core_csr_new_mip_lo_lo_hi , core_csr_new_mip_lo_lo_lo }; 
    wire[1:0] core_csr_new_mip_lo_hi_lo ={ core_csr_reg_mip_stip , core_csr_reg_mip_utip }; 
    wire[1:0] core_csr_new_mip_lo_hi_hi ={ core_csr_reg_mip_mtip , core_csr_reg_mip_vstip }; 
    wire[3:0] core_csr_new_mip_lo_hi ={ core_csr_new_mip_lo_hi_hi , core_csr_new_mip_lo_hi_lo }; 
    wire[7:0] core_csr_new_mip_lo ={ core_csr_new_mip_lo_hi , core_csr_new_mip_lo_lo }; 
    wire[1:0] core_csr_new_mip_hi_lo_lo ={ core_csr_reg_mip_seip , core_csr_reg_mip_ueip }; 
    wire[1:0] core_csr_new_mip_hi_lo_hi ={ core_csr_reg_mip_meip , core_csr_reg_mip_vseip }; 
    wire[3:0] core_csr_new_mip_hi_lo ={ core_csr_new_mip_hi_lo_hi , core_csr_new_mip_hi_lo_lo }; 
    wire[1:0] core_csr_new_mip_hi_hi_lo ={ core_csr_reg_mip_rocc , core_csr_reg_mip_sgeip }; 
    wire[1:0] core_csr_new_mip_hi_hi_hi ={ core_csr_reg_mip_zero1 , core_csr_reg_mip_debug }; 
    wire[3:0] core_csr_new_mip_hi_hi ={ core_csr_new_mip_hi_hi_hi , core_csr_new_mip_hi_hi_lo }; 
    wire[7:0] core_csr_new_mip_hi ={ core_csr_new_mip_hi_hi , core_csr_new_mip_hi_lo }; 
    wire[63:0] core_csr__GEN_76 =({48'h0, core_csr_io_rw_cmd [1] ? { core_csr_new_mip_hi , core_csr_new_mip_lo }:16'h0}| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :64'h0); 
    wire[15:0] core_csr__new_mip_WIRE = core_csr__GEN_76 [15:0]; 
    wire core_csr_new_mip_usip = core_csr__new_mip_WIRE [0]; 
    wire core_csr_new_mip_ssip = core_csr__new_mip_WIRE [1]; 
    wire core_csr_new_mip_vssip = core_csr__new_mip_WIRE [2]; 
    wire core_csr_new_mip_msip = core_csr__new_mip_WIRE [3]; 
    wire core_csr_new_mip_utip = core_csr__new_mip_WIRE [4]; 
    wire core_csr_new_mip_stip = core_csr__new_mip_WIRE [5]; 
    wire core_csr_new_mip_vstip = core_csr__new_mip_WIRE [6]; 
    wire core_csr_new_mip_mtip = core_csr__new_mip_WIRE [7]; 
    wire core_csr_new_mip_ueip = core_csr__new_mip_WIRE [8]; 
    wire core_csr_new_mip_seip = core_csr__new_mip_WIRE [9]; 
    wire core_csr_new_mip_vseip = core_csr__new_mip_WIRE [10]; 
    wire core_csr_new_mip_meip = core_csr__new_mip_WIRE [11]; 
    wire core_csr_new_mip_sgeip = core_csr__new_mip_WIRE [12]; 
    wire core_csr_new_mip_rocc = core_csr__new_mip_WIRE [13]; 
    wire core_csr_new_mip_debug = core_csr__new_mip_WIRE [14]; 
    wire core_csr_new_mip_zero1 = core_csr__new_mip_WIRE [15]; 
    wire[63:0] core_csr__GEN_77 = core_csr_wdata &{48'h0, core_csr_supported_interrupts }; 
    wire[63:0] core_csr__GEN_78 =~(~ core_csr_wdata |64'h1); 
    wire[63:0] core_csr__GEN_79 = core_csr_wdata &64'h800000000000000F; 
    wire[63:0] core_csr__GEN_80 = core_csr_wdata &64'hFFFFFFFFFFFFFFFD; 
    wire[31:0] core_csr__new_dcsr_WIRE = core_csr_wdata [31:0]; 
    wire[1:0] core_csr_new_dcsr_prv = core_csr__new_dcsr_WIRE [1:0]; 
    wire core_csr_new_dcsr_step = core_csr__new_dcsr_WIRE [2]; 
    wire[1:0] core_csr_new_dcsr_zero1 = core_csr__new_dcsr_WIRE [4:3]; 
    wire core_csr_new_dcsr_v = core_csr__new_dcsr_WIRE [5]; 
    wire[2:0] core_csr_new_dcsr_cause = core_csr__new_dcsr_WIRE [8:6]; 
    wire core_csr_new_dcsr_stoptime = core_csr__new_dcsr_WIRE [9]; 
    wire core_csr_new_dcsr_stopcycle = core_csr__new_dcsr_WIRE [10]; 
    wire core_csr_new_dcsr_zero2 = core_csr__new_dcsr_WIRE [11]; 
    wire core_csr_new_dcsr_ebreaku = core_csr__new_dcsr_WIRE [12]; 
    wire core_csr_new_dcsr_ebreaks = core_csr__new_dcsr_WIRE [13]; 
    wire core_csr_new_dcsr_ebreakh = core_csr__new_dcsr_WIRE [14]; 
    wire core_csr_new_dcsr_ebreakm = core_csr__new_dcsr_WIRE [15]; 
    wire[11:0] core_csr_new_dcsr_zero3 = core_csr__new_dcsr_WIRE [27:16]; 
    wire[1:0] core_csr_new_dcsr_zero4 = core_csr__new_dcsr_WIRE [29:28]; 
    wire[1:0] core_csr_new_dcsr_xdebugver = core_csr__new_dcsr_WIRE [31:30]; 
    wire[63:0] core_csr__GEN_81 =~(~ core_csr_wdata |64'h1); 
    wire core_csr__GEN_82 =1'h0== core_csr_reg_tselect &( core_csr_reg_bp_0_control_dmode ==1'h0| core_csr_reg_debug ); 
    wire core_csr__GEN_83 = core_csr_csr_wen & core_csr__GEN_82 ; 
    wire core_csr__GEN_84 = core_csr__GEN_83 & core_csr_decoded_1 ; 
    wire core_csr__reg_bp_0_control_WIRE_r = core_csr__reg_bp_0_control_WIRE_1 [0]; 
    wire core_csr__reg_bp_0_control_WIRE_w = core_csr__reg_bp_0_control_WIRE_1 [1]; 
    wire core_csr__reg_bp_0_control_WIRE_x = core_csr__reg_bp_0_control_WIRE_1 [2]; 
    wire core_csr__reg_bp_0_control_WIRE_u = core_csr__reg_bp_0_control_WIRE_1 [3]; 
    wire core_csr__reg_bp_0_control_WIRE_s = core_csr__reg_bp_0_control_WIRE_1 [4]; 
    wire core_csr__reg_bp_0_control_WIRE_h = core_csr__reg_bp_0_control_WIRE_1 [5]; 
    wire core_csr__reg_bp_0_control_WIRE_m = core_csr__reg_bp_0_control_WIRE_1 [6]; 
    wire[1:0] core_csr__reg_bp_0_control_WIRE_tmatch = core_csr__reg_bp_0_control_WIRE_1 [8:7]; 
    wire[1:0] core_csr__reg_bp_0_control_WIRE_zero = core_csr__reg_bp_0_control_WIRE_1 [10:9]; 
    wire core_csr__reg_bp_0_control_WIRE_chain = core_csr__reg_bp_0_control_WIRE_1 [11]; 
    wire core_csr__reg_bp_0_control_WIRE_action = core_csr__reg_bp_0_control_WIRE_1 [12]; 
    wire[39:0] core_csr__reg_bp_0_control_WIRE_reserved = core_csr__reg_bp_0_control_WIRE_1 [52:13]; 
    wire[5:0] core_csr__reg_bp_0_control_WIRE_maskmax = core_csr__reg_bp_0_control_WIRE_1 [58:53]; 
    wire core_csr__reg_bp_0_control_WIRE_dmode = core_csr__reg_bp_0_control_WIRE_1 [59]; 
    wire[3:0] core_csr__reg_bp_0_control_WIRE_ttype = core_csr__reg_bp_0_control_WIRE_1 [63:60]; 
    wire[1:0] core_csr_newBPC_lo_lo_hi ={ core_csr_reg_bp_0_control_x , core_csr_reg_bp_0_control_w }; 
    wire[2:0] core_csr_newBPC_lo_lo ={ core_csr_newBPC_lo_lo_hi , core_csr_reg_bp_0_control_r }; 
    wire[1:0] core_csr_newBPC_lo_hi_lo ={ core_csr_reg_bp_0_control_s , core_csr_reg_bp_0_control_u }; 
    wire[1:0] core_csr_newBPC_lo_hi_hi ={ core_csr_reg_bp_0_control_m , core_csr_reg_bp_0_control_h }; 
    wire[3:0] core_csr_newBPC_lo_hi ={ core_csr_newBPC_lo_hi_hi , core_csr_newBPC_lo_hi_lo }; 
    wire[6:0] core_csr_newBPC_lo ={ core_csr_newBPC_lo_hi , core_csr_newBPC_lo_lo }; 
    wire[3:0] core_csr_newBPC_hi_lo_lo ={ core_csr_reg_bp_0_control_zero , core_csr_reg_bp_0_control_tmatch }; 
    wire[1:0] core_csr_newBPC_hi_lo_hi ={ core_csr_reg_bp_0_control_action , core_csr_reg_bp_0_control_chain }; 
    wire[5:0] core_csr_newBPC_hi_lo ={ core_csr_newBPC_hi_lo_hi , core_csr_newBPC_hi_lo_lo }; 
    wire[45:0] core_csr_newBPC_hi_hi_lo ={ core_csr_reg_bp_0_control_maskmax , core_csr_reg_bp_0_control_reserved }; 
    wire[4:0] core_csr_newBPC_hi_hi_hi ={ core_csr_reg_bp_0_control_ttype , core_csr_reg_bp_0_control_dmode }; 
    wire[50:0] core_csr_newBPC_hi_hi ={ core_csr_newBPC_hi_hi_hi , core_csr_newBPC_hi_hi_lo }; 
    wire[56:0] core_csr_newBPC_hi ={ core_csr_newBPC_hi_hi , core_csr_newBPC_hi_lo }; 
    wire[63:0] core_csr__newBPC_WIRE =(( core_csr_io_rw_cmd [1] ? { core_csr_newBPC_hi , core_csr_newBPC_lo }:64'h0)| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :64'h0); 
    wire core_csr_newBPC_r = core_csr__newBPC_WIRE [0]; 
    wire core_csr_newBPC_w = core_csr__newBPC_WIRE [1]; 
    wire core_csr_newBPC_x = core_csr__newBPC_WIRE [2]; 
    wire core_csr_newBPC_u = core_csr__newBPC_WIRE [3]; 
    wire core_csr_newBPC_s = core_csr__newBPC_WIRE [4]; 
    wire core_csr_newBPC_h = core_csr__newBPC_WIRE [5]; 
    wire core_csr_newBPC_m = core_csr__newBPC_WIRE [6]; 
    wire[1:0] core_csr_newBPC_tmatch = core_csr__newBPC_WIRE [8:7]; 
    wire[1:0] core_csr_newBPC_zero = core_csr__newBPC_WIRE [10:9]; 
    wire core_csr_newBPC_chain = core_csr__newBPC_WIRE [11]; 
    wire core_csr_newBPC_action = core_csr__newBPC_WIRE [12]; 
    wire[39:0] core_csr_newBPC_reserved = core_csr__newBPC_WIRE [52:13]; 
    wire[5:0] core_csr_newBPC_maskmax = core_csr__newBPC_WIRE [58:53]; 
    wire core_csr_newBPC_dmode = core_csr__newBPC_WIRE [59]; 
    wire[3:0] core_csr_newBPC_ttype = core_csr__newBPC_WIRE [63:60]; 
    wire core_csr_dMode = core_csr_newBPC_dmode & core_csr_reg_debug ; 
    wire core_csr__GEN_85 = core_csr_dMode | core_csr_newBPC_action >1'h1; 
    wire core_csr__GEN_86 =1'h1== core_csr_reg_tselect &( core_csr_reg_bp_1_control_dmode ==1'h0| core_csr_reg_debug ); 
    wire core_csr__GEN_87 = core_csr_csr_wen & core_csr__GEN_86 ; 
    wire core_csr__GEN_88 = core_csr__GEN_87 & core_csr_decoded_1 ; 
    wire core_csr__reg_bp_1_control_WIRE_r = core_csr__reg_bp_1_control_WIRE_1 [0]; 
    wire core_csr__reg_bp_1_control_WIRE_w = core_csr__reg_bp_1_control_WIRE_1 [1]; 
    wire core_csr__reg_bp_1_control_WIRE_x = core_csr__reg_bp_1_control_WIRE_1 [2]; 
    wire core_csr__reg_bp_1_control_WIRE_u = core_csr__reg_bp_1_control_WIRE_1 [3]; 
    wire core_csr__reg_bp_1_control_WIRE_s = core_csr__reg_bp_1_control_WIRE_1 [4]; 
    wire core_csr__reg_bp_1_control_WIRE_h = core_csr__reg_bp_1_control_WIRE_1 [5]; 
    wire core_csr__reg_bp_1_control_WIRE_m = core_csr__reg_bp_1_control_WIRE_1 [6]; 
    wire[1:0] core_csr__reg_bp_1_control_WIRE_tmatch = core_csr__reg_bp_1_control_WIRE_1 [8:7]; 
    wire[1:0] core_csr__reg_bp_1_control_WIRE_zero = core_csr__reg_bp_1_control_WIRE_1 [10:9]; 
    wire core_csr__reg_bp_1_control_WIRE_chain = core_csr__reg_bp_1_control_WIRE_1 [11]; 
    wire core_csr__reg_bp_1_control_WIRE_action = core_csr__reg_bp_1_control_WIRE_1 [12]; 
    wire[39:0] core_csr__reg_bp_1_control_WIRE_reserved = core_csr__reg_bp_1_control_WIRE_1 [52:13]; 
    wire[5:0] core_csr__reg_bp_1_control_WIRE_maskmax = core_csr__reg_bp_1_control_WIRE_1 [58:53]; 
    wire core_csr__reg_bp_1_control_WIRE_dmode = core_csr__reg_bp_1_control_WIRE_1 [59]; 
    wire[3:0] core_csr__reg_bp_1_control_WIRE_ttype = core_csr__reg_bp_1_control_WIRE_1 [63:60]; 
    wire[1:0] core_csr_newBPC_lo_lo_hi_1 ={ core_csr_reg_bp_1_control_x , core_csr_reg_bp_1_control_w }; 
    wire[2:0] core_csr_newBPC_lo_lo_1 ={ core_csr_newBPC_lo_lo_hi_1 , core_csr_reg_bp_1_control_r }; 
    wire[1:0] core_csr_newBPC_lo_hi_lo_1 ={ core_csr_reg_bp_1_control_s , core_csr_reg_bp_1_control_u }; 
    wire[1:0] core_csr_newBPC_lo_hi_hi_1 ={ core_csr_reg_bp_1_control_m , core_csr_reg_bp_1_control_h }; 
    wire[3:0] core_csr_newBPC_lo_hi_1 ={ core_csr_newBPC_lo_hi_hi_1 , core_csr_newBPC_lo_hi_lo_1 }; 
    wire[6:0] core_csr_newBPC_lo_1 ={ core_csr_newBPC_lo_hi_1 , core_csr_newBPC_lo_lo_1 }; 
    wire[3:0] core_csr_newBPC_hi_lo_lo_1 ={ core_csr_reg_bp_1_control_zero , core_csr_reg_bp_1_control_tmatch }; 
    wire[1:0] core_csr_newBPC_hi_lo_hi_1 ={ core_csr_reg_bp_1_control_action , core_csr_reg_bp_1_control_chain }; 
    wire[5:0] core_csr_newBPC_hi_lo_1 ={ core_csr_newBPC_hi_lo_hi_1 , core_csr_newBPC_hi_lo_lo_1 }; 
    wire[45:0] core_csr_newBPC_hi_hi_lo_1 ={ core_csr_reg_bp_1_control_maskmax , core_csr_reg_bp_1_control_reserved }; 
    wire[4:0] core_csr_newBPC_hi_hi_hi_1 ={ core_csr_reg_bp_1_control_ttype , core_csr_reg_bp_1_control_dmode }; 
    wire[50:0] core_csr_newBPC_hi_hi_1 ={ core_csr_newBPC_hi_hi_hi_1 , core_csr_newBPC_hi_hi_lo_1 }; 
    wire[56:0] core_csr_newBPC_hi_1 ={ core_csr_newBPC_hi_hi_1 , core_csr_newBPC_hi_lo_1 }; 
    wire[63:0] core_csr__newBPC_WIRE_1 =(( core_csr_io_rw_cmd [1] ? { core_csr_newBPC_hi_1 , core_csr_newBPC_lo_1 }:64'h0)| core_csr_io_rw_wdata )&~((&( core_csr_io_rw_cmd [1:0])) ?  core_csr_io_rw_wdata :64'h0); 
    wire core_csr_newBPC_1_r = core_csr__newBPC_WIRE_1 [0]; 
    wire core_csr_newBPC_1_w = core_csr__newBPC_WIRE_1 [1]; 
    wire core_csr_newBPC_1_x = core_csr__newBPC_WIRE_1 [2]; 
    wire core_csr_newBPC_1_u = core_csr__newBPC_WIRE_1 [3]; 
    wire core_csr_newBPC_1_s = core_csr__newBPC_WIRE_1 [4]; 
    wire core_csr_newBPC_1_h = core_csr__newBPC_WIRE_1 [5]; 
    wire core_csr_newBPC_1_m = core_csr__newBPC_WIRE_1 [6]; 
    wire[1:0] core_csr_newBPC_1_tmatch = core_csr__newBPC_WIRE_1 [8:7]; 
    wire[1:0] core_csr_newBPC_1_zero = core_csr__newBPC_WIRE_1 [10:9]; 
    wire core_csr_newBPC_1_chain = core_csr__newBPC_WIRE_1 [11]; 
    wire core_csr_newBPC_1_action = core_csr__newBPC_WIRE_1 [12]; 
    wire[39:0] core_csr_newBPC_1_reserved = core_csr__newBPC_WIRE_1 [52:13]; 
    wire[5:0] core_csr_newBPC_1_maskmax = core_csr__newBPC_WIRE_1 [58:53]; 
    wire core_csr_newBPC_1_dmode = core_csr__newBPC_WIRE_1 [59]; 
    wire[3:0] core_csr_newBPC_1_ttype = core_csr__newBPC_WIRE_1 [63:60]; 
    wire core_csr_dMode_1 = core_csr_newBPC_1_dmode & core_csr_reg_debug &( core_csr_reg_bp_0_control_dmode | core_csr_reg_bp_0_control_chain ==1'h0); 
    wire core_csr__GEN_89 = core_csr_dMode_1 | core_csr_newBPC_1_action >1'h1; 
    wire core_csr__GEN_90 = core_csr_decoded_109 & core_csr_reg_pmp_0_cfg_l ==1'h0; 
    wire[7:0] core_csr__newCfg_WIRE = core_csr_wdata [7:0]; 
    wire core_csr_newCfg_r = core_csr__newCfg_WIRE [0]; 
    wire core_csr_newCfg_w = core_csr__newCfg_WIRE [1]; 
    wire core_csr_newCfg_x = core_csr__newCfg_WIRE [2]; 
    wire[1:0] core_csr_newCfg_a = core_csr__newCfg_WIRE [4:3]; 
    wire[1:0] core_csr_newCfg_res = core_csr__newCfg_WIRE [6:5]; 
    wire core_csr_newCfg_l = core_csr__newCfg_WIRE [7]; 
    wire core_csr__GEN_91 = core_csr_newCfg_w & core_csr_newCfg_r ; 
    wire core_csr__GEN_92 = core_csr_decoded_111 &( core_csr_reg_pmp_0_cfg_l | core_csr_reg_pmp_1_cfg_l & core_csr_reg_pmp_1_cfg_a [1]==1'h0& core_csr_reg_pmp_1_cfg_a [0])==1'h0; 
    wire core_csr__GEN_93 = core_csr_decoded_109 & core_csr_reg_pmp_1_cfg_l ==1'h0; 
    wire[55:0] core_csr__wdata_63to8 = core_csr_wdata [63:8]; 
    wire[7:0] core_csr__newCfg_WIRE_1 = core_csr__wdata_63to8 [7:0]; 
    wire core_csr_newCfg_1_r = core_csr__newCfg_WIRE_1 [0]; 
    wire core_csr_newCfg_1_w = core_csr__newCfg_WIRE_1 [1]; 
    wire core_csr_newCfg_1_x = core_csr__newCfg_WIRE_1 [2]; 
    wire[1:0] core_csr_newCfg_1_a = core_csr__newCfg_WIRE_1 [4:3]; 
    wire[1:0] core_csr_newCfg_1_res = core_csr__newCfg_WIRE_1 [6:5]; 
    wire core_csr_newCfg_1_l = core_csr__newCfg_WIRE_1 [7]; 
    wire core_csr__GEN_94 = core_csr_newCfg_1_w & core_csr_newCfg_1_r ; 
    wire core_csr__GEN_95 = core_csr_decoded_112 &( core_csr_reg_pmp_1_cfg_l | core_csr_reg_pmp_2_cfg_l & core_csr_reg_pmp_2_cfg_a [1]==1'h0& core_csr_reg_pmp_2_cfg_a [0])==1'h0; 
    wire core_csr__GEN_96 = core_csr_decoded_109 & core_csr_reg_pmp_2_cfg_l ==1'h0; 
    wire[47:0] core_csr__wdata_63to16 = core_csr_wdata [63:16]; 
    wire[7:0] core_csr__newCfg_WIRE_2 = core_csr__wdata_63to16 [7:0]; 
    wire core_csr_newCfg_2_r = core_csr__newCfg_WIRE_2 [0]; 
    wire core_csr_newCfg_2_w = core_csr__newCfg_WIRE_2 [1]; 
    wire core_csr_newCfg_2_x = core_csr__newCfg_WIRE_2 [2]; 
    wire[1:0] core_csr_newCfg_2_a = core_csr__newCfg_WIRE_2 [4:3]; 
    wire[1:0] core_csr_newCfg_2_res = core_csr__newCfg_WIRE_2 [6:5]; 
    wire core_csr_newCfg_2_l = core_csr__newCfg_WIRE_2 [7]; 
    wire core_csr__GEN_97 = core_csr_newCfg_2_w & core_csr_newCfg_2_r ; 
    wire core_csr__GEN_98 = core_csr_decoded_113 &( core_csr_reg_pmp_2_cfg_l | core_csr_reg_pmp_3_cfg_l & core_csr_reg_pmp_3_cfg_a [1]==1'h0& core_csr_reg_pmp_3_cfg_a [0])==1'h0; 
    wire core_csr__GEN_99 = core_csr_decoded_109 & core_csr_reg_pmp_3_cfg_l ==1'h0; 
    wire[39:0] core_csr__wdata_63to24 = core_csr_wdata [63:24]; 
    wire[7:0] core_csr__newCfg_WIRE_3 = core_csr__wdata_63to24 [7:0]; 
    wire core_csr_newCfg_3_r = core_csr__newCfg_WIRE_3 [0]; 
    wire core_csr_newCfg_3_w = core_csr__newCfg_WIRE_3 [1]; 
    wire core_csr_newCfg_3_x = core_csr__newCfg_WIRE_3 [2]; 
    wire[1:0] core_csr_newCfg_3_a = core_csr__newCfg_WIRE_3 [4:3]; 
    wire[1:0] core_csr_newCfg_3_res = core_csr__newCfg_WIRE_3 [6:5]; 
    wire core_csr_newCfg_3_l = core_csr__newCfg_WIRE_3 [7]; 
    wire core_csr__GEN_100 = core_csr_newCfg_3_w & core_csr_newCfg_3_r ; 
    wire core_csr__GEN_101 = core_csr_decoded_114 &( core_csr_reg_pmp_3_cfg_l | core_csr_reg_pmp_4_cfg_l & core_csr_reg_pmp_4_cfg_a [1]==1'h0& core_csr_reg_pmp_4_cfg_a [0])==1'h0; 
    wire core_csr__GEN_102 = core_csr_decoded_109 & core_csr_reg_pmp_4_cfg_l ==1'h0; 
    wire[31:0] core_csr__wdata_63to32 = core_csr_wdata [63:32]; 
    wire[7:0] core_csr__newCfg_WIRE_4 = core_csr__wdata_63to32 [7:0]; 
    wire core_csr_newCfg_4_r = core_csr__newCfg_WIRE_4 [0]; 
    wire core_csr_newCfg_4_w = core_csr__newCfg_WIRE_4 [1]; 
    wire core_csr_newCfg_4_x = core_csr__newCfg_WIRE_4 [2]; 
    wire[1:0] core_csr_newCfg_4_a = core_csr__newCfg_WIRE_4 [4:3]; 
    wire[1:0] core_csr_newCfg_4_res = core_csr__newCfg_WIRE_4 [6:5]; 
    wire core_csr_newCfg_4_l = core_csr__newCfg_WIRE_4 [7]; 
    wire core_csr__GEN_103 = core_csr_newCfg_4_w & core_csr_newCfg_4_r ; 
    wire core_csr__GEN_104 = core_csr_decoded_115 &( core_csr_reg_pmp_4_cfg_l | core_csr_reg_pmp_5_cfg_l & core_csr_reg_pmp_5_cfg_a [1]==1'h0& core_csr_reg_pmp_5_cfg_a [0])==1'h0; 
    wire core_csr__GEN_105 = core_csr_decoded_109 & core_csr_reg_pmp_5_cfg_l ==1'h0; 
    wire[23:0] core_csr__wdata_63to40 = core_csr_wdata [63:40]; 
    wire[7:0] core_csr__newCfg_WIRE_5 = core_csr__wdata_63to40 [7:0]; 
    wire core_csr_newCfg_5_r = core_csr__newCfg_WIRE_5 [0]; 
    wire core_csr_newCfg_5_w = core_csr__newCfg_WIRE_5 [1]; 
    wire core_csr_newCfg_5_x = core_csr__newCfg_WIRE_5 [2]; 
    wire[1:0] core_csr_newCfg_5_a = core_csr__newCfg_WIRE_5 [4:3]; 
    wire[1:0] core_csr_newCfg_5_res = core_csr__newCfg_WIRE_5 [6:5]; 
    wire core_csr_newCfg_5_l = core_csr__newCfg_WIRE_5 [7]; 
    wire core_csr__GEN_106 = core_csr_newCfg_5_w & core_csr_newCfg_5_r ; 
    wire core_csr__GEN_107 = core_csr_decoded_116 &( core_csr_reg_pmp_5_cfg_l | core_csr_reg_pmp_6_cfg_l & core_csr_reg_pmp_6_cfg_a [1]==1'h0& core_csr_reg_pmp_6_cfg_a [0])==1'h0; 
    wire core_csr__GEN_108 = core_csr_decoded_109 & core_csr_reg_pmp_6_cfg_l ==1'h0; 
    wire[15:0] core_csr__wdata_63to48 = core_csr_wdata [63:48]; 
    wire[7:0] core_csr__newCfg_WIRE_6 = core_csr__wdata_63to48 [7:0]; 
    wire core_csr_newCfg_6_r = core_csr__newCfg_WIRE_6 [0]; 
    wire core_csr_newCfg_6_w = core_csr__newCfg_WIRE_6 [1]; 
    wire core_csr_newCfg_6_x = core_csr__newCfg_WIRE_6 [2]; 
    wire[1:0] core_csr_newCfg_6_a = core_csr__newCfg_WIRE_6 [4:3]; 
    wire[1:0] core_csr_newCfg_6_res = core_csr__newCfg_WIRE_6 [6:5]; 
    wire core_csr_newCfg_6_l = core_csr__newCfg_WIRE_6 [7]; 
    wire core_csr__GEN_109 = core_csr_newCfg_6_w & core_csr_newCfg_6_r ; 
    wire core_csr__GEN_110 = core_csr_decoded_117 &( core_csr_reg_pmp_6_cfg_l | core_csr_reg_pmp_7_cfg_l & core_csr_reg_pmp_7_cfg_a [1]==1'h0& core_csr_reg_pmp_7_cfg_a [0])==1'h0; 
    wire core_csr__GEN_111 = core_csr_decoded_109 & core_csr_reg_pmp_7_cfg_l ==1'h0; 
    wire[7:0] core_csr__newCfg_WIRE_7 = core_csr_wdata [63:56]; 
    wire core_csr_newCfg_7_r = core_csr__newCfg_WIRE_7 [0]; 
    wire core_csr_newCfg_7_w = core_csr__newCfg_WIRE_7 [1]; 
    wire core_csr_newCfg_7_x = core_csr__newCfg_WIRE_7 [2]; 
    wire[1:0] core_csr_newCfg_7_a = core_csr__newCfg_WIRE_7 [4:3]; 
    wire[1:0] core_csr_newCfg_7_res = core_csr__newCfg_WIRE_7 [6:5]; 
    wire core_csr_newCfg_7_l = core_csr__newCfg_WIRE_7 [7]; 
    wire core_csr__GEN_112 = core_csr_newCfg_7_w & core_csr_newCfg_7_r ; 
    wire core_csr__GEN_113 = core_csr_decoded_118 &( core_csr_reg_pmp_7_cfg_l | core_csr_reg_pmp_7_cfg_l & core_csr_reg_pmp_7_cfg_a [1]==1'h0& core_csr_reg_pmp_7_cfg_a [0])==1'h0; 
    wire[63:0] core_csr__GEN_114 = core_csr_wdata &64'h208| core_csr_reg_custom_0 &64'hFFFFFFFFFFFFFDF7; 
    wire[63:0] core_csr__GEN_115 = core_csr_reg_custom_1 |64'h0; 
    wire[63:0] core_csr__GEN_116 = core_csr_reg_custom_2 |64'h0; 
    wire[63:0] core_csr__GEN_117 = core_csr_reg_custom_3 |64'h0; 
    wire[63:0] core_csr__GEN_118 = core_csr_io_customCSRs_0_sdata &64'h208| core_csr_reg_custom_0 &64'hFFFFFFFFFFFFFDF7; 
    wire[63:0] core_csr__GEN_119 = core_csr_reg_custom_1 |64'h0; 
    wire[63:0] core_csr__GEN_120 = core_csr_reg_custom_2 |64'h0; 
    wire[63:0] core_csr__GEN_121 = core_csr_reg_custom_3 |64'h0; 
    wire core_csr__io_trace_0_exception_output = core_csr_io_retire >=1'h0& core_csr_exception ; 
  always @( posedge  core_csr_clock )
         begin 
             if ( core_csr_reset )
                 begin  
                     core_csr_reg_mstatus_debug  <= core_csr_reset_mstatus_debug ; 
                     core_csr_reg_mstatus_cease  <= core_csr_reset_mstatus_cease ; 
                     core_csr_reg_mstatus_wfi  <= core_csr_reset_mstatus_wfi ; 
                     core_csr_reg_mstatus_isa  <= core_csr_reset_mstatus_isa ; 
                     core_csr_reg_mstatus_dprv  <= core_csr_reset_mstatus_dprv ; 
                     core_csr_reg_mstatus_dv  <= core_csr_reset_mstatus_dv ; 
                     core_csr_reg_mstatus_prv  <= core_csr_reset_mstatus_prv ; 
                     core_csr_reg_mstatus_v  <= core_csr_reset_mstatus_v ; 
                     core_csr_reg_mstatus_sd  <= core_csr_reset_mstatus_sd ; 
                     core_csr_reg_mstatus_zero2  <= core_csr_reset_mstatus_zero2 ; 
                     core_csr_reg_mstatus_mpv  <= core_csr_reset_mstatus_mpv ; 
                     core_csr_reg_mstatus_gva  <= core_csr_reset_mstatus_gva ; 
                     core_csr_reg_mstatus_mbe  <= core_csr_reset_mstatus_mbe ; 
                     core_csr_reg_mstatus_sbe  <= core_csr_reset_mstatus_sbe ; 
                     core_csr_reg_mstatus_sxl  <= core_csr_reset_mstatus_sxl ; 
                     core_csr_reg_mstatus_uxl  <= core_csr_reset_mstatus_uxl ; 
                     core_csr_reg_mstatus_sd_rv32  <= core_csr_reset_mstatus_sd_rv32 ; 
                     core_csr_reg_mstatus_zero1  <= core_csr_reset_mstatus_zero1 ; 
                     core_csr_reg_mstatus_tsr  <= core_csr_reset_mstatus_tsr ; 
                     core_csr_reg_mstatus_tw  <= core_csr_reset_mstatus_tw ; 
                     core_csr_reg_mstatus_tvm  <= core_csr_reset_mstatus_tvm ; 
                     core_csr_reg_mstatus_mxr  <= core_csr_reset_mstatus_mxr ; 
                     core_csr_reg_mstatus_sum  <= core_csr_reset_mstatus_sum ; 
                     core_csr_reg_mstatus_mprv  <= core_csr_reset_mstatus_mprv ; 
                     core_csr_reg_mstatus_xs  <= core_csr_reset_mstatus_xs ; 
                     core_csr_reg_mstatus_fs  <= core_csr_reset_mstatus_fs ; 
                     core_csr_reg_mstatus_mpp  <= core_csr_reset_mstatus_mpp ; 
                     core_csr_reg_mstatus_vs  <= core_csr_reset_mstatus_vs ; 
                     core_csr_reg_mstatus_spp  <= core_csr_reset_mstatus_spp ; 
                     core_csr_reg_mstatus_mpie  <= core_csr_reset_mstatus_mpie ; 
                     core_csr_reg_mstatus_ube  <= core_csr_reset_mstatus_ube ; 
                     core_csr_reg_mstatus_spie  <= core_csr_reset_mstatus_spie ; 
                     core_csr_reg_mstatus_upie  <= core_csr_reset_mstatus_upie ; 
                     core_csr_reg_mstatus_mie  <= core_csr_reset_mstatus_mie ; 
                     core_csr_reg_mstatus_hie  <= core_csr_reset_mstatus_hie ; 
                     core_csr_reg_mstatus_sie  <= core_csr_reset_mstatus_sie ; 
                     core_csr_reg_mstatus_uie  <= core_csr_reset_mstatus_uie ; 
                     core_csr_reg_dcsr_xdebugver  <= core_csr_reset_dcsr_xdebugver ; 
                     core_csr_reg_dcsr_zero4  <= core_csr_reset_dcsr_zero4 ; 
                     core_csr_reg_dcsr_zero3  <= core_csr_reset_dcsr_zero3 ; 
                     core_csr_reg_dcsr_ebreakm  <= core_csr_reset_dcsr_ebreakm ; 
                     core_csr_reg_dcsr_ebreakh  <= core_csr_reset_dcsr_ebreakh ; 
                     core_csr_reg_dcsr_ebreaks  <= core_csr_reset_dcsr_ebreaks ; 
                     core_csr_reg_dcsr_ebreaku  <= core_csr_reset_dcsr_ebreaku ; 
                     core_csr_reg_dcsr_zero2  <= core_csr_reset_dcsr_zero2 ; 
                     core_csr_reg_dcsr_stopcycle  <= core_csr_reset_dcsr_stopcycle ; 
                     core_csr_reg_dcsr_stoptime  <= core_csr_reset_dcsr_stoptime ; 
                     core_csr_reg_dcsr_cause  <= core_csr_reset_dcsr_cause ; 
                     core_csr_reg_dcsr_v  <= core_csr_reset_dcsr_v ; 
                     core_csr_reg_dcsr_zero1  <= core_csr_reset_dcsr_zero1 ; 
                     core_csr_reg_dcsr_step  <= core_csr_reset_dcsr_step ; 
                     core_csr_reg_dcsr_prv  <= core_csr_reset_dcsr_prv ; 
                     core_csr_reg_debug  <=1'h0; 
                     core_csr_reg_mcause  <=64'h0; 
                     core_csr_reg_mtvec  <=32'h0; 
                     core_csr_reg_mncause  <=64'h0; 
                     core_csr_reg_mnstatus_mpp  <= core_csr_reset_mnstatus_mpp ; 
                     core_csr_reg_mnstatus_zero3  <= core_csr_reset_mnstatus_zero3 ; 
                     core_csr_reg_mnstatus_mpv  <= core_csr_reset_mnstatus_mpv ; 
                     core_csr_reg_mnstatus_zero2  <= core_csr_reset_mnstatus_zero2 ; 
                     core_csr_reg_mnstatus_mie  <= core_csr_reset_mnstatus_mie ; 
                     core_csr_reg_mnstatus_zero1  <= core_csr_reset_mnstatus_zero1 ; 
                     core_csr_reg_rnmie  <=1'h1; 
                     core_csr_reg_menvcfg_stce  <= core_csr__reg_menvcfg_WIRE_stce ; 
                     core_csr_reg_menvcfg_pbmte  <= core_csr__reg_menvcfg_WIRE_pbmte ; 
                     core_csr_reg_menvcfg_zero54  <= core_csr__reg_menvcfg_WIRE_zero54 ; 
                     core_csr_reg_menvcfg_cbze  <= core_csr__reg_menvcfg_WIRE_cbze ; 
                     core_csr_reg_menvcfg_cbcfe  <= core_csr__reg_menvcfg_WIRE_cbcfe ; 
                     core_csr_reg_menvcfg_cbie  <= core_csr__reg_menvcfg_WIRE_cbie ; 
                     core_csr_reg_menvcfg_zero3  <= core_csr__reg_menvcfg_WIRE_zero3 ; 
                     core_csr_reg_menvcfg_fiom  <= core_csr__reg_menvcfg_WIRE_fiom ; 
                     core_csr_reg_senvcfg_stce  <= core_csr__reg_senvcfg_WIRE_stce ; 
                     core_csr_reg_senvcfg_pbmte  <= core_csr__reg_senvcfg_WIRE_pbmte ; 
                     core_csr_reg_senvcfg_zero54  <= core_csr__reg_senvcfg_WIRE_zero54 ; 
                     core_csr_reg_senvcfg_cbze  <= core_csr__reg_senvcfg_WIRE_cbze ; 
                     core_csr_reg_senvcfg_cbcfe  <= core_csr__reg_senvcfg_WIRE_cbcfe ; 
                     core_csr_reg_senvcfg_cbie  <= core_csr__reg_senvcfg_WIRE_cbie ; 
                     core_csr_reg_senvcfg_zero3  <= core_csr__reg_senvcfg_WIRE_zero3 ; 
                     core_csr_reg_senvcfg_fiom  <= core_csr__reg_senvcfg_WIRE_fiom ; 
                     core_csr_reg_henvcfg_stce  <= core_csr__reg_henvcfg_WIRE_stce ; 
                     core_csr_reg_henvcfg_pbmte  <= core_csr__reg_henvcfg_WIRE_pbmte ; 
                     core_csr_reg_henvcfg_zero54  <= core_csr__reg_henvcfg_WIRE_zero54 ; 
                     core_csr_reg_henvcfg_cbze  <= core_csr__reg_henvcfg_WIRE_cbze ; 
                     core_csr_reg_henvcfg_cbcfe  <= core_csr__reg_henvcfg_WIRE_cbcfe ; 
                     core_csr_reg_henvcfg_cbie  <= core_csr__reg_henvcfg_WIRE_cbie ; 
                     core_csr_reg_henvcfg_zero3  <= core_csr__reg_henvcfg_WIRE_zero3 ; 
                     core_csr_reg_henvcfg_fiom  <= core_csr__reg_henvcfg_WIRE_fiom ; 
                     core_csr_reg_hstatus_zero6  <= core_csr__reg_hstatus_WIRE_zero6 ; 
                     core_csr_reg_hstatus_vsxl  <= core_csr__reg_hstatus_WIRE_vsxl ; 
                     core_csr_reg_hstatus_zero5  <= core_csr__reg_hstatus_WIRE_zero5 ; 
                     core_csr_reg_hstatus_vtsr  <= core_csr__reg_hstatus_WIRE_vtsr ; 
                     core_csr_reg_hstatus_vtw  <= core_csr__reg_hstatus_WIRE_vtw ; 
                     core_csr_reg_hstatus_vtvm  <= core_csr__reg_hstatus_WIRE_vtvm ; 
                     core_csr_reg_hstatus_zero3  <= core_csr__reg_hstatus_WIRE_zero3 ; 
                     core_csr_reg_hstatus_vgein  <= core_csr__reg_hstatus_WIRE_vgein ; 
                     core_csr_reg_hstatus_zero2  <= core_csr__reg_hstatus_WIRE_zero2 ; 
                     core_csr_reg_hstatus_hu  <= core_csr__reg_hstatus_WIRE_hu ; 
                     core_csr_reg_hstatus_spvp  <= core_csr__reg_hstatus_WIRE_spvp ; 
                     core_csr_reg_hstatus_spv  <= core_csr__reg_hstatus_WIRE_spv ; 
                     core_csr_reg_hstatus_gva  <= core_csr__reg_hstatus_WIRE_gva ; 
                     core_csr_reg_hstatus_vsbe  <= core_csr__reg_hstatus_WIRE_vsbe ; 
                     core_csr_reg_hstatus_zero1  <= core_csr__reg_hstatus_WIRE_zero1 ; 
                     core_csr_reg_mcountinhibit  <=3'h0; 
                     core_csr_small_0  <=6'h0; 
                     core_csr_large_0  <=58'h0; 
                     core_csr_reg_misa  <=64'h8000000000801105; 
                     core_csr_reg_custom_0  <=64'h208; 
                     core_csr_reg_custom_1  <=64'h1; 
                     core_csr_reg_custom_2  <=64'h0; 
                     core_csr_reg_custom_3  <=64'h20181004; 
                     core_csr_io_status_cease_r  <=1'h0;
                 end 
              else 
                 begin  
                     core_csr_reg_mstatus_prv  <=2'h3;
                     if ( core_csr_insn_ret )
                         begin  
                             core_csr_reg_mstatus_v  <=1'h0;
                             if ( core_csr__GEN_70 )
                                 begin 
                                     if ( core_csr_exception )
                                         begin 
                                             if ( core_csr_trapToDebug )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr_trapToNmiInt )
                                                     begin 
                                                     end 
                                                  else 
                                                     if ( core_csr__GEN_58 )
                                                         begin 
                                                         end 
                                                      else 
                                                         if ( core_csr__GEN_61 )
                                                             begin 
                                                             end 
                                                          else 
                                                             begin  
                                                                 core_csr_reg_mstatus_mpv  <= core_csr_reg_mstatus_v ; 
                                                                 core_csr_reg_mstatus_mpp  <=2'h3;
                                                             end 
                                         end 
                                      else 
                                         begin 
                                         end  
                                     core_csr_reg_debug  <=1'h0;
                                 end 
                              else 
                                 begin  
                                     core_csr_reg_mstatus_mpv  <=1'h0; 
                                     core_csr_reg_mstatus_mpp  <=2'h3;
                                     if ( core_csr_exception )
                                         begin 
                                             if ( core_csr_trapToDebug )
                                                 begin 
                                                     if ( core_csr__GEN_51 ) 
                                                         core_csr_reg_debug  <=1'h1;
                                                      else 
                                                         begin 
                                                         end 
                                                 end 
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else 
                                         begin 
                                         end 
                                 end 
                         end 
                      else 
                         if ( core_csr_exception )
                             begin 
                                 if ( core_csr_trapToDebug )
                                     begin 
                                         if ( core_csr__GEN_51 )
                                             begin  
                                                 core_csr_reg_mstatus_v  <=1'h0; 
                                                 core_csr_reg_debug  <=1'h1;
                                             end 
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     if ( core_csr_trapToNmiInt )
                                         begin 
                                             if ( core_csr_reg_rnmie ) 
                                                 core_csr_reg_mstatus_v  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else 
                                         begin  
                                             core_csr_reg_mstatus_v  <= core_csr__GEN_58 ;
                                             if ( core_csr__GEN_58 )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr__GEN_61 )
                                                     begin 
                                                     end 
                                                  else 
                                                     begin  
                                                         core_csr_reg_mstatus_mpv  <= core_csr_reg_mstatus_v ; 
                                                         core_csr_reg_mstatus_mpp  <=2'h3;
                                                     end 
                                         end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_exception )
                         begin 
                             if ( core_csr_trapToDebug )
                                 begin 
                                     if ( core_csr__GEN_51 )
                                         begin  
                                             core_csr_reg_dcsr_cause  <= core_csr__GEN_54 ; 
                                             core_csr_reg_dcsr_v  <= core_csr_reg_mstatus_v ; 
                                             core_csr_reg_dcsr_prv  <=2'h3;
                                         end 
                                      else 
                                         begin 
                                         end 
                                 end 
                              else 
                                 if ( core_csr_trapToNmiInt )
                                     begin 
                                         if ( core_csr_reg_rnmie )
                                             begin  
                                                 core_csr_reg_mncause  <= core_csr__GEN_56 ; 
                                                 core_csr_reg_mnstatus_mpp  <=2'h3; 
                                                 core_csr_reg_mnstatus_mpv  <= core_csr_reg_mstatus_v ; 
                                                 core_csr_reg_rnmie  <=1'h0;
                                             end 
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     if ( core_csr__GEN_58 )
                                         begin 
                                         end 
                                      else 
                                         if ( core_csr__GEN_61 )
                                             begin  
                                                 core_csr_reg_mstatus_spp  <= core_csr_reg_mstatus_prv [0]; 
                                                 core_csr_reg_mstatus_spie  <= core_csr_reg_mstatus_sie ; 
                                                 core_csr_reg_mstatus_sie  <=1'h0;
                                                 if ( core_csr_reg_mstatus_v ) 
                                                     core_csr_reg_hstatus_spvp  <= core_csr_reg_mstatus_prv [0];
                                                  else 
                                                     begin 
                                                     end  
                                                 core_csr_reg_hstatus_spv  <= core_csr_reg_mstatus_v ; 
                                                 core_csr_reg_hstatus_gva  <= core_csr_io_gva ;
                                             end 
                                          else  
                                             core_csr_reg_mstatus_gva  <= core_csr_io_gva ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr_csr_wen )
                         begin 
                             if ( core_csr_decoded_5 )
                                 begin  
                                     core_csr_reg_mstatus_vs  <=2'h0; 
                                     core_csr_reg_mstatus_mpie  <= core_csr_new_mstatus_mpie ; 
                                     core_csr_reg_mstatus_mie  <= core_csr_new_mstatus_mie ;
                                 end 
                              else 
                                 if ( core_csr_insn_ret )
                                     begin 
                                         if ( core_csr__GEN_70 )
                                             begin 
                                                 if ( core_csr_exception )
                                                     begin 
                                                         if ( core_csr_trapToDebug )
                                                             begin 
                                                             end 
                                                          else 
                                                             if ( core_csr_trapToNmiInt )
                                                                 begin 
                                                                 end 
                                                              else 
                                                                 if ( core_csr__GEN_58 )
                                                                     begin 
                                                                     end 
                                                                  else 
                                                                     if ( core_csr__GEN_61 )
                                                                         begin 
                                                                         end 
                                                                      else 
                                                                         begin  
                                                                             core_csr_reg_mstatus_mpie  <= core_csr_reg_mstatus_mie ; 
                                                                             core_csr_reg_mstatus_mie  <=1'h0;
                                                                         end 
                                                     end 
                                                  else 
                                                     begin 
                                                     end 
                                             end 
                                          else 
                                             begin  
                                                 core_csr_reg_mstatus_mpie  <=1'h1; 
                                                 core_csr_reg_mstatus_mie  <= core_csr_reg_mstatus_mpie ;
                                             end 
                                     end 
                                  else 
                                     if ( core_csr_exception )
                                         begin 
                                             if ( core_csr_trapToDebug )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr_trapToNmiInt )
                                                     begin 
                                                     end 
                                                  else 
                                                     if ( core_csr__GEN_58 )
                                                         begin 
                                                         end 
                                                      else 
                                                         if ( core_csr__GEN_61 )
                                                             begin 
                                                             end 
                                                          else 
                                                             begin  
                                                                 core_csr_reg_mstatus_mpie  <= core_csr_reg_mstatus_mie ; 
                                                                 core_csr_reg_mstatus_mie  <=1'h0;
                                                             end 
                                         end 
                                      else 
                                         begin 
                                         end 
                             if ( core_csr_decoded_14 )
                                 begin  
                                     core_csr_reg_dcsr_ebreakm  <= core_csr_new_dcsr_ebreakm ; 
                                     core_csr_reg_dcsr_step  <= core_csr_new_dcsr_step ;
                                 end 
                              else 
                                 begin 
                                 end 
                             if ( core_csr_decoded_12 ) 
                                 core_csr_reg_mcause  <= core_csr__GEN_79 ;
                              else 
                                 if ( core_csr_exception )
                                     begin 
                                         if ( core_csr_trapToDebug )
                                             begin 
                                             end 
                                          else 
                                             if ( core_csr_trapToNmiInt )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr__GEN_58 )
                                                     begin 
                                                     end 
                                                  else 
                                                     if ( core_csr__GEN_61 )
                                                         begin 
                                                         end 
                                                      else  
                                                         core_csr_reg_mcause  <= core_csr_cause ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             if ( core_csr_decoded_6 ) 
                                 core_csr_reg_mtvec  <= core_csr_wdata [31:0];
                              else 
                                 begin 
                                 end 
                             if ( core_csr_decoded_17 ) 
                                 core_csr_reg_mcountinhibit  <= core_csr__GEN_80 [2:0];
                              else 
                                 begin 
                                 end 
                             if ( core_csr_decoded_19 )
                                 begin  
                                     core_csr_small_0  <= core_csr_wdata [5:0]; 
                                     core_csr_large_0  <= core_csr_wdata [63:6];
                                 end 
                              else 
                                 begin 
                                     if ( core_csr__GEN_0 ) 
                                         core_csr_small_0  <= core_csr_nextSmall [5:0];
                                      else 
                                         begin 
                                         end 
                                     if ( core_csr__GEN_2 ) 
                                         core_csr_large_0  <= core_csr__GEN_3 [57:0];
                                      else 
                                         begin 
                                         end 
                                 end 
                             if ( core_csr_decoded_4 )
                                 begin 
                                     if ( core_csr__GEN_74 ) 
                                         core_csr_reg_misa  <= core_csr__GEN_75 ;
                                      else 
                                         begin 
                                         end 
                                 end 
                              else 
                                 begin 
                                 end 
                         end 
                      else 
                         begin 
                             if ( core_csr_insn_ret )
                                 begin 
                                     if ( core_csr__GEN_70 )
                                         begin 
                                             if ( core_csr_exception )
                                                 begin 
                                                     if ( core_csr_trapToDebug )
                                                         begin 
                                                         end 
                                                      else 
                                                         if ( core_csr_trapToNmiInt )
                                                             begin 
                                                             end 
                                                          else 
                                                             if ( core_csr__GEN_58 )
                                                                 begin 
                                                                 end 
                                                              else 
                                                                 if ( core_csr__GEN_61 )
                                                                     begin 
                                                                     end 
                                                                  else 
                                                                     begin  
                                                                         core_csr_reg_mstatus_mpie  <= core_csr_reg_mstatus_mie ; 
                                                                         core_csr_reg_mstatus_mie  <=1'h0;
                                                                     end 
                                                 end 
                                              else 
                                                 begin 
                                                 end 
                                         end 
                                      else 
                                         begin  
                                             core_csr_reg_mstatus_mpie  <=1'h1; 
                                             core_csr_reg_mstatus_mie  <= core_csr_reg_mstatus_mpie ;
                                         end 
                                 end 
                              else 
                                 if ( core_csr_exception )
                                     begin 
                                         if ( core_csr_trapToDebug )
                                             begin 
                                             end 
                                          else 
                                             if ( core_csr_trapToNmiInt )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr__GEN_58 )
                                                     begin 
                                                     end 
                                                  else 
                                                     if ( core_csr__GEN_61 )
                                                         begin 
                                                         end 
                                                      else 
                                                         begin  
                                                             core_csr_reg_mstatus_mpie  <= core_csr_reg_mstatus_mie ; 
                                                             core_csr_reg_mstatus_mie  <=1'h0;
                                                         end 
                                     end 
                                  else 
                                     begin 
                                     end 
                             if ( core_csr_exception )
                                 begin 
                                     if ( core_csr_trapToDebug )
                                         begin 
                                         end 
                                      else 
                                         if ( core_csr_trapToNmiInt )
                                             begin 
                                             end 
                                          else 
                                             if ( core_csr__GEN_58 )
                                                 begin 
                                                 end 
                                              else 
                                                 if ( core_csr__GEN_61 )
                                                     begin 
                                                     end 
                                                  else  
                                                     core_csr_reg_mcause  <= core_csr_cause ;
                                 end 
                              else 
                                 begin 
                                 end 
                             if ( core_csr__GEN_0 ) 
                                 core_csr_small_0  <= core_csr_nextSmall [5:0];
                              else 
                                 begin 
                                 end 
                             if ( core_csr__GEN_2 ) 
                                 core_csr_large_0  <= core_csr__GEN_3 [57:0];
                              else 
                                 begin 
                                 end 
                         end 
                     if ( core_csr_io_customCSRs_0_set ) 
                         core_csr_reg_custom_0  <= core_csr__GEN_118 ;
                      else 
                         if ( core_csr_csr_wen )
                             begin 
                                 if ( core_csr_decoded_127 ) 
                                     core_csr_reg_custom_0  <= core_csr__GEN_114 ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_io_customCSRs_1_set ) 
                         core_csr_reg_custom_1  <= core_csr__GEN_119 ;
                      else 
                         if ( core_csr_csr_wen )
                             begin 
                                 if ( core_csr_decoded_128 ) 
                                     core_csr_reg_custom_1  <= core_csr__GEN_115 ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_io_customCSRs_2_set ) 
                         core_csr_reg_custom_2  <= core_csr__GEN_120 ;
                      else 
                         if ( core_csr_csr_wen )
                             begin 
                                 if ( core_csr_decoded_129 ) 
                                     core_csr_reg_custom_2  <= core_csr__GEN_116 ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_io_customCSRs_3_set ) 
                         core_csr_reg_custom_3  <= core_csr__GEN_121 ;
                      else 
                         if ( core_csr_csr_wen )
                             begin 
                                 if ( core_csr_decoded_130 ) 
                                     core_csr_reg_custom_3  <= core_csr__GEN_117 ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_insn_cease ) 
                         core_csr_io_status_cease_r  <=1'h1;
                      else 
                         begin 
                         end 
                 end 
         end
  always @( posedge  core_csr_clock )
         begin 
             if ( core_csr_csr_wen )
                 begin 
                     if ( core_csr_decoded_15 ) 
                         core_csr_reg_dpc  <= core_csr__GEN_81 [33:0];
                      else 
                         if ( core_csr_exception )
                             begin 
                                 if ( core_csr_trapToDebug )
                                     begin 
                                         if ( core_csr__GEN_51 ) 
                                             core_csr_reg_dpc  <= core_csr_epc ;
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_decoded_16 ) 
                         core_csr_reg_dscratch0  <= core_csr_wdata ;
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_82 )
                         begin 
                             if ( core_csr_decoded_1 ) 
                                 core_csr_reg_bp_0_control_tmatch  <= core_csr__reg_bp_0_control_WIRE_tmatch ;
                              else 
                                 begin 
                                 end 
                             if ( core_csr_decoded_2 ) 
                                 core_csr_reg_bp_0_address  <= core_csr_wdata [32:0];
                              else 
                                 begin 
                                 end 
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_90 )
                         begin  
                             core_csr_reg_pmp_0_cfg_x  <= core_csr_newCfg_x ; 
                             core_csr_reg_pmp_0_cfg_w  <= core_csr__GEN_91 ; 
                             core_csr_reg_pmp_0_cfg_r  <= core_csr_newCfg_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_92 ) 
                         core_csr_reg_pmp_0_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_93 )
                         begin  
                             core_csr_reg_pmp_1_cfg_x  <= core_csr_newCfg_1_x ; 
                             core_csr_reg_pmp_1_cfg_w  <= core_csr__GEN_94 ; 
                             core_csr_reg_pmp_1_cfg_r  <= core_csr_newCfg_1_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_95 ) 
                         core_csr_reg_pmp_1_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_96 )
                         begin  
                             core_csr_reg_pmp_2_cfg_x  <= core_csr_newCfg_2_x ; 
                             core_csr_reg_pmp_2_cfg_w  <= core_csr__GEN_97 ; 
                             core_csr_reg_pmp_2_cfg_r  <= core_csr_newCfg_2_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_98 ) 
                         core_csr_reg_pmp_2_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_99 )
                         begin  
                             core_csr_reg_pmp_3_cfg_x  <= core_csr_newCfg_3_x ; 
                             core_csr_reg_pmp_3_cfg_w  <= core_csr__GEN_100 ; 
                             core_csr_reg_pmp_3_cfg_r  <= core_csr_newCfg_3_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_101 ) 
                         core_csr_reg_pmp_3_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_102 )
                         begin  
                             core_csr_reg_pmp_4_cfg_x  <= core_csr_newCfg_4_x ; 
                             core_csr_reg_pmp_4_cfg_w  <= core_csr__GEN_103 ; 
                             core_csr_reg_pmp_4_cfg_r  <= core_csr_newCfg_4_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_104 ) 
                         core_csr_reg_pmp_4_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_105 )
                         begin  
                             core_csr_reg_pmp_5_cfg_x  <= core_csr_newCfg_5_x ; 
                             core_csr_reg_pmp_5_cfg_w  <= core_csr__GEN_106 ; 
                             core_csr_reg_pmp_5_cfg_r  <= core_csr_newCfg_5_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_107 ) 
                         core_csr_reg_pmp_5_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_108 )
                         begin  
                             core_csr_reg_pmp_6_cfg_x  <= core_csr_newCfg_6_x ; 
                             core_csr_reg_pmp_6_cfg_w  <= core_csr__GEN_109 ; 
                             core_csr_reg_pmp_6_cfg_r  <= core_csr_newCfg_6_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_110 ) 
                         core_csr_reg_pmp_6_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_111 )
                         begin  
                             core_csr_reg_pmp_7_cfg_x  <= core_csr_newCfg_7_x ; 
                             core_csr_reg_pmp_7_cfg_w  <= core_csr__GEN_112 ; 
                             core_csr_reg_pmp_7_cfg_r  <= core_csr_newCfg_7_r ;
                         end 
                      else 
                         begin 
                         end 
                     if ( core_csr__GEN_113 ) 
                         core_csr_reg_pmp_7_addr  <= core_csr_wdata [29:0];
                      else 
                         begin 
                         end 
                     if ( core_csr_decoded_8 ) 
                         core_csr_reg_mie  <= core_csr__GEN_77 ;
                      else 
                         begin 
                         end 
                     if ( core_csr_decoded_10 ) 
                         core_csr_reg_mepc  <= core_csr__GEN_78 [33:0];
                      else 
                         if ( core_csr_exception )
                             begin 
                                 if ( core_csr_trapToDebug )
                                     begin 
                                     end 
                                  else 
                                     if ( core_csr_trapToNmiInt )
                                         begin 
                                         end 
                                      else 
                                         if ( core_csr__GEN_58 )
                                             begin 
                                             end 
                                          else 
                                             if ( core_csr__GEN_61 )
                                                 begin 
                                                 end 
                                              else  
                                                 core_csr_reg_mepc  <= core_csr_epc ;
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_decoded_11 ) 
                         core_csr_reg_mtval  <= core_csr_wdata [33:0];
                      else 
                         if ( core_csr_exception )
                             begin 
                                 if ( core_csr_trapToDebug )
                                     begin 
                                     end 
                                  else 
                                     if ( core_csr_trapToNmiInt )
                                         begin 
                                         end 
                                      else 
                                         if ( core_csr__GEN_58 )
                                             begin 
                                             end 
                                          else 
                                             if ( core_csr__GEN_61 )
                                                 begin 
                                                 end 
                                              else  
                                                 core_csr_reg_mtval  <= core_csr_tval ;
                             end 
                          else 
                             begin 
                             end 
                     if ( core_csr_decoded_9 ) 
                         core_csr_reg_mscratch  <= core_csr_wdata ;
                      else 
                         begin 
                         end 
                 end 
              else 
                 if ( core_csr_exception )
                     begin 
                         if ( core_csr_trapToDebug )
                             begin 
                                 if ( core_csr__GEN_51 ) 
                                     core_csr_reg_dpc  <= core_csr_epc ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             if ( core_csr_trapToNmiInt )
                                 begin 
                                 end 
                              else 
                                 if ( core_csr__GEN_58 )
                                     begin 
                                     end 
                                  else 
                                     if ( core_csr__GEN_61 )
                                         begin 
                                         end 
                                      else 
                                         begin  
                                             core_csr_reg_mepc  <= core_csr_epc ; 
                                             core_csr_reg_mtval  <= core_csr_tval ;
                                         end 
                     end 
                  else 
                     begin 
                     end 
             if ( core_csr__GEN_48 ) 
                 core_csr_reg_singleStepped  <=1'h0;
              else 
                 if ( core_csr__GEN_47 ) 
                     core_csr_reg_singleStepped  <=1'h1;
                  else 
                     begin 
                     end  
             core_csr_reg_tselect  <=1'h0; 
             core_csr_reg_bp_0_control_ttype  <=4'h2;
             if ( core_csr_reset )
                 begin  
                     core_csr_reg_bp_0_control_dmode  <=1'h0; 
                     core_csr_reg_bp_0_control_action  <=1'h0; 
                     core_csr_reg_bp_0_control_chain  <=1'h0; 
                     core_csr_reg_bp_0_control_x  <=1'h0; 
                     core_csr_reg_bp_0_control_w  <=1'h0; 
                     core_csr_reg_bp_0_control_r  <=1'h0; 
                     core_csr_reg_pmp_0_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_0_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_1_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_1_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_2_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_2_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_3_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_3_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_4_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_4_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_5_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_5_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_6_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_6_cfg_a  <=2'h0; 
                     core_csr_reg_pmp_7_cfg_l  <=1'h0; 
                     core_csr_reg_pmp_7_cfg_a  <=2'h0;
                 end 
              else 
                 if ( core_csr_csr_wen )
                     begin 
                         if ( core_csr__GEN_82 )
                             begin 
                                 if ( core_csr_decoded_1 )
                                     begin  
                                         core_csr_reg_bp_0_control_dmode  <= core_csr_dMode ;
                                         if ( core_csr__GEN_85 ) 
                                             core_csr_reg_bp_0_control_action  <= core_csr_newBPC_action ;
                                          else  
                                             core_csr_reg_bp_0_control_action  <=1'h0; 
                                         core_csr_reg_bp_0_control_chain  <=1'h0; 
                                         core_csr_reg_bp_0_control_x  <= core_csr__reg_bp_0_control_WIRE_x ; 
                                         core_csr_reg_bp_0_control_w  <= core_csr__reg_bp_0_control_WIRE_w ; 
                                         core_csr_reg_bp_0_control_r  <= core_csr__reg_bp_0_control_WIRE_r ;
                                     end 
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_90 )
                             begin  
                                 core_csr_reg_pmp_0_cfg_l  <= core_csr_newCfg_l ; 
                                 core_csr_reg_pmp_0_cfg_a  <= core_csr_newCfg_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_93 )
                             begin  
                                 core_csr_reg_pmp_1_cfg_l  <= core_csr_newCfg_1_l ; 
                                 core_csr_reg_pmp_1_cfg_a  <= core_csr_newCfg_1_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_96 )
                             begin  
                                 core_csr_reg_pmp_2_cfg_l  <= core_csr_newCfg_2_l ; 
                                 core_csr_reg_pmp_2_cfg_a  <= core_csr_newCfg_2_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_99 )
                             begin  
                                 core_csr_reg_pmp_3_cfg_l  <= core_csr_newCfg_3_l ; 
                                 core_csr_reg_pmp_3_cfg_a  <= core_csr_newCfg_3_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_102 )
                             begin  
                                 core_csr_reg_pmp_4_cfg_l  <= core_csr_newCfg_4_l ; 
                                 core_csr_reg_pmp_4_cfg_a  <= core_csr_newCfg_4_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_105 )
                             begin  
                                 core_csr_reg_pmp_5_cfg_l  <= core_csr_newCfg_5_l ; 
                                 core_csr_reg_pmp_5_cfg_a  <= core_csr_newCfg_5_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_108 )
                             begin  
                                 core_csr_reg_pmp_6_cfg_l  <= core_csr_newCfg_6_l ; 
                                 core_csr_reg_pmp_6_cfg_a  <= core_csr_newCfg_6_a ;
                             end 
                          else 
                             begin 
                             end 
                         if ( core_csr__GEN_111 )
                             begin  
                                 core_csr_reg_pmp_7_cfg_l  <= core_csr_newCfg_7_l ; 
                                 core_csr_reg_pmp_7_cfg_a  <= core_csr_newCfg_7_a ;
                             end 
                          else 
                             begin 
                             end 
                     end 
                  else 
                     begin 
                     end  
             core_csr_reg_bp_0_control_maskmax  <=6'h4; 
             core_csr_reg_bp_0_control_reserved  <=40'h0; 
             core_csr_reg_bp_0_control_zero  <=2'h0; 
             core_csr_reg_bp_0_control_m  <=1'h1; 
             core_csr_reg_bp_0_control_h  <=1'h0; 
             core_csr_reg_bp_0_control_s  <=1'h0; 
             core_csr_reg_bp_0_control_u  <=1'h0; 
             core_csr_reg_bp_0_textra_mselect  <=1'h0; 
             core_csr_reg_bp_0_textra_sselect  <=1'h0; 
             core_csr_reg_bp_1_control_ttype  <= core_csr__reg_bp_1_WIRE_control_ttype ; 
             core_csr_reg_bp_1_control_dmode  <= core_csr__reg_bp_1_WIRE_control_dmode ; 
             core_csr_reg_bp_1_control_maskmax  <= core_csr__reg_bp_1_WIRE_control_maskmax ; 
             core_csr_reg_bp_1_control_reserved  <= core_csr__reg_bp_1_WIRE_control_reserved ; 
             core_csr_reg_bp_1_control_action  <= core_csr__reg_bp_1_WIRE_control_action ; 
             core_csr_reg_bp_1_control_chain  <= core_csr__reg_bp_1_WIRE_control_chain ; 
             core_csr_reg_bp_1_control_zero  <= core_csr__reg_bp_1_WIRE_control_zero ; 
             core_csr_reg_bp_1_control_tmatch  <= core_csr__reg_bp_1_WIRE_control_tmatch ; 
             core_csr_reg_bp_1_control_m  <= core_csr__reg_bp_1_WIRE_control_m ; 
             core_csr_reg_bp_1_control_h  <= core_csr__reg_bp_1_WIRE_control_h ; 
             core_csr_reg_bp_1_control_s  <= core_csr__reg_bp_1_WIRE_control_s ; 
             core_csr_reg_bp_1_control_u  <= core_csr__reg_bp_1_WIRE_control_u ; 
             core_csr_reg_bp_1_control_x  <= core_csr__reg_bp_1_WIRE_control_x ; 
             core_csr_reg_bp_1_control_w  <= core_csr__reg_bp_1_WIRE_control_w ; 
             core_csr_reg_bp_1_control_r  <= core_csr__reg_bp_1_WIRE_control_r ; 
             core_csr_reg_bp_1_address  <= core_csr__reg_bp_1_WIRE_address ; 
             core_csr_reg_bp_1_textra_mselect  <= core_csr__reg_bp_1_WIRE_textra_mselect ; 
             core_csr_reg_bp_1_textra_pad2  <= core_csr__reg_bp_1_WIRE_textra_pad2 ; 
             core_csr_reg_bp_1_textra_pad1  <= core_csr__reg_bp_1_WIRE_textra_pad1 ; 
             core_csr_reg_bp_1_textra_sselect  <= core_csr__reg_bp_1_WIRE_textra_sselect ; 
             core_csr_reg_pmp_0_cfg_res  <=2'h0; 
             core_csr_reg_pmp_1_cfg_res  <=2'h0; 
             core_csr_reg_pmp_2_cfg_res  <=2'h0; 
             core_csr_reg_pmp_3_cfg_res  <=2'h0; 
             core_csr_reg_pmp_4_cfg_res  <=2'h0; 
             core_csr_reg_pmp_5_cfg_res  <=2'h0; 
             core_csr_reg_pmp_6_cfg_res  <=2'h0; 
             core_csr_reg_pmp_7_cfg_res  <=2'h0;
             if ( core_csr_exception )
                 begin 
                     if ( core_csr_trapToDebug )
                         begin 
                         end 
                      else 
                         if ( core_csr_trapToNmiInt )
                             begin 
                                 if ( core_csr_reg_rnmie ) 
                                     core_csr_reg_mnepc  <= core_csr_epc ;
                                  else 
                                     begin 
                                     end 
                             end 
                          else 
                             if ( core_csr__GEN_58 )
                                 begin  
                                     core_csr_reg_vsstatus_spp  <= core_csr_reg_mstatus_prv [0]; 
                                     core_csr_reg_vsstatus_spie  <= core_csr_reg_vsstatus_sie ; 
                                     core_csr_reg_vsstatus_sie  <=1'h0; 
                                     core_csr_reg_vsepc  <= core_csr_epc ; 
                                     core_csr_reg_vscause  <= core_csr__GEN_59 ; 
                                     core_csr_reg_vstval  <= core_csr_tval ;
                                 end 
                              else 
                                 if ( core_csr__GEN_61 )
                                     begin  
                                         core_csr_reg_htval  <= core_csr_io_htval ; 
                                         core_csr_reg_sepc  <= core_csr_epc ; 
                                         core_csr_reg_scause  <= core_csr_cause ; 
                                         core_csr_reg_stval  <= core_csr_tval ;
                                     end 
                                  else  
                                     core_csr_reg_mtval2  <= core_csr_io_htval ;
                 end 
              else 
                 begin 
                 end  
             core_csr_reg_hgatp_mode  <=4'h0; 
             core_csr_reg_hgatp_asid  <=16'h0; 
             core_csr_reg_hgatp_ppn  <=44'h0; 
             core_csr_reg_vsstatus_xs  <=2'h0; 
             core_csr_reg_vsatp_mode  <=4'h0; 
             core_csr_reg_vsatp_asid  <=16'h0; 
             core_csr_reg_vsatp_ppn  <=44'h0; 
             core_csr_reg_satp_mode  <=4'h0; 
             core_csr_reg_satp_asid  <=16'h0; 
             core_csr_reg_satp_ppn  <=44'h0;
             if ( core_csr_io_fcsr_flags_valid ) 
                 core_csr_reg_fflags  <= core_csr__GEN_73 ;
              else 
                 begin 
                 end 
         end
  always @( posedge  core_csr_io_ungated_clock )
         begin 
             if ( core_csr_reset )
                 begin  
                     core_csr_reg_wfi  <=1'h0; 
                     core_csr_small_1  <=6'h0; 
                     core_csr_large_1  <=58'h0;
                 end 
              else 
                 begin 
                     if ( core_csr__GEN_46 ) 
                         core_csr_reg_wfi  <=1'h0;
                      else 
                         if ( core_csr__GEN_45 ) 
                             core_csr_reg_wfi  <=1'h1;
                          else 
                             begin 
                             end 
                     if ( core_csr_csr_wen )
                         begin 
                             if ( core_csr_decoded_18 )
                                 begin  
                                     core_csr_small_1  <= core_csr_wdata [5:0]; 
                                     core_csr_large_1  <= core_csr_wdata [63:6];
                                 end 
                              else 
                                 begin 
                                     if ( core_csr__GEN_5 ) 
                                         core_csr_small_1  <= core_csr_nextSmall_1 [5:0];
                                      else 
                                         begin 
                                         end 
                                     if ( core_csr__GEN_7 ) 
                                         core_csr_large_1  <= core_csr__GEN_8 [57:0];
                                      else 
                                         begin 
                                         end 
                                 end 
                         end 
                      else 
                         begin 
                             if ( core_csr__GEN_5 ) 
                                 core_csr_small_1  <= core_csr_nextSmall_1 [5:0];
                              else 
                                 begin 
                                 end 
                             if ( core_csr__GEN_7 ) 
                                 core_csr_large_1  <= core_csr__GEN_8 [57:0];
                              else 
                                 begin 
                                 end 
                         end 
                 end 
         end
  assign  core_csr_io_rw_rdata = core_csr__io_rw_rdata_output ; 
  assign  core_csr_io_decode_0_fp_illegal = core_csr__io_decode_0_fp_illegal_output ; 
  assign  core_csr_io_decode_0_vector_illegal = core_csr__io_decode_0_vector_illegal_output ; 
  assign  core_csr_io_decode_0_fp_csr = core_csr__io_decode_0_fp_csr_output ; 
  assign  core_csr_io_decode_0_rocc_illegal = core_csr__io_status_xs_output ==2'h0| core_csr_reg_mstatus_v & core_csr_reg_vsstatus_xs ==2'h0| core_csr_reg_misa [23]==1'h0; 
  assign  core_csr_io_decode_0_read_illegal = core_csr_csr_addr_legal ==1'h0| core_csr_csr_exists ==1'h0|( core_csr_addr_1 ==12'h180| core_csr_addr_1 ==12'h680)& core_csr_allow_sfence_vma ==1'h0| core_csr_is_counter & core_csr_allow_counter ==1'h0| core_csr_io_decode_0_read_illegal_plaOutput & core_csr_reg_debug ==1'h0| core_csr_io_decode_0_read_illegal_plaOutput_1 & core_csr__io_decode_0_vector_illegal_output | core_csr__io_decode_0_fp_csr_output & core_csr__io_decode_0_fp_illegal_output ; 
  assign  core_csr_io_decode_0_write_illegal =&( core_csr_addr_1 [11:10]); 
  assign  core_csr_io_decode_0_write_flush =( core_csr_io_decode_0_write_flush_addr_m >=12'h340& core_csr_io_decode_0_write_flush_addr_m <=12'h343)==1'h0; 
  assign  core_csr_io_decode_0_system_illegal = core_csr_csr_addr_legal ==1'h0& core_csr_is_hlsv ==1'h0| core_csr_is_wfi & core_csr_allow_wfi ==1'h0| core_csr_is_ret & core_csr_allow_sret ==1'h0| core_csr_is_ret & core_csr_addr_1 [10]& core_csr_addr_1 [7]& core_csr_reg_debug ==1'h0|( core_csr_is_sfence | core_csr_is_hfence_gvma )& core_csr_allow_sfence_vma ==1'h0| core_csr_is_hfence_vvma & core_csr_allow_hfence_vvma ==1'h0| core_csr_is_hlsv & core_csr_allow_hlsv ==1'h0; 
  assign  core_csr_io_decode_0_virtual_access_illegal = core_csr_reg_mstatus_v & core_csr_csr_exists &( core_csr_addr_1 [9:8]==2'h2| core_csr_is_counter & core_csr__GEN_35 [0]&( core_csr__GEN_36 [0]==1'h0| core_csr_reg_mstatus_prv [0]==1'h0& core_csr__GEN_37 [0]==1'h0)| core_csr_addr_1 [9:8]==2'h1& core_csr_reg_mstatus_prv [0]==1'h0| core_csr_addr_1 ==12'h180& core_csr_reg_mstatus_prv [0]& core_csr_reg_hstatus_vtvm ); 
  assign  core_csr_io_decode_0_virtual_system_illegal = core_csr_reg_mstatus_v &( core_csr_is_hfence_vvma | core_csr_is_hfence_gvma | core_csr_is_hlsv | core_csr_is_wfi &( core_csr_reg_mstatus_prv [0]==1'h0| core_csr_reg_mstatus_tw ==1'h0& core_csr_reg_hstatus_vtw )| core_csr_is_ret & core_csr_addr_1 [9:8]==2'h1&( core_csr_reg_mstatus_prv [0]==1'h0| core_csr_reg_hstatus_vtsr )| core_csr_is_sfence &( core_csr_reg_mstatus_prv [0]==1'h0| core_csr_reg_hstatus_vtvm )); 
  assign  core_csr_io_csr_stall = core_csr__io_csr_stall_output ; 
  assign  core_csr_io_rw_stall = core_csr__io_rw_stall_output ; 
  assign  core_csr_io_eret = core_csr_insn_call | core_csr_insn_break | core_csr_insn_ret ; 
  assign  core_csr_io_singleStep = core_csr__io_singleStep_output ; 
  assign  core_csr_io_status_debug = core_csr__io_status_debug_output ; 
  assign  core_csr_io_status_cease = core_csr__io_status_cease_output ; 
  assign  core_csr_io_status_wfi = core_csr__io_status_wfi_output ; 
  assign  core_csr_io_status_isa = core_csr__io_status_isa_output ; 
  assign  core_csr_io_status_dprv = core_csr__io_status_dprv_output ; 
  assign  core_csr_io_status_dv = core_csr__io_status_dv_output ; 
  assign  core_csr_io_status_prv = core_csr__io_status_prv_output ; 
  assign  core_csr_io_status_v = core_csr__io_status_v_output ; 
  assign  core_csr_io_status_sd = core_csr__io_status_sd_output ; 
  assign  core_csr_io_status_zero2 = core_csr__io_status_zero2_output ; 
  assign  core_csr_io_status_mpv = core_csr__io_status_mpv_output ; 
  assign  core_csr_io_status_gva = core_csr__io_status_gva_output ; 
  assign  core_csr_io_status_mbe = core_csr__io_status_mbe_output ; 
  assign  core_csr_io_status_sbe = core_csr__io_status_sbe_output ; 
  assign  core_csr_io_status_sxl = core_csr__io_status_sxl_output ; 
  assign  core_csr_io_status_uxl = core_csr__io_status_uxl_output ; 
  assign  core_csr_io_status_sd_rv32 = core_csr__io_status_sd_rv32_output ; 
  assign  core_csr_io_status_zero1 = core_csr__io_status_zero1_output ; 
  assign  core_csr_io_status_tsr = core_csr__io_status_tsr_output ; 
  assign  core_csr_io_status_tw = core_csr__io_status_tw_output ; 
  assign  core_csr_io_status_tvm = core_csr__io_status_tvm_output ; 
  assign  core_csr_io_status_mxr = core_csr__io_status_mxr_output ; 
  assign  core_csr_io_status_sum = core_csr__io_status_sum_output ; 
  assign  core_csr_io_status_mprv = core_csr__io_status_mprv_output ; 
  assign  core_csr_io_status_xs = core_csr__io_status_xs_output ; 
  assign  core_csr_io_status_fs = core_csr__io_status_fs_output ; 
  assign  core_csr_io_status_mpp = core_csr__io_status_mpp_output ; 
  assign  core_csr_io_status_vs = core_csr__io_status_vs_output ; 
  assign  core_csr_io_status_spp = core_csr__io_status_spp_output ; 
  assign  core_csr_io_status_mpie = core_csr__io_status_mpie_output ; 
  assign  core_csr_io_status_ube = core_csr__io_status_ube_output ; 
  assign  core_csr_io_status_spie = core_csr__io_status_spie_output ; 
  assign  core_csr_io_status_upie = core_csr__io_status_upie_output ; 
  assign  core_csr_io_status_mie = core_csr__io_status_mie_output ; 
  assign  core_csr_io_status_hie = core_csr__io_status_hie_output ; 
  assign  core_csr_io_status_sie = core_csr__io_status_sie_output ; 
  assign  core_csr_io_status_uie = core_csr__io_status_uie_output ; 
  assign  core_csr_io_hstatus_zero6 = core_csr_reg_hstatus_zero6 ; 
  assign  core_csr_io_hstatus_vsxl =2'h0; 
  assign  core_csr_io_hstatus_zero5 = core_csr_reg_hstatus_zero5 ; 
  assign  core_csr_io_hstatus_vtsr = core_csr_reg_hstatus_vtsr ; 
  assign  core_csr_io_hstatus_vtw = core_csr_reg_hstatus_vtw ; 
  assign  core_csr_io_hstatus_vtvm = core_csr_reg_hstatus_vtvm ; 
  assign  core_csr_io_hstatus_zero3 = core_csr_reg_hstatus_zero3 ; 
  assign  core_csr_io_hstatus_vgein = core_csr_reg_hstatus_vgein ; 
  assign  core_csr_io_hstatus_zero2 = core_csr_reg_hstatus_zero2 ; 
  assign  core_csr_io_hstatus_hu = core_csr_reg_hstatus_hu ; 
  assign  core_csr_io_hstatus_spvp = core_csr_reg_hstatus_spvp ; 
  assign  core_csr_io_hstatus_spv = core_csr_reg_hstatus_spv ; 
  assign  core_csr_io_hstatus_gva = core_csr_reg_hstatus_gva ; 
  assign  core_csr_io_hstatus_vsbe = core_csr_reg_hstatus_vsbe ; 
  assign  core_csr_io_hstatus_zero1 = core_csr_reg_hstatus_zero1 ; 
  assign  core_csr_io_gstatus_debug = core_csr_reg_vsstatus_debug ; 
  assign  core_csr_io_gstatus_cease = core_csr_reg_vsstatus_cease ; 
  assign  core_csr_io_gstatus_wfi = core_csr_reg_vsstatus_wfi ; 
  assign  core_csr_io_gstatus_isa = core_csr_reg_vsstatus_isa ; 
  assign  core_csr_io_gstatus_dprv = core_csr_reg_vsstatus_dprv ; 
  assign  core_csr_io_gstatus_dv = core_csr_reg_vsstatus_dv ; 
  assign  core_csr_io_gstatus_prv = core_csr_reg_vsstatus_prv ; 
  assign  core_csr_io_gstatus_v = core_csr_reg_vsstatus_v ; 
  assign  core_csr_io_gstatus_sd = core_csr__io_gstatus_sd_output ; 
  assign  core_csr_io_gstatus_zero2 = core_csr_reg_vsstatus_zero2 ; 
  assign  core_csr_io_gstatus_mpv = core_csr_reg_vsstatus_mpv ; 
  assign  core_csr_io_gstatus_gva = core_csr_reg_vsstatus_gva ; 
  assign  core_csr_io_gstatus_mbe = core_csr_reg_vsstatus_mbe ; 
  assign  core_csr_io_gstatus_sbe = core_csr_reg_vsstatus_sbe ; 
  assign  core_csr_io_gstatus_sxl = core_csr_reg_vsstatus_sxl ; 
  assign  core_csr_io_gstatus_uxl =2'h0; 
  assign  core_csr_io_gstatus_sd_rv32 =1'h0; 
  assign  core_csr_io_gstatus_zero1 = core_csr_reg_vsstatus_zero1 ; 
  assign  core_csr_io_gstatus_tsr = core_csr_reg_vsstatus_tsr ; 
  assign  core_csr_io_gstatus_tw = core_csr_reg_vsstatus_tw ; 
  assign  core_csr_io_gstatus_tvm = core_csr_reg_vsstatus_tvm ; 
  assign  core_csr_io_gstatus_mxr = core_csr_reg_vsstatus_mxr ; 
  assign  core_csr_io_gstatus_sum = core_csr_reg_vsstatus_sum ; 
  assign  core_csr_io_gstatus_mprv = core_csr_reg_vsstatus_mprv ; 
  assign  core_csr_io_gstatus_xs = core_csr__io_gstatus_xs_output ; 
  assign  core_csr_io_gstatus_fs = core_csr__io_gstatus_fs_output ; 
  assign  core_csr_io_gstatus_mpp = core_csr_reg_vsstatus_mpp ; 
  assign  core_csr_io_gstatus_vs = core_csr__io_gstatus_vs_output ; 
  assign  core_csr_io_gstatus_spp = core_csr_reg_vsstatus_spp ; 
  assign  core_csr_io_gstatus_mpie = core_csr_reg_vsstatus_mpie ; 
  assign  core_csr_io_gstatus_ube = core_csr_reg_vsstatus_ube ; 
  assign  core_csr_io_gstatus_spie = core_csr_reg_vsstatus_spie ; 
  assign  core_csr_io_gstatus_upie = core_csr_reg_vsstatus_upie ; 
  assign  core_csr_io_gstatus_mie = core_csr_reg_vsstatus_mie ; 
  assign  core_csr_io_gstatus_hie = core_csr_reg_vsstatus_hie ; 
  assign  core_csr_io_gstatus_sie = core_csr_reg_vsstatus_sie ; 
  assign  core_csr_io_gstatus_uie = core_csr_reg_vsstatus_uie ; 
  assign  core_csr_io_ptbr_mode = core_csr_reg_satp_mode ; 
  assign  core_csr_io_ptbr_asid = core_csr_reg_satp_asid ; 
  assign  core_csr_io_ptbr_ppn = core_csr_reg_satp_ppn ; 
  assign  core_csr_io_hgatp_mode = core_csr_reg_hgatp_mode ; 
  assign  core_csr_io_hgatp_asid = core_csr_reg_hgatp_asid ; 
  assign  core_csr_io_hgatp_ppn = core_csr_reg_hgatp_ppn ; 
  assign  core_csr_io_vsatp_mode = core_csr_reg_vsatp_mode ; 
  assign  core_csr_io_vsatp_asid = core_csr_reg_vsatp_asid ; 
  assign  core_csr_io_vsatp_ppn = core_csr_reg_vsatp_ppn ; 
  assign  core_csr_io_evec = core_csr_insn_ret  ? ( core_csr__GEN_70  ? ~(~ core_csr_reg_dpc |{32'h0, core_csr_reg_misa [2] ? 2'h1:2'h3}):~(~ core_csr_reg_mepc |{32'h0, core_csr_reg_misa [2] ? 2'h1:2'h3})): core_csr_tvec [33:0]; 
  assign  core_csr_io_time = core_csr_value_1 ; 
  assign  core_csr_io_fcsr_rm = core_csr_reg_frm ; 
  assign  core_csr_io_interrupt =( core_csr_anyInterrupt & core_csr__io_singleStep_output ==1'h0| core_csr_reg_singleStepped )&( core_csr_reg_debug | core_csr__io_status_cease_output )==1'h0; 
  assign  core_csr_io_interrupt_cause = core_csr_interruptCause ; 
  assign  core_csr_io_bp_0_control_ttype = core_csr_reg_bp_0_control_ttype ; 
  assign  core_csr_io_bp_0_control_dmode = core_csr_reg_bp_0_control_dmode ; 
  assign  core_csr_io_bp_0_control_maskmax = core_csr_reg_bp_0_control_maskmax ; 
  assign  core_csr_io_bp_0_control_reserved = core_csr_reg_bp_0_control_reserved ; 
  assign  core_csr_io_bp_0_control_action = core_csr_reg_bp_0_control_action ; 
  assign  core_csr_io_bp_0_control_chain = core_csr_reg_bp_0_control_chain ; 
  assign  core_csr_io_bp_0_control_zero = core_csr_reg_bp_0_control_zero ; 
  assign  core_csr_io_bp_0_control_tmatch = core_csr_reg_bp_0_control_tmatch ; 
  assign  core_csr_io_bp_0_control_m = core_csr_reg_bp_0_control_m ; 
  assign  core_csr_io_bp_0_control_h = core_csr_reg_bp_0_control_h ; 
  assign  core_csr_io_bp_0_control_s = core_csr_reg_bp_0_control_s ; 
  assign  core_csr_io_bp_0_control_u = core_csr_reg_bp_0_control_u ; 
  assign  core_csr_io_bp_0_control_x = core_csr_reg_bp_0_control_x ; 
  assign  core_csr_io_bp_0_control_w = core_csr_reg_bp_0_control_w ; 
  assign  core_csr_io_bp_0_control_r = core_csr_reg_bp_0_control_r ; 
  assign  core_csr_io_bp_0_address = core_csr_reg_bp_0_address ; 
  assign  core_csr_io_bp_0_textra_mselect = core_csr_reg_bp_0_textra_mselect ; 
  assign  core_csr_io_bp_0_textra_pad2 = core_csr_reg_bp_0_textra_pad2 ; 
  assign  core_csr_io_bp_0_textra_pad1 = core_csr_reg_bp_0_textra_pad1 ; 
  assign  core_csr_io_bp_0_textra_sselect = core_csr_reg_bp_0_textra_sselect ; 
  assign  core_csr_io_pmp_0_cfg_l = core_csr_pmp_cfg_l ; 
  assign  core_csr_io_pmp_0_cfg_res = core_csr_pmp_cfg_res ; 
  assign  core_csr_io_pmp_0_cfg_a = core_csr_pmp_cfg_a ; 
  assign  core_csr_io_pmp_0_cfg_x = core_csr_pmp_cfg_x ; 
  assign  core_csr_io_pmp_0_cfg_w = core_csr_pmp_cfg_w ; 
  assign  core_csr_io_pmp_0_cfg_r = core_csr_pmp_cfg_r ; 
  assign  core_csr_io_pmp_0_addr = core_csr_pmp_addr ; 
  assign  core_csr_io_pmp_0_mask = core_csr_pmp_mask ; 
  assign  core_csr_io_pmp_1_cfg_l = core_csr_pmp_1_cfg_l ; 
  assign  core_csr_io_pmp_1_cfg_res = core_csr_pmp_1_cfg_res ; 
  assign  core_csr_io_pmp_1_cfg_a = core_csr_pmp_1_cfg_a ; 
  assign  core_csr_io_pmp_1_cfg_x = core_csr_pmp_1_cfg_x ; 
  assign  core_csr_io_pmp_1_cfg_w = core_csr_pmp_1_cfg_w ; 
  assign  core_csr_io_pmp_1_cfg_r = core_csr_pmp_1_cfg_r ; 
  assign  core_csr_io_pmp_1_addr = core_csr_pmp_1_addr ; 
  assign  core_csr_io_pmp_1_mask = core_csr_pmp_1_mask ; 
  assign  core_csr_io_pmp_2_cfg_l = core_csr_pmp_2_cfg_l ; 
  assign  core_csr_io_pmp_2_cfg_res = core_csr_pmp_2_cfg_res ; 
  assign  core_csr_io_pmp_2_cfg_a = core_csr_pmp_2_cfg_a ; 
  assign  core_csr_io_pmp_2_cfg_x = core_csr_pmp_2_cfg_x ; 
  assign  core_csr_io_pmp_2_cfg_w = core_csr_pmp_2_cfg_w ; 
  assign  core_csr_io_pmp_2_cfg_r = core_csr_pmp_2_cfg_r ; 
  assign  core_csr_io_pmp_2_addr = core_csr_pmp_2_addr ; 
  assign  core_csr_io_pmp_2_mask = core_csr_pmp_2_mask ; 
  assign  core_csr_io_pmp_3_cfg_l = core_csr_pmp_3_cfg_l ; 
  assign  core_csr_io_pmp_3_cfg_res = core_csr_pmp_3_cfg_res ; 
  assign  core_csr_io_pmp_3_cfg_a = core_csr_pmp_3_cfg_a ; 
  assign  core_csr_io_pmp_3_cfg_x = core_csr_pmp_3_cfg_x ; 
  assign  core_csr_io_pmp_3_cfg_w = core_csr_pmp_3_cfg_w ; 
  assign  core_csr_io_pmp_3_cfg_r = core_csr_pmp_3_cfg_r ; 
  assign  core_csr_io_pmp_3_addr = core_csr_pmp_3_addr ; 
  assign  core_csr_io_pmp_3_mask = core_csr_pmp_3_mask ; 
  assign  core_csr_io_pmp_4_cfg_l = core_csr_pmp_4_cfg_l ; 
  assign  core_csr_io_pmp_4_cfg_res = core_csr_pmp_4_cfg_res ; 
  assign  core_csr_io_pmp_4_cfg_a = core_csr_pmp_4_cfg_a ; 
  assign  core_csr_io_pmp_4_cfg_x = core_csr_pmp_4_cfg_x ; 
  assign  core_csr_io_pmp_4_cfg_w = core_csr_pmp_4_cfg_w ; 
  assign  core_csr_io_pmp_4_cfg_r = core_csr_pmp_4_cfg_r ; 
  assign  core_csr_io_pmp_4_addr = core_csr_pmp_4_addr ; 
  assign  core_csr_io_pmp_4_mask = core_csr_pmp_4_mask ; 
  assign  core_csr_io_pmp_5_cfg_l = core_csr_pmp_5_cfg_l ; 
  assign  core_csr_io_pmp_5_cfg_res = core_csr_pmp_5_cfg_res ; 
  assign  core_csr_io_pmp_5_cfg_a = core_csr_pmp_5_cfg_a ; 
  assign  core_csr_io_pmp_5_cfg_x = core_csr_pmp_5_cfg_x ; 
  assign  core_csr_io_pmp_5_cfg_w = core_csr_pmp_5_cfg_w ; 
  assign  core_csr_io_pmp_5_cfg_r = core_csr_pmp_5_cfg_r ; 
  assign  core_csr_io_pmp_5_addr = core_csr_pmp_5_addr ; 
  assign  core_csr_io_pmp_5_mask = core_csr_pmp_5_mask ; 
  assign  core_csr_io_pmp_6_cfg_l = core_csr_pmp_6_cfg_l ; 
  assign  core_csr_io_pmp_6_cfg_res = core_csr_pmp_6_cfg_res ; 
  assign  core_csr_io_pmp_6_cfg_a = core_csr_pmp_6_cfg_a ; 
  assign  core_csr_io_pmp_6_cfg_x = core_csr_pmp_6_cfg_x ; 
  assign  core_csr_io_pmp_6_cfg_w = core_csr_pmp_6_cfg_w ; 
  assign  core_csr_io_pmp_6_cfg_r = core_csr_pmp_6_cfg_r ; 
  assign  core_csr_io_pmp_6_addr = core_csr_pmp_6_addr ; 
  assign  core_csr_io_pmp_6_mask = core_csr_pmp_6_mask ; 
  assign  core_csr_io_pmp_7_cfg_l = core_csr_pmp_7_cfg_l ; 
  assign  core_csr_io_pmp_7_cfg_res = core_csr_pmp_7_cfg_res ; 
  assign  core_csr_io_pmp_7_cfg_a = core_csr_pmp_7_cfg_a ; 
  assign  core_csr_io_pmp_7_cfg_x = core_csr_pmp_7_cfg_x ; 
  assign  core_csr_io_pmp_7_cfg_w = core_csr_pmp_7_cfg_w ; 
  assign  core_csr_io_pmp_7_cfg_r = core_csr_pmp_7_cfg_r ; 
  assign  core_csr_io_pmp_7_addr = core_csr_pmp_7_addr ; 
  assign  core_csr_io_pmp_7_mask = core_csr_pmp_7_mask ; 
  assign  core_csr_io_csrw_counter = core_csr_csr_wen &1'h1&( core_csr_io_rw_addr >=12'hB00& core_csr_io_rw_addr <12'hB20| core_csr_io_rw_addr >=12'hB80& core_csr_io_rw_addr <12'hBA0) ? 32'h1<< core_csr_io_rw_addr [4:0]:32'h0; 
  assign  core_csr_io_inhibit_cycle = core_csr_reg_mcountinhibit [0]; 
  assign  core_csr_io_trace_0_valid = core_csr_io_retire >1'h0| core_csr__io_trace_0_exception_output ; 
  assign  core_csr_io_trace_0_iaddr = core_csr_io_pc ; 
  assign  core_csr_io_trace_0_insn = core_csr_io_inst_0 ; 
  assign  core_csr_io_trace_0_priv ={ core_csr_reg_debug , core_csr_reg_mstatus_prv }; 
  assign  core_csr_io_trace_0_exception = core_csr__io_trace_0_exception_output ; 
  assign  core_csr_io_trace_0_interrupt = core_csr_cause [63]; 
  assign  core_csr_io_trace_0_cause = core_csr_cause ; 
  assign  core_csr_io_trace_0_tval = core_csr_io_tval ; 
  assign  core_csr_io_fiom = core_csr_reg_mstatus_prv <2'h3& core_csr_reg_menvcfg_fiom | core_csr_reg_mstatus_prv <2'h1& core_csr_reg_senvcfg_fiom | core_csr_reg_mstatus_v & core_csr_reg_henvcfg_fiom ; 
  assign  core_csr_io_customCSRs_0_ren = core_csr_reg_custom_read ; 
  assign  core_csr_io_customCSRs_0_wen = core_csr_csr_wen  ?  core_csr_decoded_127 :1'h0; 
  assign  core_csr_io_customCSRs_0_wdata = core_csr_wdata ; 
  assign  core_csr_io_customCSRs_0_value = core_csr_reg_custom_0 ; 
  assign  core_csr_io_customCSRs_1_ren = core_csr_reg_custom_read_1 ; 
  assign  core_csr_io_customCSRs_1_wen = core_csr_csr_wen  ?  core_csr_decoded_128 :1'h0; 
  assign  core_csr_io_customCSRs_1_wdata = core_csr_wdata ; 
  assign  core_csr_io_customCSRs_1_value = core_csr_reg_custom_1 ; 
  assign  core_csr_io_customCSRs_2_ren = core_csr_reg_custom_read_2 ; 
  assign  core_csr_io_customCSRs_2_wen = core_csr_csr_wen  ?  core_csr_decoded_129 :1'h0; 
  assign  core_csr_io_customCSRs_2_wdata = core_csr_wdata ; 
  assign  core_csr_io_customCSRs_2_value = core_csr_reg_custom_2 ; 
  assign  core_csr_io_customCSRs_3_ren = core_csr_reg_custom_read_3 ; 
  assign  core_csr_io_customCSRs_3_wen = core_csr_csr_wen  ?  core_csr_decoded_130 :1'h0; 
  assign  core_csr_io_customCSRs_3_wdata = core_csr_wdata ; 
  assign  core_csr_io_customCSRs_3_value = core_csr_reg_custom_3 ;
    assign core_csr_clock = core_clock;
    assign core_csr_reset = core_reset;
    assign core_csr_io_ungated_clock = core_clock;
    assign core_csr_io_interrupts_debug = core_io_interrupts_debug;
    assign core_csr_io_interrupts_mtip = core_io_interrupts_mtip;
    assign core_csr_io_interrupts_msip = core_io_interrupts_msip;
    assign core_csr_io_interrupts_meip = core_io_interrupts_meip;
    assign core_csr_io_hartid = core_io_hartid;
    assign core_csr_io_rw_addr = core__wb_reg_inst_31to20;
    assign core_csr_io_rw_cmd = core__GEN_0;
    assign core__csr_io_rw_rdata = core_csr_io_rw_rdata;
    assign core_csr_io_rw_wdata = core_wb_reg_wdata;
    assign core_csr_io_decode_0_inst = core__ibuf_io_inst_0_bits_inst_bits;
    assign core__csr_io_decode_0_fp_illegal = core_csr_io_decode_0_fp_illegal;
    assign core__csr_io_decode_0_fp_csr = core_csr_io_decode_0_fp_csr;
    assign core__csr_io_decode_0_rocc_illegal = core_csr_io_decode_0_rocc_illegal;
    assign core__csr_io_decode_0_read_illegal = core_csr_io_decode_0_read_illegal;
    assign core__csr_io_decode_0_write_illegal = core_csr_io_decode_0_write_illegal;
    assign core__csr_io_decode_0_write_flush = core_csr_io_decode_0_write_flush;
    assign core__csr_io_decode_0_system_illegal = core_csr_io_decode_0_system_illegal;
    assign core__csr_io_decode_0_virtual_access_illegal = core_csr_io_decode_0_virtual_access_illegal;
    assign core__csr_io_decode_0_virtual_system_illegal = core_csr_io_decode_0_virtual_system_illegal;
    assign core__csr_io_csr_stall = core_csr_io_csr_stall;
    assign core__csr_io_rw_stall = core_csr_io_rw_stall;
    assign core__csr_io_eret = core_csr_io_eret;
    assign core__csr_io_singleStep = core_csr_io_singleStep;
    assign core__csr_io_status_debug = core_csr_io_status_debug;
    assign core__csr_io_status_cease = core_csr_io_status_cease;
    assign core__csr_io_status_wfi = core_csr_io_status_wfi;
    assign core__csr_io_status_isa = core_csr_io_status_isa;
    assign core__csr_io_status_dprv = core_csr_io_status_dprv;
    assign core__csr_io_status_dv = core_csr_io_status_dv;
    assign core__csr_io_status_prv = core_csr_io_status_prv;
    assign core__csr_io_status_v = core_csr_io_status_v;
    assign core__csr_io_status_sd = core_csr_io_status_sd;
    assign core__csr_io_status_zero2 = core_csr_io_status_zero2;
    assign core__csr_io_status_mpv = core_csr_io_status_mpv;
    assign core__csr_io_status_gva = core_csr_io_status_gva;
    assign core__csr_io_status_mbe = core_csr_io_status_mbe;
    assign core__csr_io_status_sbe = core_csr_io_status_sbe;
    assign core__csr_io_status_sxl = core_csr_io_status_sxl;
    assign core__csr_io_status_uxl = core_csr_io_status_uxl;
    assign core__csr_io_status_sd_rv32 = core_csr_io_status_sd_rv32;
    assign core__csr_io_status_zero1 = core_csr_io_status_zero1;
    assign core__csr_io_status_tsr = core_csr_io_status_tsr;
    assign core__csr_io_status_tw = core_csr_io_status_tw;
    assign core__csr_io_status_tvm = core_csr_io_status_tvm;
    assign core__csr_io_status_mxr = core_csr_io_status_mxr;
    assign core__csr_io_status_sum = core_csr_io_status_sum;
    assign core__csr_io_status_mprv = core_csr_io_status_mprv;
    assign core__csr_io_status_xs = core_csr_io_status_xs;
    assign core__csr_io_status_fs = core_csr_io_status_fs;
    assign core__csr_io_status_mpp = core_csr_io_status_mpp;
    assign core__csr_io_status_vs = core_csr_io_status_vs;
    assign core__csr_io_status_spp = core_csr_io_status_spp;
    assign core__csr_io_status_mpie = core_csr_io_status_mpie;
    assign core__csr_io_status_ube = core_csr_io_status_ube;
    assign core__csr_io_status_spie = core_csr_io_status_spie;
    assign core__csr_io_status_upie = core_csr_io_status_upie;
    assign core__csr_io_status_mie = core_csr_io_status_mie;
    assign core__csr_io_status_hie = core_csr_io_status_hie;
    assign core__csr_io_status_sie = core_csr_io_status_sie;
    assign core__csr_io_status_uie = core_csr_io_status_uie;
    assign core_io_ptw_hstatus_zero6 = core_csr_io_hstatus_zero6;
    assign core_io_ptw_hstatus_vsxl = core_csr_io_hstatus_vsxl;
    assign core_io_ptw_hstatus_zero5 = core_csr_io_hstatus_zero5;
    assign core_io_ptw_hstatus_vtsr = core_csr_io_hstatus_vtsr;
    assign core_io_ptw_hstatus_vtw = core_csr_io_hstatus_vtw;
    assign core_io_ptw_hstatus_vtvm = core_csr_io_hstatus_vtvm;
    assign core_io_ptw_hstatus_zero3 = core_csr_io_hstatus_zero3;
    assign core_io_ptw_hstatus_vgein = core_csr_io_hstatus_vgein;
    assign core_io_ptw_hstatus_zero2 = core_csr_io_hstatus_zero2;
    assign core_io_ptw_hstatus_hu = core_csr_io_hstatus_hu;
    assign core__csr_io_hstatus_spvp = core_csr_io_hstatus_spvp;
    assign core_io_ptw_hstatus_spv = core_csr_io_hstatus_spv;
    assign core_io_ptw_hstatus_gva = core_csr_io_hstatus_gva;
    assign core_io_ptw_hstatus_vsbe = core_csr_io_hstatus_vsbe;
    assign core_io_ptw_hstatus_zero1 = core_csr_io_hstatus_zero1;
    assign core_io_ptw_gstatus_debug = core_csr_io_gstatus_debug;
    assign core_io_ptw_gstatus_cease = core_csr_io_gstatus_cease;
    assign core_io_ptw_gstatus_wfi = core_csr_io_gstatus_wfi;
    assign core_io_ptw_gstatus_isa = core_csr_io_gstatus_isa;
    assign core_io_ptw_gstatus_dprv = core_csr_io_gstatus_dprv;
    assign core_io_ptw_gstatus_dv = core_csr_io_gstatus_dv;
    assign core_io_ptw_gstatus_prv = core_csr_io_gstatus_prv;
    assign core_io_ptw_gstatus_v = core_csr_io_gstatus_v;
    assign core_io_ptw_gstatus_sd = core_csr_io_gstatus_sd;
    assign core_io_ptw_gstatus_zero2 = core_csr_io_gstatus_zero2;
    assign core_io_ptw_gstatus_mpv = core_csr_io_gstatus_mpv;
    assign core_io_ptw_gstatus_gva = core_csr_io_gstatus_gva;
    assign core_io_ptw_gstatus_mbe = core_csr_io_gstatus_mbe;
    assign core_io_ptw_gstatus_sbe = core_csr_io_gstatus_sbe;
    assign core_io_ptw_gstatus_sxl = core_csr_io_gstatus_sxl;
    assign core_io_ptw_gstatus_uxl = core_csr_io_gstatus_uxl;
    assign core_io_ptw_gstatus_sd_rv32 = core_csr_io_gstatus_sd_rv32;
    assign core_io_ptw_gstatus_zero1 = core_csr_io_gstatus_zero1;
    assign core_io_ptw_gstatus_tsr = core_csr_io_gstatus_tsr;
    assign core_io_ptw_gstatus_tw = core_csr_io_gstatus_tw;
    assign core_io_ptw_gstatus_tvm = core_csr_io_gstatus_tvm;
    assign core_io_ptw_gstatus_mxr = core_csr_io_gstatus_mxr;
    assign core_io_ptw_gstatus_sum = core_csr_io_gstatus_sum;
    assign core_io_ptw_gstatus_mprv = core_csr_io_gstatus_mprv;
    assign core_io_ptw_gstatus_xs = core_csr_io_gstatus_xs;
    assign core_io_ptw_gstatus_fs = core_csr_io_gstatus_fs;
    assign core_io_ptw_gstatus_mpp = core_csr_io_gstatus_mpp;
    assign core_io_ptw_gstatus_vs = core_csr_io_gstatus_vs;
    assign core_io_ptw_gstatus_spp = core_csr_io_gstatus_spp;
    assign core_io_ptw_gstatus_mpie = core_csr_io_gstatus_mpie;
    assign core_io_ptw_gstatus_ube = core_csr_io_gstatus_ube;
    assign core_io_ptw_gstatus_spie = core_csr_io_gstatus_spie;
    assign core_io_ptw_gstatus_upie = core_csr_io_gstatus_upie;
    assign core_io_ptw_gstatus_mie = core_csr_io_gstatus_mie;
    assign core_io_ptw_gstatus_hie = core_csr_io_gstatus_hie;
    assign core_io_ptw_gstatus_sie = core_csr_io_gstatus_sie;
    assign core_io_ptw_gstatus_uie = core_csr_io_gstatus_uie;
    assign core_io_ptw_ptbr_mode = core_csr_io_ptbr_mode;
    assign core_io_ptw_ptbr_asid = core_csr_io_ptbr_asid;
    assign core_io_ptw_ptbr_ppn = core_csr_io_ptbr_ppn;
    assign core_io_ptw_hgatp_mode = core_csr_io_hgatp_mode;
    assign core_io_ptw_hgatp_asid = core_csr_io_hgatp_asid;
    assign core_io_ptw_hgatp_ppn = core_csr_io_hgatp_ppn;
    assign core_io_ptw_vsatp_mode = core_csr_io_vsatp_mode;
    assign core_io_ptw_vsatp_asid = core_csr_io_vsatp_asid;
    assign core_io_ptw_vsatp_ppn = core_csr_io_vsatp_ppn;
    assign core__csr_io_evec = core_csr_io_evec;
    assign core_csr_io_exception = core_wb_xcpt;
    assign core_csr_io_retire = core_wb_valid;
    assign core_csr_io_cause = core_wb_cause;
    assign core_csr_io_pc = core_wb_reg_pc;
    assign core_csr_io_tval = core__GEN_2;
    assign core_csr_io_htval = core__GEN_1;
    assign core_csr_io_gva = core__GEN_3;
    assign core__csr_io_time = core_csr_io_time;
    assign core_io_fpu_fcsr_rm = core_csr_io_fcsr_rm;
    assign core_csr_io_fcsr_flags_valid = core_io_fpu_fcsr_flags_valid;
    assign core_csr_io_fcsr_flags_bits = core_io_fpu_fcsr_flags_bits;
    assign core_csr_io_rocc_interrupt = core_io_rocc_interrupt;
    assign core__csr_io_interrupt = core_csr_io_interrupt;
    assign core__csr_io_interrupt_cause = core_csr_io_interrupt_cause;
    assign core__csr_io_bp_0_control_ttype = core_csr_io_bp_0_control_ttype;
    assign core__csr_io_bp_0_control_dmode = core_csr_io_bp_0_control_dmode;
    assign core__csr_io_bp_0_control_maskmax = core_csr_io_bp_0_control_maskmax;
    assign core__csr_io_bp_0_control_reserved = core_csr_io_bp_0_control_reserved;
    assign core__csr_io_bp_0_control_action = core_csr_io_bp_0_control_action;
    assign core__csr_io_bp_0_control_chain = core_csr_io_bp_0_control_chain;
    assign core__csr_io_bp_0_control_zero = core_csr_io_bp_0_control_zero;
    assign core__csr_io_bp_0_control_tmatch = core_csr_io_bp_0_control_tmatch;
    assign core__csr_io_bp_0_control_m = core_csr_io_bp_0_control_m;
    assign core__csr_io_bp_0_control_h = core_csr_io_bp_0_control_h;
    assign core__csr_io_bp_0_control_s = core_csr_io_bp_0_control_s;
    assign core__csr_io_bp_0_control_u = core_csr_io_bp_0_control_u;
    assign core__csr_io_bp_0_control_x = core_csr_io_bp_0_control_x;
    assign core__csr_io_bp_0_control_w = core_csr_io_bp_0_control_w;
    assign core__csr_io_bp_0_control_r = core_csr_io_bp_0_control_r;
    assign core__csr_io_bp_0_address = core_csr_io_bp_0_address;
    assign core__csr_io_bp_0_textra_mselect = core_csr_io_bp_0_textra_mselect;
    assign core__csr_io_bp_0_textra_pad2 = core_csr_io_bp_0_textra_pad2;
    assign core__csr_io_bp_0_textra_pad1 = core_csr_io_bp_0_textra_pad1;
    assign core__csr_io_bp_0_textra_sselect = core_csr_io_bp_0_textra_sselect;
    assign core_io_ptw_pmp_0_cfg_l = core_csr_io_pmp_0_cfg_l;
    assign core_io_ptw_pmp_0_cfg_res = core_csr_io_pmp_0_cfg_res;
    assign core_io_ptw_pmp_0_cfg_a = core_csr_io_pmp_0_cfg_a;
    assign core_io_ptw_pmp_0_cfg_x = core_csr_io_pmp_0_cfg_x;
    assign core_io_ptw_pmp_0_cfg_w = core_csr_io_pmp_0_cfg_w;
    assign core_io_ptw_pmp_0_cfg_r = core_csr_io_pmp_0_cfg_r;
    assign core_io_ptw_pmp_0_addr = core_csr_io_pmp_0_addr;
    assign core_io_ptw_pmp_0_mask = core_csr_io_pmp_0_mask;
    assign core_io_ptw_pmp_1_cfg_l = core_csr_io_pmp_1_cfg_l;
    assign core_io_ptw_pmp_1_cfg_res = core_csr_io_pmp_1_cfg_res;
    assign core_io_ptw_pmp_1_cfg_a = core_csr_io_pmp_1_cfg_a;
    assign core_io_ptw_pmp_1_cfg_x = core_csr_io_pmp_1_cfg_x;
    assign core_io_ptw_pmp_1_cfg_w = core_csr_io_pmp_1_cfg_w;
    assign core_io_ptw_pmp_1_cfg_r = core_csr_io_pmp_1_cfg_r;
    assign core_io_ptw_pmp_1_addr = core_csr_io_pmp_1_addr;
    assign core_io_ptw_pmp_1_mask = core_csr_io_pmp_1_mask;
    assign core_io_ptw_pmp_2_cfg_l = core_csr_io_pmp_2_cfg_l;
    assign core_io_ptw_pmp_2_cfg_res = core_csr_io_pmp_2_cfg_res;
    assign core_io_ptw_pmp_2_cfg_a = core_csr_io_pmp_2_cfg_a;
    assign core_io_ptw_pmp_2_cfg_x = core_csr_io_pmp_2_cfg_x;
    assign core_io_ptw_pmp_2_cfg_w = core_csr_io_pmp_2_cfg_w;
    assign core_io_ptw_pmp_2_cfg_r = core_csr_io_pmp_2_cfg_r;
    assign core_io_ptw_pmp_2_addr = core_csr_io_pmp_2_addr;
    assign core_io_ptw_pmp_2_mask = core_csr_io_pmp_2_mask;
    assign core_io_ptw_pmp_3_cfg_l = core_csr_io_pmp_3_cfg_l;
    assign core_io_ptw_pmp_3_cfg_res = core_csr_io_pmp_3_cfg_res;
    assign core_io_ptw_pmp_3_cfg_a = core_csr_io_pmp_3_cfg_a;
    assign core_io_ptw_pmp_3_cfg_x = core_csr_io_pmp_3_cfg_x;
    assign core_io_ptw_pmp_3_cfg_w = core_csr_io_pmp_3_cfg_w;
    assign core_io_ptw_pmp_3_cfg_r = core_csr_io_pmp_3_cfg_r;
    assign core_io_ptw_pmp_3_addr = core_csr_io_pmp_3_addr;
    assign core_io_ptw_pmp_3_mask = core_csr_io_pmp_3_mask;
    assign core_io_ptw_pmp_4_cfg_l = core_csr_io_pmp_4_cfg_l;
    assign core_io_ptw_pmp_4_cfg_res = core_csr_io_pmp_4_cfg_res;
    assign core_io_ptw_pmp_4_cfg_a = core_csr_io_pmp_4_cfg_a;
    assign core_io_ptw_pmp_4_cfg_x = core_csr_io_pmp_4_cfg_x;
    assign core_io_ptw_pmp_4_cfg_w = core_csr_io_pmp_4_cfg_w;
    assign core_io_ptw_pmp_4_cfg_r = core_csr_io_pmp_4_cfg_r;
    assign core_io_ptw_pmp_4_addr = core_csr_io_pmp_4_addr;
    assign core_io_ptw_pmp_4_mask = core_csr_io_pmp_4_mask;
    assign core_io_ptw_pmp_5_cfg_l = core_csr_io_pmp_5_cfg_l;
    assign core_io_ptw_pmp_5_cfg_res = core_csr_io_pmp_5_cfg_res;
    assign core_io_ptw_pmp_5_cfg_a = core_csr_io_pmp_5_cfg_a;
    assign core_io_ptw_pmp_5_cfg_x = core_csr_io_pmp_5_cfg_x;
    assign core_io_ptw_pmp_5_cfg_w = core_csr_io_pmp_5_cfg_w;
    assign core_io_ptw_pmp_5_cfg_r = core_csr_io_pmp_5_cfg_r;
    assign core_io_ptw_pmp_5_addr = core_csr_io_pmp_5_addr;
    assign core_io_ptw_pmp_5_mask = core_csr_io_pmp_5_mask;
    assign core_io_ptw_pmp_6_cfg_l = core_csr_io_pmp_6_cfg_l;
    assign core_io_ptw_pmp_6_cfg_res = core_csr_io_pmp_6_cfg_res;
    assign core_io_ptw_pmp_6_cfg_a = core_csr_io_pmp_6_cfg_a;
    assign core_io_ptw_pmp_6_cfg_x = core_csr_io_pmp_6_cfg_x;
    assign core_io_ptw_pmp_6_cfg_w = core_csr_io_pmp_6_cfg_w;
    assign core_io_ptw_pmp_6_cfg_r = core_csr_io_pmp_6_cfg_r;
    assign core_io_ptw_pmp_6_addr = core_csr_io_pmp_6_addr;
    assign core_io_ptw_pmp_6_mask = core_csr_io_pmp_6_mask;
    assign core_io_ptw_pmp_7_cfg_l = core_csr_io_pmp_7_cfg_l;
    assign core_io_ptw_pmp_7_cfg_res = core_csr_io_pmp_7_cfg_res;
    assign core_io_ptw_pmp_7_cfg_a = core_csr_io_pmp_7_cfg_a;
    assign core_io_ptw_pmp_7_cfg_x = core_csr_io_pmp_7_cfg_x;
    assign core_io_ptw_pmp_7_cfg_w = core_csr_io_pmp_7_cfg_w;
    assign core_io_ptw_pmp_7_cfg_r = core_csr_io_pmp_7_cfg_r;
    assign core_io_ptw_pmp_7_addr = core_csr_io_pmp_7_addr;
    assign core_io_ptw_pmp_7_mask = core_csr_io_pmp_7_mask;
    assign core__csr_io_inhibit_cycle = core_csr_io_inhibit_cycle;
    assign core_csr_io_inst_0 = core__GEN_4;
    assign core__csr_io_trace_0_valid = core_csr_io_trace_0_valid;
    assign core__csr_io_trace_0_iaddr = core_csr_io_trace_0_iaddr;
    assign core__csr_io_trace_0_insn = core_csr_io_trace_0_insn;
    assign core__csr_io_trace_0_priv = core_csr_io_trace_0_priv;
    assign core__csr_io_trace_0_exception = core_csr_io_trace_0_exception;
    assign core_io_trace_insns_0_interrupt = core_csr_io_trace_0_interrupt;
    assign core_io_trace_insns_0_cause = core_csr_io_trace_0_cause;
    assign core_io_trace_insns_0_tval = core_csr_io_trace_0_tval;
    assign core_io_ptw_customCSRs_csrs_0_ren = core_csr_io_customCSRs_0_ren;
    assign core_io_ptw_customCSRs_csrs_0_wen = core_csr_io_customCSRs_0_wen;
    assign core_io_ptw_customCSRs_csrs_0_wdata = core_csr_io_customCSRs_0_wdata;
    assign core__io_ptw_customCSRs_csrs_0_value_output = core_csr_io_customCSRs_0_value;
    assign core_csr_io_customCSRs_0_stall = core_io_ptw_customCSRs_csrs_0_stall;
    assign core_csr_io_customCSRs_0_set = core_io_ptw_customCSRs_csrs_0_set;
    assign core_csr_io_customCSRs_0_sdata = core_io_ptw_customCSRs_csrs_0_sdata;
    assign core_io_ptw_customCSRs_csrs_1_ren = core_csr_io_customCSRs_1_ren;
    assign core_io_ptw_customCSRs_csrs_1_wen = core_csr_io_customCSRs_1_wen;
    assign core_io_ptw_customCSRs_csrs_1_wdata = core_csr_io_customCSRs_1_wdata;
    assign core_io_ptw_customCSRs_csrs_1_value = core_csr_io_customCSRs_1_value;
    assign core_csr_io_customCSRs_1_stall = core_io_ptw_customCSRs_csrs_1_stall;
    assign core_csr_io_customCSRs_1_set = core_io_ptw_customCSRs_csrs_1_set;
    assign core_csr_io_customCSRs_1_sdata = core_io_ptw_customCSRs_csrs_1_sdata;
    assign core_io_ptw_customCSRs_csrs_2_ren = core_csr_io_customCSRs_2_ren;
    assign core_io_ptw_customCSRs_csrs_2_wen = core_csr_io_customCSRs_2_wen;
    assign core_io_ptw_customCSRs_csrs_2_wdata = core_csr_io_customCSRs_2_wdata;
    assign core_io_ptw_customCSRs_csrs_2_value = core_csr_io_customCSRs_2_value;
    assign core_csr_io_customCSRs_2_stall = core_io_ptw_customCSRs_csrs_2_stall;
    assign core_csr_io_customCSRs_2_set = core_io_ptw_customCSRs_csrs_2_set;
    assign core_csr_io_customCSRs_2_sdata = core_io_ptw_customCSRs_csrs_2_sdata;
    assign core_io_ptw_customCSRs_csrs_3_ren = core_csr_io_customCSRs_3_ren;
    assign core_io_ptw_customCSRs_csrs_3_wen = core_csr_io_customCSRs_3_wen;
    assign core_io_ptw_customCSRs_csrs_3_wdata = core_csr_io_customCSRs_3_wdata;
    assign core_io_ptw_customCSRs_csrs_3_value = core_csr_io_customCSRs_3_value;
    assign core_csr_io_customCSRs_3_stall = core_io_ptw_customCSRs_csrs_3_stall;
    assign core_csr_io_customCSRs_3_set = core_io_ptw_customCSRs_csrs_3_set;
    assign core_csr_io_customCSRs_3_sdata = core_io_ptw_customCSRs_csrs_3_sdata;
     
    wire core_coreMonitorBundle_excpt ; 
  assign  core_coreMonitorBundle_excpt = core__csr_io_trace_0_exception ; 
    wire[2:0] core_coreMonitorBundle_priv_mode ; 
  assign  core_coreMonitorBundle_priv_mode = core__csr_io_trace_0_priv ; 
    wire[31:0] core_coreMonitorBundle_inst ; 
  assign  core_coreMonitorBundle_inst = core__csr_io_trace_0_insn ; 
    wire[2:0] core_xrfWriteBundle_priv_mode ; 
  assign  core_xrfWriteBundle_priv_mode = core__csr_io_trace_0_priv ; 
    wire core_id_csr_en = core_id_ctrl_csr ==3'h6|(& core_id_ctrl_csr )| core_id_ctrl_csr ==3'h5; 
    wire core_id_system_insn = core_id_ctrl_csr ==3'h4; 
    wire core_id_csr_ren =( core_id_ctrl_csr ==3'h6|(& core_id_ctrl_csr ))& core__ibuf_io_inst_0_bits_inst_rs1 ==5'h0; 
    wire[2:0] core_id_csr = core_id_system_insn & core_id_ctrl_mem  ? 3'h0: core_id_csr_ren  ? 3'h2: core_id_ctrl_csr ; 
    wire core_id_csr_flush = core_id_system_insn | core_id_csr_en & core_id_csr_ren ==1'h0& core__csr_io_decode_0_write_flush ; 
    wire core_id_illegal_insn = core_id_ctrl_legal ==1'h0|( core_id_ctrl_mul | core_id_ctrl_div )& core__csr_io_status_isa [12]==1'h0| core_id_ctrl_amo & core__csr_io_status_isa [0]==1'h0| core_id_ctrl_fp &( core__csr_io_decode_0_fp_illegal | core_io_fpu_illegal_rm )| core_id_ctrl_dp & core__csr_io_status_isa [3]==1'h0| core__ibuf_io_inst_0_bits_rvc & core__csr_io_status_isa [2]==1'h0| core_id_ctrl_rocc & core__csr_io_decode_0_rocc_illegal | core_id_csr_en &( core__csr_io_decode_0_read_illegal | core_id_csr_ren ==1'h0& core__csr_io_decode_0_write_illegal )| core__ibuf_io_inst_0_bits_rvc ==1'h0& core_id_system_insn & core__csr_io_decode_0_system_illegal ; 
    wire core_id_virtual_insn = core_id_ctrl_legal &( core_id_csr_en &( core_id_csr_ren ==1'h0& core__csr_io_decode_0_write_illegal )==1'h0& core__csr_io_decode_0_virtual_access_illegal | core__ibuf_io_inst_0_bits_rvc ==1'h0& core_id_system_insn & core__csr_io_decode_0_virtual_system_illegal ); 
    wire core_id_amo_aq = core__ibuf_io_inst_0_bits_inst_bits [26]; 
    wire core_id_amo_rl = core__ibuf_io_inst_0_bits_inst_bits [25]; 
    wire[3:0] core_id_fence_pred = core__ibuf_io_inst_0_bits_inst_bits [27:24]; 
    wire[3:0] core_id_fence_succ = core__ibuf_io_inst_0_bits_inst_bits [23:20]; 
    wire core_id_fence_next = core_id_ctrl_fence | core_id_ctrl_amo & core_id_amo_aq ; 
    wire core__io_dmem_req_valid_output ; 
    wire core_id_mem_busy = core_io_dmem_ordered ==1'h0| core__io_dmem_req_valid_output ; 
    wire core__GEN_59 = core_id_mem_busy ==1'h0; 
    wire core__GEN_60 = core__GEN_59  ? 1'h0: core_id_reg_fence ; 
    wire core_id_do_fence = core_id_rocc_busy & core_id_ctrl_fence | core_id_mem_busy &( core_id_ctrl_amo & core_id_amo_rl | core_id_ctrl_fence_i | core_id_reg_fence &( core_id_ctrl_mem | core_id_ctrl_rocc ));  
    wire core_bpu_clock;
    wire core_bpu_reset;
    wire core_bpu_io_status_debug;
    wire core_bpu_io_status_cease;
    wire core_bpu_io_status_wfi;
    wire[31:0] core_bpu_io_status_isa;
    wire[1:0] core_bpu_io_status_dprv;
    wire core_bpu_io_status_dv;
    wire[1:0] core_bpu_io_status_prv;
    wire core_bpu_io_status_v;
    wire core_bpu_io_status_sd;
    wire[22:0] core_bpu_io_status_zero2;
    wire core_bpu_io_status_mpv;
    wire core_bpu_io_status_gva;
    wire core_bpu_io_status_mbe;
    wire core_bpu_io_status_sbe;
    wire[1:0] core_bpu_io_status_sxl;
    wire[1:0] core_bpu_io_status_uxl;
    wire core_bpu_io_status_sd_rv32;
    wire[7:0] core_bpu_io_status_zero1;
    wire core_bpu_io_status_tsr;
    wire core_bpu_io_status_tw;
    wire core_bpu_io_status_tvm;
    wire core_bpu_io_status_mxr;
    wire core_bpu_io_status_sum;
    wire core_bpu_io_status_mprv;
    wire[1:0] core_bpu_io_status_xs;
    wire[1:0] core_bpu_io_status_fs;
    wire[1:0] core_bpu_io_status_mpp;
    wire[1:0] core_bpu_io_status_vs;
    wire core_bpu_io_status_spp;
    wire core_bpu_io_status_mpie;
    wire core_bpu_io_status_ube;
    wire core_bpu_io_status_spie;
    wire core_bpu_io_status_upie;
    wire core_bpu_io_status_mie;
    wire core_bpu_io_status_hie;
    wire core_bpu_io_status_sie;
    wire core_bpu_io_status_uie;
    wire[3:0] core_bpu_io_bp_0_control_ttype;
    wire core_bpu_io_bp_0_control_dmode;
    wire[5:0] core_bpu_io_bp_0_control_maskmax;
    wire[39:0] core_bpu_io_bp_0_control_reserved;
    wire core_bpu_io_bp_0_control_action;
    wire core_bpu_io_bp_0_control_chain;
    wire[1:0] core_bpu_io_bp_0_control_zero;
    wire[1:0] core_bpu_io_bp_0_control_tmatch;
    wire core_bpu_io_bp_0_control_m;
    wire core_bpu_io_bp_0_control_h;
    wire core_bpu_io_bp_0_control_s;
    wire core_bpu_io_bp_0_control_u;
    wire core_bpu_io_bp_0_control_x;
    wire core_bpu_io_bp_0_control_w;
    wire core_bpu_io_bp_0_control_r;
    wire[32:0] core_bpu_io_bp_0_address;
    wire core_bpu_io_bp_0_textra_mselect;
    wire[47:0] core_bpu_io_bp_0_textra_pad2;
    wire core_bpu_io_bp_0_textra_pad1;
    wire core_bpu_io_bp_0_textra_sselect;
    wire[32:0] core_bpu_io_pc;
    wire[32:0] core_bpu_io_ea;
    wire core_bpu_io_xcpt_if;
    wire core_bpu_io_xcpt_ld;
    wire core_bpu_io_xcpt_st;
    wire core_bpu_io_debug_if;
    wire core_bpu_io_debug_ld;
    wire core_bpu_io_debug_st;
    wire core_bpu_io_bpwatch_0_valid_0;
    wire core_bpu_io_bpwatch_0_rvalid_0;
    wire core_bpu_io_bpwatch_0_wvalid_0;
    wire core_bpu_io_bpwatch_0_ivalid_0;
    wire[2:0] core_bpu_io_bpwatch_0_action;

    wire core_bpu_cx =1'h1; 
    wire[1:0] core_bpu_en_lo ={ core_bpu_io_bp_0_control_s , core_bpu_io_bp_0_control_u }; 
    wire[1:0] core_bpu_en_hi ={ core_bpu_io_bp_0_control_m , core_bpu_io_bp_0_control_h }; 
    wire[3:0] core_bpu__GEN ={ core_bpu_en_hi , core_bpu_en_lo }>> core_bpu_io_status_prv ; 
    wire core_bpu_en = core_bpu_io_status_debug ==1'h0& core_bpu__GEN [0]; 
    wire core_bpu__GEN_0 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_1 = core_bpu__GEN_0 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_r_lo ={ core_bpu__GEN_0 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_r_hi ={ core_bpu__GEN_1 & core_bpu_io_bp_0_address [2], core_bpu__GEN_1 }; 
    wire core_bpu__GEN_2 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_3 = core_bpu__GEN_2 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_r_lo_1 ={ core_bpu__GEN_2 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_r_hi_1 ={ core_bpu__GEN_3 & core_bpu_io_bp_0_address [2], core_bpu__GEN_3 }; 
    wire core_bpu_r = core_bpu_en & core_bpu_io_bp_0_control_r &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu_io_ea >= core_bpu_io_bp_0_address ^ core_bpu_io_bp_0_control_tmatch [0]:(~ core_bpu_io_ea |{29'h0,{ core_bpu_r_hi , core_bpu_r_lo }})==(~ core_bpu_io_bp_0_address |{29'h0,{ core_bpu_r_hi_1 , core_bpu_r_lo_1 }}))& core_bpu_cx ; 
    wire core_bpu__GEN_4 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_5 = core_bpu__GEN_4 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_w_lo ={ core_bpu__GEN_4 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_w_hi ={ core_bpu__GEN_5 & core_bpu_io_bp_0_address [2], core_bpu__GEN_5 }; 
    wire core_bpu__GEN_6 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_7 = core_bpu__GEN_6 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_w_lo_1 ={ core_bpu__GEN_6 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_w_hi_1 ={ core_bpu__GEN_7 & core_bpu_io_bp_0_address [2], core_bpu__GEN_7 }; 
    wire core_bpu_w = core_bpu_en & core_bpu_io_bp_0_control_w &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu_io_ea >= core_bpu_io_bp_0_address ^ core_bpu_io_bp_0_control_tmatch [0]:(~ core_bpu_io_ea |{29'h0,{ core_bpu_w_hi , core_bpu_w_lo }})==(~ core_bpu_io_bp_0_address |{29'h0,{ core_bpu_w_hi_1 , core_bpu_w_lo_1 }}))& core_bpu_cx ; 
    wire core_bpu__GEN_8 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_9 = core_bpu__GEN_8 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_x_lo ={ core_bpu__GEN_8 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_x_hi ={ core_bpu__GEN_9 & core_bpu_io_bp_0_address [2], core_bpu__GEN_9 }; 
    wire core_bpu__GEN_10 = core_bpu_io_bp_0_control_tmatch [0]& core_bpu_io_bp_0_address [0]; 
    wire core_bpu__GEN_11 = core_bpu__GEN_10 & core_bpu_io_bp_0_address [1]; 
    wire[1:0] core_bpu_x_lo_1 ={ core_bpu__GEN_10 , core_bpu_io_bp_0_control_tmatch [0]}; 
    wire[1:0] core_bpu_x_hi_1 ={ core_bpu__GEN_11 & core_bpu_io_bp_0_address [2], core_bpu__GEN_11 }; 
    wire core_bpu_x = core_bpu_en & core_bpu_io_bp_0_control_x &( core_bpu_io_bp_0_control_tmatch [1] ?  core_bpu_io_pc >= core_bpu_io_bp_0_address ^ core_bpu_io_bp_0_control_tmatch [0]:(~ core_bpu_io_pc |{29'h0,{ core_bpu_x_hi , core_bpu_x_lo }})==(~ core_bpu_io_bp_0_address |{29'h0,{ core_bpu_x_hi_1 , core_bpu_x_lo_1 }}))& core_bpu_cx ; 
    wire core_bpu_end_0 = core_bpu_io_bp_0_control_chain ==1'h0; 
    wire core_bpu__GEN_12 = core_bpu_end_0 & core_bpu_r ; 
    wire core_bpu__GEN_13 = core_bpu_end_0 & core_bpu_w ; 
    wire core_bpu__GEN_14 = core_bpu_end_0 & core_bpu_x ; 
  assign  core_bpu_io_xcpt_if = core_bpu__GEN_14  ?  core_bpu_io_bp_0_control_action ==1'h0:1'h0; 
  assign  core_bpu_io_xcpt_ld = core_bpu__GEN_12  ?  core_bpu_io_bp_0_control_action ==1'h0:1'h0; 
  assign  core_bpu_io_xcpt_st = core_bpu__GEN_13  ?  core_bpu_io_bp_0_control_action ==1'h0:1'h0; 
  assign  core_bpu_io_debug_if = core_bpu__GEN_14  ? (& core_bpu_io_bp_0_control_action ):1'h0; 
  assign  core_bpu_io_debug_ld = core_bpu__GEN_12  ? (& core_bpu_io_bp_0_control_action ):1'h0; 
  assign  core_bpu_io_debug_st = core_bpu__GEN_13  ? (& core_bpu_io_bp_0_control_action ):1'h0; 
  assign  core_bpu_io_bpwatch_0_valid_0 = core_bpu__GEN_14  ? 1'h1: core_bpu__GEN_13  ? 1'h1: core_bpu__GEN_12 ; 
  assign  core_bpu_io_bpwatch_0_rvalid_0 = core_bpu__GEN_12 ; 
  assign  core_bpu_io_bpwatch_0_wvalid_0 = core_bpu__GEN_13 ; 
  assign  core_bpu_io_bpwatch_0_ivalid_0 = core_bpu__GEN_14 ; 
  assign  core_bpu_io_bpwatch_0_action ={2'h0, core_bpu_io_bp_0_control_action };
    assign core_bpu_clock = core_clock;
    assign core_bpu_reset = core_reset;
    assign core_bpu_io_status_debug = core__csr_io_status_debug;
    assign core_bpu_io_status_cease = core__csr_io_status_cease;
    assign core_bpu_io_status_wfi = core__csr_io_status_wfi;
    assign core_bpu_io_status_isa = core__csr_io_status_isa;
    assign core_bpu_io_status_dprv = core__csr_io_status_dprv;
    assign core_bpu_io_status_dv = core__csr_io_status_dv;
    assign core_bpu_io_status_prv = core__csr_io_status_prv;
    assign core_bpu_io_status_v = core__csr_io_status_v;
    assign core_bpu_io_status_sd = core__csr_io_status_sd;
    assign core_bpu_io_status_zero2 = core__csr_io_status_zero2;
    assign core_bpu_io_status_mpv = core__csr_io_status_mpv;
    assign core_bpu_io_status_gva = core__csr_io_status_gva;
    assign core_bpu_io_status_mbe = core__csr_io_status_mbe;
    assign core_bpu_io_status_sbe = core__csr_io_status_sbe;
    assign core_bpu_io_status_sxl = core__csr_io_status_sxl;
    assign core_bpu_io_status_uxl = core__csr_io_status_uxl;
    assign core_bpu_io_status_sd_rv32 = core__csr_io_status_sd_rv32;
    assign core_bpu_io_status_zero1 = core__csr_io_status_zero1;
    assign core_bpu_io_status_tsr = core__csr_io_status_tsr;
    assign core_bpu_io_status_tw = core__csr_io_status_tw;
    assign core_bpu_io_status_tvm = core__csr_io_status_tvm;
    assign core_bpu_io_status_mxr = core__csr_io_status_mxr;
    assign core_bpu_io_status_sum = core__csr_io_status_sum;
    assign core_bpu_io_status_mprv = core__csr_io_status_mprv;
    assign core_bpu_io_status_xs = core__csr_io_status_xs;
    assign core_bpu_io_status_fs = core__csr_io_status_fs;
    assign core_bpu_io_status_mpp = core__csr_io_status_mpp;
    assign core_bpu_io_status_vs = core__csr_io_status_vs;
    assign core_bpu_io_status_spp = core__csr_io_status_spp;
    assign core_bpu_io_status_mpie = core__csr_io_status_mpie;
    assign core_bpu_io_status_ube = core__csr_io_status_ube;
    assign core_bpu_io_status_spie = core__csr_io_status_spie;
    assign core_bpu_io_status_upie = core__csr_io_status_upie;
    assign core_bpu_io_status_mie = core__csr_io_status_mie;
    assign core_bpu_io_status_hie = core__csr_io_status_hie;
    assign core_bpu_io_status_sie = core__csr_io_status_sie;
    assign core_bpu_io_status_uie = core__csr_io_status_uie;
    assign core_bpu_io_bp_0_control_ttype = core__csr_io_bp_0_control_ttype;
    assign core_bpu_io_bp_0_control_dmode = core__csr_io_bp_0_control_dmode;
    assign core_bpu_io_bp_0_control_maskmax = core__csr_io_bp_0_control_maskmax;
    assign core_bpu_io_bp_0_control_reserved = core__csr_io_bp_0_control_reserved;
    assign core_bpu_io_bp_0_control_action = core__csr_io_bp_0_control_action;
    assign core_bpu_io_bp_0_control_chain = core__csr_io_bp_0_control_chain;
    assign core_bpu_io_bp_0_control_zero = core__csr_io_bp_0_control_zero;
    assign core_bpu_io_bp_0_control_tmatch = core__csr_io_bp_0_control_tmatch;
    assign core_bpu_io_bp_0_control_m = core__csr_io_bp_0_control_m;
    assign core_bpu_io_bp_0_control_h = core__csr_io_bp_0_control_h;
    assign core_bpu_io_bp_0_control_s = core__csr_io_bp_0_control_s;
    assign core_bpu_io_bp_0_control_u = core__csr_io_bp_0_control_u;
    assign core_bpu_io_bp_0_control_x = core__csr_io_bp_0_control_x;
    assign core_bpu_io_bp_0_control_w = core__csr_io_bp_0_control_w;
    assign core_bpu_io_bp_0_control_r = core__csr_io_bp_0_control_r;
    assign core_bpu_io_bp_0_address = core__csr_io_bp_0_address;
    assign core_bpu_io_bp_0_textra_mselect = core__csr_io_bp_0_textra_mselect;
    assign core_bpu_io_bp_0_textra_pad2 = core__csr_io_bp_0_textra_pad2;
    assign core_bpu_io_bp_0_textra_pad1 = core__csr_io_bp_0_textra_pad1;
    assign core_bpu_io_bp_0_textra_sselect = core__csr_io_bp_0_textra_sselect;
    assign core_bpu_io_pc = core__ibuf_io_pc_32to0;
    assign core_bpu_io_ea = core__mem_reg_wdata_32to0;
    assign core__bpu_io_xcpt_if = core_bpu_io_xcpt_if;
    assign core__bpu_io_xcpt_ld = core_bpu_io_xcpt_ld;
    assign core__bpu_io_xcpt_st = core_bpu_io_xcpt_st;
    assign core__bpu_io_debug_if = core_bpu_io_debug_if;
    assign core__bpu_io_debug_ld = core_bpu_io_debug_ld;
    assign core__bpu_io_debug_st = core_bpu_io_debug_st;
    assign core__bpu_io_bpwatch_0_rvalid_0 = core_bpu_io_bpwatch_0_rvalid_0;
    assign core__bpu_io_bpwatch_0_wvalid_0 = core_bpu_io_bpwatch_0_wvalid_0;
    assign core__bpu_io_bpwatch_0_ivalid_0 = core_bpu_io_bpwatch_0_ivalid_0;
     
  assign  core__ibuf_io_pc_32to0 = core__ibuf_io_pc [32:0]; 
  assign  core__mem_reg_wdata_32to0 = core_mem_reg_wdata [32:0]; 
    wire core_id_xcpt = core__csr_io_interrupt | core__bpu_io_debug_if | core__bpu_io_xcpt_if | core__ibuf_io_inst_0_bits_xcpt0_pf_inst | core__ibuf_io_inst_0_bits_xcpt0_gf_inst | core__ibuf_io_inst_0_bits_xcpt0_ae_inst | core__ibuf_io_inst_0_bits_xcpt1_pf_inst | core__ibuf_io_inst_0_bits_xcpt1_gf_inst | core__ibuf_io_inst_0_bits_xcpt1_ae_inst | core_id_virtual_insn | core_id_illegal_insn ; 
    wire[63:0] core_id_cause = core__csr_io_interrupt  ?  core__csr_io_interrupt_cause :{59'h0, core__bpu_io_debug_if  ? 5'hE: core__bpu_io_xcpt_if  ? 5'h3: core__ibuf_io_inst_0_bits_xcpt0_pf_inst  ? 5'hC: core__ibuf_io_inst_0_bits_xcpt0_gf_inst  ? 5'h14: core__ibuf_io_inst_0_bits_xcpt0_ae_inst  ? 5'h1: core__ibuf_io_inst_0_bits_xcpt1_pf_inst  ? 5'hC: core__ibuf_io_inst_0_bits_xcpt1_gf_inst  ? 5'h14: core__ibuf_io_inst_0_bits_xcpt1_ae_inst  ? 5'h1: core_id_virtual_insn  ? 5'h16:5'h2}; 
    wire[4:0] core_ex_waddr = core_ex_reg_inst [11:7]; 
    wire[4:0] core_mem_waddr = core_mem_reg_inst [11:7]; 
    wire[4:0] core_wb_waddr = core_wb_reg_inst [11:7]; 
    wire[4:0] core_coreMonitorBundle_wrdst = core_wb_waddr ; 
    wire core__GEN_61 = core_ex_reg_valid & core_ex_ctrl_wxd ; 
    wire core__GEN_62 = core_mem_reg_valid & core_mem_ctrl_wxd & core_mem_ctrl_mem ==1'h0; 
    wire core__GEN_63 = core_mem_reg_valid & core_mem_ctrl_wxd ; 
    wire core_id_bypass_src_0_0 =5'h0== core_id_raddr1 &1'h1; 
    wire core_id_bypass_src_0_1 = core__GEN_61 & core_ex_waddr == core_id_raddr1 ; 
    wire core_id_bypass_src_0_2 = core__GEN_62 & core_mem_waddr == core_id_raddr1 ; 
    wire core_id_bypass_src_0_3 = core__GEN_63 & core_mem_waddr == core_id_raddr1 ; 
    wire core_id_bypass_src_1_0 =5'h0== core_id_raddr2 &1'h1; 
    wire core_id_bypass_src_1_1 = core__GEN_61 & core_ex_waddr == core_id_raddr2 ; 
    wire core_id_bypass_src_1_2 = core__GEN_62 & core_mem_waddr == core_id_raddr2 ; 
    wire core_id_bypass_src_1_3 = core__GEN_63 & core_mem_waddr == core_id_raddr2 ; 
    reg core_ex_reg_rs_bypass_0 ; 
    reg core_ex_reg_rs_bypass_1 ; reg[1:0] core_ex_reg_rs_lsb_0 ; reg[1:0] core_ex_reg_rs_lsb_1 ; reg[61:0] core_ex_reg_rs_msb_0 ; reg[61:0] core_ex_reg_rs_msb_1 ; 
    wire[63:0] core_ex_rs_0 = core_ex_reg_rs_bypass_0  ? ((& core_ex_reg_rs_lsb_0 ) ?  core_dcache_bypass_data : core_ex_reg_rs_lsb_0 ==2'h2 ?  core_wb_reg_wdata : core_ex_reg_rs_lsb_0 ==2'h1 ?  core_mem_reg_wdata :64'h0):{ core_ex_reg_rs_msb_0 , core_ex_reg_rs_lsb_0 }; 
    wire[63:0] core_ex_rs_1 = core_ex_reg_rs_bypass_1  ? ((& core_ex_reg_rs_lsb_1 ) ?  core_dcache_bypass_data : core_ex_reg_rs_lsb_1 ==2'h2 ?  core_wb_reg_wdata : core_ex_reg_rs_lsb_1 ==2'h1 ?  core_mem_reg_wdata :64'h0):{ core_ex_reg_rs_msb_1 , core_ex_reg_rs_lsb_1 }; 
    wire core_ex_imm_sign = core_ex_ctrl_sel_imm ==3'h5 ? 1'h0: core_ex_reg_inst [31]; 
    wire core_ex_imm_hi_hi_hi = core_ex_imm_sign ; 
    wire[10:0] core_ex_imm_b30_20 = core_ex_ctrl_sel_imm ==3'h2 ?  core_ex_reg_inst [30:20]:{{10{ core_ex_imm_sign }}, core_ex_imm_sign }; 
    wire[10:0] core_ex_imm_hi_hi_lo = core_ex_imm_b30_20 ; 
    wire[7:0] core_ex_imm_b19_12 = core_ex_ctrl_sel_imm !=3'h2& core_ex_ctrl_sel_imm !=3'h3 ? {{7{ core_ex_imm_sign }}, core_ex_imm_sign }: core_ex_reg_inst [19:12]; 
    wire[7:0] core_ex_imm_hi_lo_hi = core_ex_imm_b19_12 ; 
    wire core_ex_imm_b11 = core_ex_ctrl_sel_imm ==3'h2| core_ex_ctrl_sel_imm ==3'h5 ? 1'h0: core_ex_ctrl_sel_imm ==3'h3 ?  core_ex_reg_inst [20]: core_ex_ctrl_sel_imm ==3'h1 ?  core_ex_reg_inst [7]: core_ex_imm_sign ; 
    wire core_ex_imm_hi_lo_lo = core_ex_imm_b11 ; 
    wire[5:0] core_ex_imm_b10_5 = core_ex_ctrl_sel_imm ==3'h2| core_ex_ctrl_sel_imm ==3'h5 ? 6'h0: core_ex_reg_inst [30:25]; 
    wire[3:0] core_ex_imm_b4_1 = core_ex_ctrl_sel_imm ==3'h2 ? 4'h0: core_ex_ctrl_sel_imm ==3'h0| core_ex_ctrl_sel_imm ==3'h1 ?  core_ex_reg_inst [11:8]: core_ex_ctrl_sel_imm ==3'h5 ?  core_ex_reg_inst [19:16]: core_ex_reg_inst [24:21]; 
    wire core_ex_imm_b0 = core_ex_ctrl_sel_imm ==3'h0 ?  core_ex_reg_inst [7]: core_ex_ctrl_sel_imm ==3'h4 ?  core_ex_reg_inst [20]: core_ex_ctrl_sel_imm ==3'h5 ?  core_ex_reg_inst [15]:1'h0; 
    wire[9:0] core_ex_imm_lo_hi ={ core_ex_imm_b10_5 , core_ex_imm_b4_1 }; 
    wire[10:0] core_ex_imm_lo ={ core_ex_imm_lo_hi , core_ex_imm_b0 }; 
    wire[8:0] core_ex_imm_hi_lo ={ core_ex_imm_hi_lo_hi , core_ex_imm_hi_lo_lo }; 
    wire[11:0] core_ex_imm_hi_hi ={ core_ex_imm_hi_hi_hi , core_ex_imm_hi_hi_lo }; 
    wire[20:0] core_ex_imm_hi ={ core_ex_imm_hi_hi , core_ex_imm_hi_lo }; 
    wire[31:0] core_ex_imm ={ core_ex_imm_hi , core_ex_imm_lo }; 
    wire[63:0] core_ex_op1 =2'h2== core_ex_ctrl_sel_alu1  ? {{30{ core_ex_reg_pc [33]}}, core_ex_reg_pc }:2'h1== core_ex_ctrl_sel_alu1  ?  core_ex_rs_0 :64'h0; 
    wire[3:0] core__GEN_64 = core_ex_reg_rvc  ? 4'h2:4'h4; 
    wire[63:0] core_ex_op2 =2'h1== core_ex_ctrl_sel_alu2  ? {{60{ core__GEN_64 [3]}}, core__GEN_64 }:2'h3== core_ex_ctrl_sel_alu2  ? {{32{ core_ex_imm [31]}}, core_ex_imm }:2'h2== core_ex_ctrl_sel_alu2  ?  core_ex_rs_1 :64'h0;  
    wire core_alu_clock;
    wire core_alu_reset;
    wire core_alu_io_dw;
    wire[3:0] core_alu_io_fn;
    wire[63:0] core_alu_io_in2;
    wire[63:0] core_alu_io_in1;
    wire[63:0] core_alu_io_out;
    wire[63:0] core_alu_io_adder_out;
    wire core_alu_io_cmp_out;

    wire[63:0] core_alu_in2_inv = core_alu_io_fn [3] ? ~ core_alu_io_in2 : core_alu_io_in2 ; 
    wire[63:0] core_alu_in1_xor_in2 = core_alu_io_in1 ^ core_alu_in2_inv ; 
    wire[64:0] core_alu__GEN ={1'h0, core_alu_io_in1 }+{1'h0, core_alu_in2_inv }; 
    wire[64:0] core_alu__GEN_0 ={1'h0, core_alu__GEN [63:0]}+{64'h0, core_alu_io_fn [3]}; 
    wire[63:0] core_alu__io_adder_out_output = core_alu__GEN_0 [63:0]; 
    wire core_alu_slt = core_alu_io_in1 [63]== core_alu_io_in2 [63] ?  core_alu__io_adder_out_output [63]: core_alu_io_fn [1] ?  core_alu_io_in2 [63]: core_alu_io_in1 [63]; 
    wire[31:0] core_alu_shin_hi_32 = core_alu_io_fn [3]& core_alu_io_in1 [31] ? 32'hFFFFFFFF:32'h0; 
    wire[31:0] core_alu_shin_hi =(& core_alu_io_dw ) ?  core_alu_io_in1 [63:32]: core_alu_shin_hi_32 ; 
    wire[5:0] core_alu_shamt ={ core_alu_io_in2 [5]&(& core_alu_io_dw ), core_alu_io_in2 [4:0]}; 
    wire[63:0] core_alu_shin_r ={ core_alu_shin_hi , core_alu_io_in1 [31:0]}; 
    wire[63:0] core_alu__GEN_1 ={32'h0, core_alu_shin_r [63:32]}&64'hFFFFFFFF|{ core_alu_shin_r [31:0],32'h0}&64'hFFFFFFFF00000000; 
    wire[63:0] core_alu__GEN_2 ={16'h0, core_alu__GEN_1 [63:16]}&64'hFFFF0000FFFF|{ core_alu__GEN_1 [47:0],16'h0}&64'hFFFF0000FFFF0000; 
    wire[63:0] core_alu__GEN_3 ={8'h0, core_alu__GEN_2 [63:8]}&64'hFF00FF00FF00FF|{ core_alu__GEN_2 [55:0],8'h0}&64'hFF00FF00FF00FF00; 
    wire[63:0] core_alu__GEN_4 ={4'h0, core_alu__GEN_3 [63:4]}&64'hF0F0F0F0F0F0F0F|{ core_alu__GEN_3 [59:0],4'h0}&64'hF0F0F0F0F0F0F0F0; 
    wire[63:0] core_alu__GEN_5 ={2'h0, core_alu__GEN_4 [63:2]}&64'h3333333333333333|{ core_alu__GEN_4 [61:0],2'h0}&64'hCCCCCCCCCCCCCCCC; 
    wire[63:0] core_alu_shin = core_alu_io_fn ==4'h5| core_alu_io_fn ==4'hB ?  core_alu_shin_r :{1'h0, core_alu__GEN_5 [63:1]}&64'h5555555555555555|{ core_alu__GEN_5 [62:0],1'h0}&64'hAAAAAAAAAAAAAAAA; 
    wire[64:0] core_alu__GEN_6 =$signed($signed({ core_alu_io_fn [3]& core_alu_shin [63], core_alu_shin })>>> core_alu_shamt ); 
    wire[63:0] core_alu_shout_r = core_alu__GEN_6 [63:0]; 
    wire[63:0] core_alu__GEN_7 ={32'h0, core_alu_shout_r [63:32]}&64'hFFFFFFFF|{ core_alu_shout_r [31:0],32'h0}&64'hFFFFFFFF00000000; 
    wire[63:0] core_alu__GEN_8 ={16'h0, core_alu__GEN_7 [63:16]}&64'hFFFF0000FFFF|{ core_alu__GEN_7 [47:0],16'h0}&64'hFFFF0000FFFF0000; 
    wire[63:0] core_alu__GEN_9 ={8'h0, core_alu__GEN_8 [63:8]}&64'hFF00FF00FF00FF|{ core_alu__GEN_8 [55:0],8'h0}&64'hFF00FF00FF00FF00; 
    wire[63:0] core_alu__GEN_10 ={4'h0, core_alu__GEN_9 [63:4]}&64'hF0F0F0F0F0F0F0F|{ core_alu__GEN_9 [59:0],4'h0}&64'hF0F0F0F0F0F0F0F0; 
    wire[63:0] core_alu__GEN_11 ={2'h0, core_alu__GEN_10 [63:2]}&64'h3333333333333333|{ core_alu__GEN_10 [61:0],2'h0}&64'hCCCCCCCCCCCCCCCC; 
    wire[63:0] core_alu_shout_l ={1'h0, core_alu__GEN_11 [63:1]}&64'h5555555555555555|{ core_alu__GEN_11 [62:0],1'h0}&64'hAAAAAAAAAAAAAAAA; 
    wire[63:0] core_alu_shout =( core_alu_io_fn ==4'h5| core_alu_io_fn ==4'hB ?  core_alu_shout_r :64'h0)|( core_alu_io_fn ==4'h1 ?  core_alu_shout_l :64'h0); 
    wire core_alu_in2_not_zero =| core_alu_io_in2 ; 
    wire[63:0] core_alu_logic_0 =( core_alu_io_fn ==4'h4| core_alu_io_fn ==4'h6 ?  core_alu_in1_xor_in2 :64'h0)|( core_alu_io_fn ==4'h6| core_alu_io_fn ==4'h7 ?  core_alu_io_in1 & core_alu_io_in2 :64'h0); 
    wire[63:0] core_alu_shift_logic ={63'h0, core_alu_io_fn >=4'hC& core_alu_slt }| core_alu_logic_0 | core_alu_shout ; 
    wire[63:0] core_alu_out = core_alu_io_fn ==4'h0| core_alu_io_fn ==4'hA ?  core_alu__io_adder_out_output : core_alu_shift_logic ; 
  assign  core_alu_io_out = core_alu_io_dw ==1'h0 ? { core_alu_out [31] ? 32'hFFFFFFFF:32'h0, core_alu_out [31:0]}: core_alu_out ; 
  assign  core_alu_io_adder_out = core_alu__io_adder_out_output ; 
  assign  core_alu_io_cmp_out = core_alu_io_fn [0]^( core_alu_io_fn [3]==1'h0 ?  core_alu_in1_xor_in2 ==64'h0: core_alu_slt );
    assign core_alu_clock = core_clock;
    assign core_alu_reset = core_reset;
    assign core_alu_io_dw = core_ex_ctrl_alu_dw;
    assign core_alu_io_fn = core_ex_ctrl_alu_fn;
    assign core_alu_io_in2 = core_ex_op2;
    assign core_alu_io_in1 = core_ex_op1;
    assign core__alu_io_out = core_alu_io_out;
    assign core__alu_io_adder_out = core_alu_io_adder_out;
    assign core__alu_io_cmp_out = core_alu_io_cmp_out;
      
    wire core_div_clock;
    wire core_div_reset;
    wire core_div_io_req_ready;
    wire core_div_io_req_valid;
    wire[3:0] core_div_io_req_bits_fn;
    wire core_div_io_req_bits_dw;
    wire[63:0] core_div_io_req_bits_in1;
    wire[63:0] core_div_io_req_bits_in2;
    wire[4:0] core_div_io_req_bits_tag;
    wire core_div_io_kill;
    wire core_div_io_resp_ready;
    wire core_div_io_resp_valid;
    wire[63:0] core_div_io_resp_bits_data;
    wire[4:0] core_div_io_resp_bits_tag;

    wire core_div_eOut =1'h0; reg[2:0] core_div_state ; reg[3:0] core_div_req_fn ; 
    reg core_div_req_dw ; reg[63:0] core_div_req_in1 ; reg[63:0] core_div_req_in2 ; reg[4:0] core_div_req_tag ; reg[6:0] core_div_count ; 
    reg core_div_neg_out ; 
    reg core_div_isHi ; 
    reg core_div_resHi ; reg[64:0] core_div_divisor ; 
    wire[64:0] core_div_mpcand = core_div_divisor ; reg[129:0] core_div_remainder ; 
    wire[2:0] core_div_decoded_plaInput ; 
    wire[2:0] core_div_decoded_invInputs =~ core_div_decoded_plaInput ; 
    wire[3:0] core_div_decoded_invMatrixOutputs ; 
    wire core_div_decoded_andMatrixInput_0 = core_div_decoded_invInputs [0]; 
    wire core_div_decoded_andMatrixInput_0_1 = core_div_decoded_invInputs [2]; 
    wire core_div_decoded_andMatrixInput_0_2 = core_div_decoded_invInputs [1]; 
    wire core_div_decoded_andMatrixInput_1 = core_div_decoded_invInputs [2]; 
    wire core_div__GEN =&{ core_div_decoded_andMatrixInput_0_2 , core_div_decoded_andMatrixInput_1 }; 
    wire core_div_decoded_andMatrixInput_0_3 = core_div_decoded_plaInput [0]; 
    wire core_div_decoded_andMatrixInput_1_1 = core_div_decoded_invInputs [2]; 
    wire core_div_decoded_andMatrixInput_0_4 = core_div_decoded_plaInput [1]; 
    wire core_div_decoded_andMatrixInput_0_5 = core_div_decoded_invInputs [0]; 
    wire core_div_decoded_andMatrixInput_1_2 = core_div_decoded_plaInput [2]; 
    wire[1:0] core_div_decoded_orMatrixOutputs_lo ={|{& core_div_decoded_andMatrixInput_0 , core_div__GEN },|{ core_div__GEN ,&{ core_div_decoded_andMatrixInput_0_5 , core_div_decoded_andMatrixInput_1_2 }}}; 
    wire[1:0] core_div_decoded_orMatrixOutputs_hi ={|(& core_div_decoded_andMatrixInput_0_1 ),|{&{ core_div_decoded_andMatrixInput_0_3 , core_div_decoded_andMatrixInput_1_1 },& core_div_decoded_andMatrixInput_0_4 }}; 
    wire[3:0] core_div_decoded_orMatrixOutputs ={ core_div_decoded_orMatrixOutputs_hi , core_div_decoded_orMatrixOutputs_lo }; 
    wire[1:0] core_div_decoded_invMatrixOutputs_lo ={ core_div_decoded_orMatrixOutputs [1], core_div_decoded_orMatrixOutputs [0]}; 
    wire[1:0] core_div_decoded_invMatrixOutputs_hi ={ core_div_decoded_orMatrixOutputs [3], core_div_decoded_orMatrixOutputs [2]}; 
  assign  core_div_decoded_invMatrixOutputs ={ core_div_decoded_invMatrixOutputs_hi , core_div_decoded_invMatrixOutputs_lo }; 
    wire[3:0] core_div_decoded = core_div_decoded_invMatrixOutputs ; 
  assign  core_div_decoded_plaInput = core_div_io_req_bits_fn [2:0]; 
    wire core_div_cmdMul = core_div_decoded [3]; 
    wire core_div_cmdHi = core_div_decoded [2]; 
    wire core_div_lhsSigned = core_div_decoded [1]; 
    wire core_div_rhsSigned = core_div_decoded [0]; 
    wire core_div__GEN_0 = core_div_io_req_bits_dw ==1'h0&1'h1; 
    wire core_div_lhs_sign = core_div_lhsSigned &( core_div__GEN_0  ?  core_div_io_req_bits_in1 [31]: core_div_io_req_bits_in1 [63]); 
    wire[31:0] core_div_hi = core_div__GEN_0  ? ( core_div_lhs_sign  ? 32'hFFFFFFFF:32'h0): core_div_io_req_bits_in1 [63:32]; 
    wire[63:0] core_div_lhs_in ={ core_div_hi , core_div_io_req_bits_in1 [31:0]}; 
    wire core_div__GEN_1 = core_div_io_req_bits_dw ==1'h0&1'h1; 
    wire core_div_rhs_sign = core_div_rhsSigned &( core_div__GEN_1  ?  core_div_io_req_bits_in2 [31]: core_div_io_req_bits_in2 [63]); 
    wire[31:0] core_div_hi_1 = core_div__GEN_1  ? ( core_div_rhs_sign  ? 32'hFFFFFFFF:32'h0): core_div_io_req_bits_in2 [63:32]; 
    wire[63:0] core_div_rhs_in ={ core_div_hi_1 , core_div_io_req_bits_in2 [31:0]}; 
    wire[65:0] core_div__GEN_2 ={1'h0, core_div_remainder [128:64]}-{1'h0, core_div_divisor }; 
    wire[64:0] core_div_subtractor = core_div__GEN_2 [64:0]; 
    wire[63:0] core_div_result = core_div_resHi  ?  core_div_remainder [128:65]: core_div_remainder [63:0]; 
    wire[64:0] core_div__GEN_3 =65'h0-{1'h0, core_div_result }; 
    wire[63:0] core_div_negated_remainder = core_div__GEN_3 [63:0]; 
    wire core_div__GEN_4 = core_div_state ==3'h1; 
    wire[129:0] core_div__GEN_5 ={66'h0, core_div_negated_remainder }; 
    wire core_div__GEN_6 = core_div_state ==3'h5; 
    wire[129:0] core_div__GEN_7 ={66'h0, core_div_negated_remainder }; 
    wire[2:0] core_div__GEN_8 = core_div__GEN_6  ? 3'h7: core_div__GEN_4  ? 3'h3: core_div_state ; 
    wire core_div__GEN_9 = core_div__GEN_6  ? 1'h0: core_div_resHi ; 
    wire core_div__GEN_10 = core_div_state ==3'h2; 
    wire[128:0] core_div_mulReg ={ core_div_remainder [129:65], core_div_remainder [63:0]}; 
    wire core_div_mplierSign = core_div_remainder [64]; 
    wire[63:0] core_div_mplier = core_div_mulReg [63:0]; 
    wire[64:0] core_div_accum = core_div_mulReg [128:64]; 
    wire[1:0] core_div__GEN_11 ={ core_div_mplierSign , core_div_mplier [0]}; 
    wire[66:0] core_div__GEN_12 ={{65{ core_div__GEN_11 [1]}}, core_div__GEN_11 }*{{2{ core_div_mpcand [64]}}, core_div_mpcand }; 
    wire[67:0] core_div__GEN_13 ={ core_div__GEN_12 [66], core_div__GEN_12 }+{{3{ core_div_accum [64]}}, core_div_accum }; 
    wire[66:0] core_div_prod = core_div__GEN_13 [66:0]; 
    wire[66:0] core_div_nextMulReg_hi = core_div_prod ; 
    wire[129:0] core_div_nextMulReg ={ core_div_nextMulReg_hi , core_div_mplier [63:1]}; 
    wire core_div_nextMplierSign = core_div_count ==7'h3E& core_div_neg_out ; 
    wire[7:0] core_div__GEN_14 ={1'h0, core_div_count }*8'h1; 
    wire[64:0] core_div__GEN_15 =$signed(65'sh10000000000000000>>> core_div__GEN_14 [5:0]); 
    wire[63:0] core_div_eOutMask = core_div__GEN_15 [63:0]; 
    wire[8:0] core_div__GEN_16 =9'h40-{1'h0,{1'h0, core_div_count }*8'h1}; 
    wire[7:0] core_div__GEN_17 = core_div__GEN_16 [7:0]; 
    wire[128:0] core_div_eOutRes = core_div_mulReg >> core_div__GEN_17 [5:0]; 
    wire[129:0] core_div__GEN_18 = core_div_eOut  ? {1'h0, core_div_eOutRes }: core_div_nextMulReg ; 
    wire[128:0] core_div_nextMulReg1 ={ core_div_nextMulReg [128:64], core_div__GEN_18 [63:0]}; 
    wire[65:0] core_div_remainder_hi ={ core_div_nextMulReg1 [128:64], core_div_nextMplierSign }; 
    wire[129:0] core_div__GEN_19 ={ core_div_remainder_hi , core_div_nextMulReg1 [63:0]}; 
    wire[7:0] core_div__GEN_20 ={1'h0, core_div_count }+8'h1; 
    wire core_div__GEN_21 = core_div_eOut | core_div_count ==7'h3F; 
    wire[2:0] core_div__GEN_22 = core_div__GEN_10  ? ( core_div__GEN_21  ? 3'h6: core_div__GEN_8 ): core_div__GEN_8 ; 
    wire core_div__GEN_23 = core_div__GEN_10  ? ( core_div__GEN_21  ?  core_div_isHi : core_div__GEN_9 ): core_div__GEN_9 ; 
    wire core_div__GEN_24 = core_div_state ==3'h3; 
    wire core_div_unrolls_less = core_div_subtractor [64]; 
    wire[127:0] core_div_unrolls_hi ={ core_div_unrolls_less  ?  core_div_remainder [127:64]: core_div_subtractor [63:0], core_div_remainder [63:0]}; 
    wire[128:0] core_div_unrolls_0 ={ core_div_unrolls_hi , core_div_unrolls_less ==1'h0}; 
    wire[129:0] core_div__GEN_25 ={1'h0, core_div_unrolls_0 }; 
    wire core_div__GEN_26 = core_div_count ==7'h40; 
    wire[2:0] core_div__GEN_27 = core_div_neg_out  ? 3'h5:3'h7; 
    wire[7:0] core_div__GEN_28 ={1'h0, core_div_count }+8'h1; 
    wire core_div_divby0 = core_div_count ==7'h0& core_div_subtractor [64]==1'h0; 
    wire core_div__GEN_29 = core_div_divby0 & core_div_isHi ==1'h0; 
    wire core_div__io_resp_valid_output ; 
    wire core_div__GEN_30 = core_div_io_resp_ready & core_div__io_resp_valid_output | core_div_io_kill ; 
    wire core_div__io_req_ready_output ; 
    wire core_div__GEN_31 = core_div__io_req_ready_output & core_div_io_req_valid ; 
    wire[2:0] core_div__GEN_32 = core_div_cmdMul  ? 3'h2: core_div_lhs_sign | core_div_rhs_sign  ? 3'h1:3'h3; 
    wire[6:0] core_div__GEN_33 ={1'h0, core_div_cmdMul & core_div_io_req_bits_dw ==1'h0&1'h1 ? 6'h20:6'h0}; 
    wire core_div__GEN_34 = core_div_cmdHi  ?  core_div_lhs_sign : core_div_lhs_sign != core_div_rhs_sign ; 
    wire[64:0] core_div__GEN_35 ={ core_div_rhs_sign , core_div_rhs_in }; 
    wire[129:0] core_div__GEN_36 ={66'h0, core_div_lhs_in }; 
    wire core_div_outMul =( core_div_state &3'h1)==3'h0; 
    wire[31:0] core_div_loOut = core_div_req_dw ==1'h0&1'h1&1'h1& core_div_outMul  ?  core_div_result [63:32]: core_div_result [31:0]; 
    wire[31:0] core_div_hiOut = core_div_req_dw ==1'h0&1'h1 ? ( core_div_loOut [31] ? 32'hFFFFFFFF:32'h0): core_div_result [63:32]; 
  assign  core_div__io_resp_valid_output = core_div_state ==3'h6|(& core_div_state ); 
  assign  core_div__io_req_ready_output = core_div_state ==3'h0; 
  always @( posedge  core_div_clock )
         begin 
             if ( core_div_reset ) 
                 core_div_state  <=3'h0;
              else 
                 if ( core_div__GEN_31 ) 
                     core_div_state  <= core_div__GEN_32 ;
                  else 
                     if ( core_div__GEN_30 ) 
                         core_div_state  <=3'h0;
                      else 
                         if ( core_div__GEN_24 )
                             begin 
                                 if ( core_div__GEN_26 ) 
                                     core_div_state  <= core_div__GEN_27 ;
                                  else 
                                     if ( core_div__GEN_10 )
                                         begin 
                                             if ( core_div__GEN_21 ) 
                                                 core_div_state  <=3'h6;
                                              else 
                                                 if ( core_div__GEN_6 ) 
                                                     core_div_state  <=3'h7;
                                                  else 
                                                     if ( core_div__GEN_4 ) 
                                                         core_div_state  <=3'h3;
                                                      else 
                                                         begin 
                                                         end 
                                         end 
                                      else 
                                         if ( core_div__GEN_6 ) 
                                             core_div_state  <=3'h7;
                                          else 
                                             if ( core_div__GEN_4 ) 
                                                 core_div_state  <=3'h3;
                                              else 
                                                 begin 
                                                 end 
                             end 
                          else 
                             if ( core_div__GEN_10 )
                                 begin 
                                     if ( core_div__GEN_21 ) 
                                         core_div_state  <=3'h6;
                                      else 
                                         if ( core_div__GEN_6 ) 
                                             core_div_state  <=3'h7;
                                          else 
                                             if ( core_div__GEN_4 ) 
                                                 core_div_state  <=3'h3;
                                              else 
                                                 begin 
                                                 end 
                                 end 
                              else 
                                 if ( core_div__GEN_6 ) 
                                     core_div_state  <=3'h7;
                                  else 
                                     if ( core_div__GEN_4 ) 
                                         core_div_state  <=3'h3;
                                      else 
                                         begin 
                                         end 
         end
  always @( posedge  core_div_clock )
         begin 
             if ( core_div__GEN_31 )
                 begin  
                     core_div_req_fn  <= core_div_io_req_bits_fn ; 
                     core_div_req_dw  <= core_div_io_req_bits_dw ; 
                     core_div_req_in1  <= core_div_io_req_bits_in1 ; 
                     core_div_req_in2  <= core_div_io_req_bits_in2 ; 
                     core_div_req_tag  <= core_div_io_req_bits_tag ; 
                     core_div_count  <= core_div__GEN_33 ; 
                     core_div_neg_out  <= core_div__GEN_34 ; 
                     core_div_isHi  <= core_div_cmdHi ; 
                     core_div_resHi  <=1'h0; 
                     core_div_divisor  <= core_div__GEN_35 ; 
                     core_div_remainder  <= core_div__GEN_36 ;
                 end 
              else 
                 begin 
                     if ( core_div__GEN_24 )
                         begin  
                             core_div_count  <= core_div__GEN_28 [6:0];
                             if ( core_div__GEN_29 ) 
                                 core_div_neg_out  <=1'h0;
                              else 
                                 begin 
                                 end 
                             if ( core_div__GEN_26 ) 
                                 core_div_resHi  <= core_div_isHi ;
                              else 
                                 if ( core_div__GEN_10 )
                                     begin 
                                         if ( core_div__GEN_21 ) 
                                             core_div_resHi  <= core_div_isHi ;
                                          else 
                                             if ( core_div__GEN_6 ) 
                                                 core_div_resHi  <=1'h0;
                                              else 
                                                 begin 
                                                 end 
                                     end 
                                  else 
                                     if ( core_div__GEN_6 ) 
                                         core_div_resHi  <=1'h0;
                                      else 
                                         begin 
                                         end  
                             core_div_remainder  <= core_div__GEN_25 ;
                         end 
                      else 
                         if ( core_div__GEN_10 )
                             begin  
                                 core_div_count  <= core_div__GEN_20 [6:0];
                                 if ( core_div__GEN_21 ) 
                                     core_div_resHi  <= core_div_isHi ;
                                  else 
                                     if ( core_div__GEN_6 ) 
                                         core_div_resHi  <=1'h0;
                                      else 
                                         begin 
                                         end  
                                 core_div_remainder  <= core_div__GEN_19 ;
                             end 
                          else 
                             if ( core_div__GEN_6 )
                                 begin  
                                     core_div_resHi  <=1'h0; 
                                     core_div_remainder  <= core_div__GEN_7 ;
                                 end 
                              else 
                                 if ( core_div__GEN_4 )
                                     begin 
                                         if ( core_div_remainder [63]) 
                                             core_div_remainder  <= core_div__GEN_5 ;
                                          else 
                                             begin 
                                             end 
                                     end 
                                  else 
                                     begin 
                                     end 
                     if ( core_div__GEN_4 )
                         begin 
                             if ( core_div_divisor [63]) 
                                 core_div_divisor  <= core_div_subtractor ;
                              else 
                                 begin 
                                 end 
                         end 
                      else 
                         begin 
                         end 
                 end 
         end
  assign  core_div_io_req_ready = core_div__io_req_ready_output ; 
  assign  core_div_io_resp_valid = core_div__io_resp_valid_output ; 
  assign  core_div_io_resp_bits_data ={ core_div_hiOut , core_div_loOut }; 
  assign  core_div_io_resp_bits_tag = core_div_req_tag ;
    assign core_div_clock = core_clock;
    assign core_div_reset = core_reset;
    assign core__div_io_req_ready = core_div_io_req_ready;
    assign core_div_io_req_valid = core__GEN_9;
    assign core_div_io_req_bits_fn = core_ex_ctrl_alu_fn;
    assign core_div_io_req_bits_dw = core_ex_ctrl_alu_dw;
    assign core_div_io_req_bits_in1 = core_ex_rs_0;
    assign core_div_io_req_bits_in2 = core_ex_rs_1;
    assign core_div_io_req_bits_tag = core_ex_waddr;
    assign core_div_io_kill = core__GEN_8;
    assign core_div_io_resp_ready = core__GEN_7;
    assign core__div_io_resp_valid = core_div_io_resp_valid;
    assign core_ll_wdata = core_div_io_resp_bits_data;
    assign core__div_io_resp_bits_tag = core_div_io_resp_bits_tag;
     
  assign  core__GEN_9 = core_ex_reg_valid & core_ex_ctrl_div ; 
    wire core_ctrl_killd ; 
    wire core__GEN_65 = core_ctrl_killd ==1'h0; 
    wire core__GEN_66 = core_id_ctrl_fence & core_id_fence_succ ==4'h0; 
    wire core__GEN_67 = core__GEN_65 & core_id_xcpt ; 
    wire[3:0] core__GEN_68 = core_id_xcpt  ? 4'h0: core_id_ctrl_alu_fn ; 
    wire core__GEN_69 = core_id_xcpt  ? 1'h1: core_id_ctrl_alu_dw ; 
    wire[1:0] core_hi ={ core__ibuf_io_inst_0_bits_xcpt1_pf_inst , core__ibuf_io_inst_0_bits_xcpt1_gf_inst }; 
    wire core__GEN_70 =|{ core_hi , core__ibuf_io_inst_0_bits_xcpt1_ae_inst }; 
    wire core__GEN_71 = core_id_xcpt  ? ( core__GEN_70  ? 1'h1: core__ibuf_io_inst_0_bits_rvc ): core__ibuf_io_inst_0_bits_rvc ; 
    wire[1:0] core_hi_1 ={ core__ibuf_io_inst_0_bits_xcpt0_pf_inst , core__ibuf_io_inst_0_bits_xcpt0_gf_inst }; 
    wire core__GEN_72 = core__bpu_io_xcpt_if |(|{ core_hi_1 , core__ibuf_io_inst_0_bits_xcpt0_ae_inst }); 
    wire[1:0] core__GEN_73 = core_id_xcpt  ? ( core__GEN_72  ? 2'h2: core__GEN_70  ? 2'h2:2'h1): core_id_ctrl_sel_alu1 ; 
    wire[1:0] core__GEN_74 = core_id_xcpt  ? ( core__GEN_72  ? 2'h0: core__GEN_70  ? 2'h1:2'h0): core_id_ctrl_sel_alu2 ; 
    wire core__GEN_75 = core_id_ctrl_fence_i | core_id_csr_flush ; 
    wire core_id_load_use ; 
    wire core__GEN_76 = core_id_ctrl_mem_cmd ==5'h14| core_id_ctrl_mem_cmd ==5'h15| core_id_ctrl_mem_cmd ==5'h16| core_id_ctrl_mem_cmd ==5'h5; 
    wire[1:0] core__GEN_77 = core__GEN_76  ? {| core_id_raddr2 ,| core_id_raddr1 }: core__ibuf_io_inst_0_bits_inst_bits [13:12]; 
    wire core__GEN_78 = core_id_ctrl_mem_cmd ==5'h14& core__csr_io_status_v ; 
    wire[4:0] core__GEN_79 = core__GEN_78  ? 5'h15: core_id_ctrl_mem_cmd ; 
    wire core_do_bypass = core_id_bypass_src_0_0 | core_id_bypass_src_0_1 | core_id_bypass_src_0_2 | core_id_bypass_src_0_3 ; 
    wire[1:0] core_bypass_src = core_id_bypass_src_0_0  ? 2'h0: core_id_bypass_src_0_1  ? 2'h1: core_id_bypass_src_0_2  ? 2'h2:2'h3; 
    wire core__GEN_80 = core_id_ctrl_rxs1 & core_do_bypass ==1'h0; 
    wire[63:0] core_id_rs_0 ; 
    wire core_do_bypass_1 = core_id_bypass_src_1_0 | core_id_bypass_src_1_1 | core_id_bypass_src_1_2 | core_id_bypass_src_1_3 ; 
    wire[1:0] core_bypass_src_1 = core_id_bypass_src_1_0  ? 2'h0: core_id_bypass_src_1_1  ? 2'h1: core_id_bypass_src_1_2  ? 2'h2:2'h3; 
    wire core__GEN_81 = core_id_ctrl_rxs2 & core_do_bypass_1 ==1'h0; 
    wire[63:0] core_id_rs_1 ; 
    wire[1:0] core__GEN_82 = core__GEN_81  ?  core_id_rs_1 [1:0]: core_bypass_src_1 ; 
    wire core__GEN_83 = core_id_illegal_insn | core_id_virtual_insn ; 
    wire[31:0] core_inst = core__ibuf_io_inst_0_bits_rvc  ? {16'h0, core__ibuf_io_inst_0_bits_raw [15:0]}: core__ibuf_io_inst_0_bits_raw ; 
    wire core__GEN_84 = core__GEN_83  ? 1'h0: core_do_bypass ; 
    wire[1:0] core__GEN_85 = core__GEN_83  ?  core_inst [1:0]: core__GEN_80  ?  core_id_rs_0 [1:0]: core_bypass_src ; 
    wire[61:0] core__GEN_86 ={32'h0, core_inst [31:2]}; 
    wire core__GEN_87 = core_ctrl_killd ==1'h0| core__csr_io_interrupt | core__ibuf_io_inst_0_bits_replay ; 
    wire core_ex_pc_valid = core_ex_reg_valid | core_ex_reg_replay | core_ex_reg_xcpt_interrupt ; 
    wire core_wb_dcache_miss = core_wb_ctrl_mem & core_io_dmem_resp_valid ==1'h0; 
    wire core_replay_ex_structural = core_ex_ctrl_mem & core_io_dmem_req_ready ==1'h0| core_ex_ctrl_div & core__div_io_req_ready ==1'h0; 
    wire core_replay_ex_load_use = core_wb_dcache_miss & core_ex_reg_load_use ; 
    wire core_replay_ex = core_ex_reg_replay | core_ex_reg_valid &( core_replay_ex_structural | core_replay_ex_load_use ); 
    wire core_ctrl_killx = core_take_pc_mem_wb | core_replay_ex | core_ex_reg_valid ==1'h0; 
    wire core_ex_slow_bypass = core_ex_ctrl_mem_cmd ==5'h7| core_ex_reg_mem_size <2'h2; 
    wire core_ex_xcpt = core_ex_reg_xcpt_interrupt | core_ex_reg_xcpt ; 
    wire core_mem_pc_valid = core_mem_reg_valid | core_mem_reg_replay | core_mem_reg_xcpt_interrupt ; 
    wire core_mem_br_target_sign = core_mem_reg_inst [31]; 
    wire core_mem_br_target_hi_hi_hi = core_mem_br_target_sign ; 
    wire[10:0] core_mem_br_target_b30_20 ={{10{ core_mem_br_target_sign }}, core_mem_br_target_sign }; 
    wire[10:0] core_mem_br_target_hi_hi_lo = core_mem_br_target_b30_20 ; 
    wire[7:0] core_mem_br_target_b19_12 ={{7{ core_mem_br_target_sign }}, core_mem_br_target_sign }; 
    wire[7:0] core_mem_br_target_hi_lo_hi = core_mem_br_target_b19_12 ; 
    wire core_mem_br_target_b11 = core_mem_reg_inst [7]; 
    wire core_mem_br_target_hi_lo_lo = core_mem_br_target_b11 ; 
    wire[5:0] core_mem_br_target_b10_5 = core_mem_reg_inst [30:25]; 
    wire[3:0] core_mem_br_target_b4_1 = core_mem_reg_inst [11:8]; 
    wire[9:0] core_mem_br_target_lo_hi ={ core_mem_br_target_b10_5 , core_mem_br_target_b4_1 }; 
    wire[10:0] core_mem_br_target_lo ={ core_mem_br_target_lo_hi , core_mem_br_target_b0 }; 
    wire[8:0] core_mem_br_target_hi_lo ={ core_mem_br_target_hi_lo_hi , core_mem_br_target_hi_lo_lo }; 
    wire[11:0] core_mem_br_target_hi_hi ={ core_mem_br_target_hi_hi_hi , core_mem_br_target_hi_hi_lo }; 
    wire[20:0] core_mem_br_target_hi ={ core_mem_br_target_hi_hi , core_mem_br_target_hi_lo }; 
    wire core_mem_br_target_sign_1 = core_mem_reg_inst [31]; 
    wire core_mem_br_target_hi_hi_hi_1 = core_mem_br_target_sign_1 ; 
    wire[10:0] core_mem_br_target_b30_20_1 ={{10{ core_mem_br_target_sign_1 }}, core_mem_br_target_sign_1 }; 
    wire[10:0] core_mem_br_target_hi_hi_lo_1 = core_mem_br_target_b30_20_1 ; 
    wire[7:0] core_mem_br_target_b19_12_1 = core_mem_reg_inst [19:12]; 
    wire[7:0] core_mem_br_target_hi_lo_hi_1 = core_mem_br_target_b19_12_1 ; 
    wire core_mem_br_target_b11_1 = core_mem_reg_inst [20]; 
    wire core_mem_br_target_hi_lo_lo_1 = core_mem_br_target_b11_1 ; 
    wire[5:0] core_mem_br_target_b10_5_1 = core_mem_reg_inst [30:25]; 
    wire[3:0] core_mem_br_target_b4_1_1 = core_mem_reg_inst [24:21]; 
    wire[9:0] core_mem_br_target_lo_hi_1 ={ core_mem_br_target_b10_5_1 , core_mem_br_target_b4_1_1 }; 
    wire[10:0] core_mem_br_target_lo_1 ={ core_mem_br_target_lo_hi_1 , core_mem_br_target_b0_1 }; 
    wire[8:0] core_mem_br_target_hi_lo_1 ={ core_mem_br_target_hi_lo_hi_1 , core_mem_br_target_hi_lo_lo_1 }; 
    wire[11:0] core_mem_br_target_hi_hi_1 ={ core_mem_br_target_hi_hi_hi_1 , core_mem_br_target_hi_hi_lo_1 }; 
    wire[20:0] core_mem_br_target_hi_1 ={ core_mem_br_target_hi_hi_1 , core_mem_br_target_hi_lo_1 }; 
    wire[3:0] core__GEN_88 = core_mem_reg_rvc  ? 4'h2:4'h4; 
    wire[31:0] core__GEN_89 = core_mem_ctrl_branch & core_mem_br_taken  ? { core_mem_br_target_hi , core_mem_br_target_lo }: core_mem_ctrl_jal  ? { core_mem_br_target_hi_1 , core_mem_br_target_lo_1 }:{{28{ core__GEN_88 [3]}}, core__GEN_88 }; 
    wire[34:0] core__GEN_90 ={ core_mem_reg_pc [33], core_mem_reg_pc }+{{3{ core__GEN_89 [31]}}, core__GEN_89 }; 
    wire[33:0] core_mem_br_target = core__GEN_90 [33:0]; 
    wire[30:0] core_mem_npc_a = core_mem_reg_wdata [63:33]; 
    wire core_mem_npc_msb = core_mem_npc_a ==31'h0|(& core_mem_npc_a ) ?  core_mem_reg_wdata [33]: core_mem_reg_wdata [32]==1'h0; 
    wire[33:0] core_mem_npc =( core_mem_ctrl_jalr | core_mem_reg_sfence  ? { core_mem_npc_msb , core_mem_reg_wdata [32:0]}: core_mem_br_target )&34'h3FFFFFFFE; 
    wire core_mem_wrong_npc = core_ex_pc_valid  ?  core_mem_npc != core_ex_reg_pc : core__ibuf_io_inst_0_valid | core_io_imem_resp_valid  ?  core_mem_npc != core__ibuf_io_pc :1'h1; 
    wire core_mem_npc_misaligned = core__csr_io_status_isa [2]==1'h0& core_mem_npc [1]& core_mem_reg_sfence ==1'h0; 
    wire[63:0] core_mem_int_wdata = core_mem_reg_xcpt ==1'h0&( core_mem_ctrl_jalr ^ core_mem_npc_misaligned ) ? {{30{ core_mem_br_target [33]}}, core_mem_br_target }: core_mem_reg_wdata ; 
    wire core_mem_cfi = core_mem_ctrl_branch | core_mem_ctrl_jalr | core_mem_ctrl_jal ; 
    wire core_mem_cfi_taken = core_mem_ctrl_branch & core_mem_br_taken | core_mem_ctrl_jalr | core_mem_ctrl_jal ; 
    wire core_mem_direction_misprediction = core_mem_ctrl_branch &(| core_mem_br_taken ); 
  assign  core_take_pc_mem = core_mem_reg_valid & core_mem_reg_xcpt ==1'h0&( core_mem_cfi_taken | core_mem_reg_sfence ); 
    wire core__GEN_91 = core_mem_reg_valid & core_mem_reg_flush_pipe ; 
    wire core__GEN_92 =~ core__GEN_91 & core_ex_pc_valid ; 
    wire core__GEN_93 = core_ex_ctrl_mem &( core_ex_ctrl_mem_cmd ==5'h0| core_ex_ctrl_mem_cmd ==5'h10| core_ex_ctrl_mem_cmd ==5'h6| core_ex_ctrl_mem_cmd ==5'h7| core_ex_ctrl_mem_cmd ==5'h4| core_ex_ctrl_mem_cmd ==5'h9| core_ex_ctrl_mem_cmd ==5'hA| core_ex_ctrl_mem_cmd ==5'hB| core_ex_ctrl_mem_cmd ==5'h8| core_ex_ctrl_mem_cmd ==5'hC| core_ex_ctrl_mem_cmd ==5'hD| core_ex_ctrl_mem_cmd ==5'hE| core_ex_ctrl_mem_cmd ==5'hF); 
    wire core__GEN_94 = core_ex_ctrl_mem &( core_ex_ctrl_mem_cmd ==5'h1| core_ex_ctrl_mem_cmd ==5'h11| core_ex_ctrl_mem_cmd ==5'h7| core_ex_ctrl_mem_cmd ==5'h4| core_ex_ctrl_mem_cmd ==5'h9| core_ex_ctrl_mem_cmd ==5'hA| core_ex_ctrl_mem_cmd ==5'hB| core_ex_ctrl_mem_cmd ==5'h8| core_ex_ctrl_mem_cmd ==5'hC| core_ex_ctrl_mem_cmd ==5'hD| core_ex_ctrl_mem_cmd ==5'hE| core_ex_ctrl_mem_cmd ==5'hF); 
    wire core__io_dmem_req_bits_dv_output ; 
    wire core__GEN_95 = core_ex_ctrl_rxs2 &( core_ex_ctrl_mem | core_ex_ctrl_rocc | core_ex_sfence ); 
    wire[1:0] core_size = core_ex_ctrl_rocc  ? 2'h3: core_ex_reg_mem_size ; 
    wire[1:0] core_mem_reg_rs2_size = core_size ; 
    wire[15:0] core__GEN_96 ={ core_ex_rs_1 [7:0], core_ex_rs_1 [7:0]}; 
    wire[31:0] core__GEN_97 ={ core__GEN_96 , core__GEN_96 }; 
    wire[31:0] core__GEN_98 ={ core_ex_rs_1 [15:0], core_ex_rs_1 [15:0]}; 
    wire[63:0] core__GEN_99 = core_mem_reg_rs2_size ==2'h0 ? { core__GEN_97 , core__GEN_97 }: core_mem_reg_rs2_size ==2'h1 ? { core__GEN_98 , core__GEN_98 }: core_mem_reg_rs2_size ==2'h2 ? { core_ex_rs_1 [31:0], core_ex_rs_1 [31:0]}: core_ex_rs_1 ; 
    wire core__GEN_100 = core_ex_ctrl_jalr & core__csr_io_status_debug ; 
    wire core__GEN_101 = core__GEN_100  ? 1'h1: core_ex_ctrl_fence_i ; 
    wire core__GEN_102 = core__GEN_100  ? 1'h1: core_ex_reg_flush_pipe ; 
    wire core_mem_breakpoint = core_mem_reg_load & core__bpu_io_xcpt_ld | core_mem_reg_store & core__bpu_io_xcpt_st ; 
    wire core_mem_debug_breakpoint = core_mem_reg_load & core__bpu_io_debug_ld | core_mem_reg_store & core__bpu_io_debug_st ; 
    wire core_mem_ldst_xcpt = core_mem_debug_breakpoint | core_mem_breakpoint ; 
    wire[3:0] core_mem_ldst_cause = core_mem_debug_breakpoint  ? 4'hE:4'h3; 
    wire core__GEN_103 = core_mem_reg_xcpt_interrupt | core_mem_reg_xcpt ; 
    wire core__GEN_104 = core_mem_reg_valid & core_mem_npc_misaligned ; 
    wire core_mem_xcpt = core__GEN_103 | core__GEN_104 | core_mem_reg_valid & core_mem_ldst_xcpt ; 
    wire[63:0] core_mem_cause = core__GEN_103  ?  core_mem_reg_cause :{60'h0, core__GEN_104  ? 4'h0: core_mem_ldst_cause }; 
    wire core_dcache_kill_mem = core_mem_reg_valid & core_mem_ctrl_wxd & core_io_dmem_replay_next ; 
    wire core_fpu_kill_mem = core_mem_reg_valid & core_mem_ctrl_fp & core_io_fpu_nack_mem ; 
    wire core_replay_mem = core_dcache_kill_mem | core_mem_reg_replay | core_fpu_kill_mem ; 
    wire core_killm_common = core_dcache_kill_mem | core_take_pc_wb | core_mem_reg_xcpt | core_mem_reg_valid ==1'h0; 
    reg core_div_io_kill_REG ; 
  assign  core__GEN_8 = core_killm_common & core_div_io_kill_REG ; 
    wire core_ctrl_killm = core_killm_common | core_mem_xcpt | core_fpu_kill_mem ; 
    wire[63:0] core__GEN_105 = core_mem_reg_xcpt ==1'h0& core_mem_ctrl_fp & core_mem_ctrl_wxd  ?  core_io_fpu_toint_data : core_mem_int_wdata ; 
    wire core__GEN_106 = core_mem_ctrl_rocc | core_mem_reg_sfence ; 
    wire core__GEN_107 = core_mem_ctrl_mem_cmd ==5'h15; 
    wire core__GEN_108 = core_mem_ctrl_mem_cmd ==5'h16; 
    wire core__GEN_109 = core_mem_reg_wphit_0 | core__bpu_io_bpwatch_0_rvalid_0 & core_mem_reg_load | core__bpu_io_bpwatch_0_wvalid_0 & core_mem_reg_store ; 
    wire core__GEN_110 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_pf_st ; 
    wire core__GEN_111 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_pf_ld ; 
    wire core__GEN_112 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_gf_st ; 
    wire core__GEN_113 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_gf_ld ; 
    wire core__GEN_114 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_ae_st ; 
    wire core__GEN_115 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_ae_ld ; 
    wire core__GEN_116 = core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_ma_st ; 
  assign  core_wb_xcpt = core_wb_reg_xcpt | core__GEN_110 | core__GEN_111 | core__GEN_112 | core__GEN_113 | core__GEN_114 | core__GEN_115 | core__GEN_116 | core_wb_reg_valid & core_wb_ctrl_mem & core_io_dmem_s2_xcpt_ma_ld ; 
  assign  core_wb_cause = core_wb_reg_xcpt  ?  core_wb_reg_cause :{59'h0, core__GEN_110  ? 5'hF: core__GEN_111  ? 5'hD: core__GEN_112  ? 5'h17: core__GEN_113  ? 5'h15:{2'h0, core__GEN_114  ? 3'h7: core__GEN_115  ? 3'h5: core__GEN_116  ? 3'h6:3'h4}}; 
    wire core_wb_pc_valid = core_wb_reg_valid | core_wb_reg_replay | core_wb_reg_xcpt ; 
    wire core_wb_wxd = core_wb_reg_valid & core_wb_ctrl_wxd ; 
    wire core_wb_set_sboard = core_wb_ctrl_div | core_wb_dcache_miss | core_wb_ctrl_rocc ; 
    wire core_replay_wb_common = core_io_dmem_s2_nack | core_wb_reg_replay ; 
    wire core_replay_wb_rocc = core_wb_reg_valid & core_wb_ctrl_rocc & core_io_rocc_cmd_ready ==1'h0; 
    wire core_replay_wb_csr = core_wb_reg_valid & core__csr_io_rw_stall ; 
    wire core_replay_wb = core_replay_wb_common | core_replay_wb_rocc | core_replay_wb_csr ; 
  assign  core_take_pc_wb = core_replay_wb | core_wb_xcpt | core__csr_io_eret | core_wb_reg_flush_pipe ; 
    wire core_dmem_resp_xpu = core_io_dmem_resp_bits_tag [0]==1'h0; 
    wire core_dmem_resp_fpu = core_io_dmem_resp_bits_tag [0]; 
    wire[4:0] core_dmem_resp_waddr = core_io_dmem_resp_bits_tag [5:1]; 
    wire core_dmem_resp_valid = core_io_dmem_resp_valid & core_io_dmem_resp_bits_has_data ; 
    wire core_dmem_resp_replay = core_dmem_resp_valid & core_io_dmem_resp_bits_replay ; 
    wire core__GEN_117 = core_dmem_resp_replay & core_dmem_resp_xpu ; 
  assign  core__GEN_7 = core__GEN_117  ? 1'h0: core_wb_wxd ==1'h0; 
    wire[4:0] core_ll_waddr = core__GEN_117  ?  core_dmem_resp_waddr : core__div_io_resp_bits_tag ; 
    wire core_ll_wen = core__GEN_117  ? 1'h1: core__GEN_7 & core__div_io_resp_valid ; 
  assign  core_wb_valid = core_wb_reg_valid & core_replay_wb ==1'h0& core_wb_xcpt ==1'h0; 
    wire core_wb_wen = core_wb_valid & core_wb_ctrl_wxd ; 
    wire core_rf_wen = core_wb_wen | core_ll_wen ; 
    wire[4:0] core_rf_waddr = core_ll_wen  ?  core_ll_waddr : core_wb_waddr ; 
    wire[4:0] core_xrfWriteBundle_wrdst = core_rf_waddr ; 
  assign  core_rf_wdata = core_dmem_resp_valid & core_dmem_resp_xpu  ?  core_io_dmem_resp_bits_data : core_ll_wen  ?  core_ll_wdata :(| core_wb_ctrl_csr ) ?  core__csr_io_rw_rdata : core_wb_reg_wdata ; 
    wire[63:0] core_coreMonitorBundle_wrdata = core_rf_wdata ; 
    wire[63:0] core_xrfWriteBundle_wrdata = core_rf_wdata ; 
    wire core__GEN_118 =| core_rf_waddr ; 
    wire core__GEN_119 = core_rf_wen & core__GEN_118 ; 
  assign  core__GEN_6 =~ core_rf_waddr ; 
  assign  core__GEN_5 = core_rf_wen  ?  core__GEN_118 :1'h0; 
    wire core__GEN_120 = core_rf_waddr == core_id_raddr1 ; 
  assign  core_id_rs_0 = core_rf_wen  ? ( core__GEN_118  ? ( core__GEN_120  ?  core_rf_wdata : core__rf_ext_R1_data ): core__rf_ext_R1_data ): core__rf_ext_R1_data ; 
    wire core__GEN_121 = core_rf_waddr == core_id_raddr2 ; 
  assign  core_id_rs_1 = core_rf_wen  ? ( core__GEN_118  ? ( core__GEN_121  ?  core_rf_wdata : core__rf_ext_R0_data ): core__rf_ext_R0_data ): core__rf_ext_R0_data ; 
  assign  core__GEN_4 ={(&( core_wb_reg_raw_inst [1:0])) ?  core_wb_reg_inst [31:16]:16'h0, core_wb_reg_raw_inst [15:0]}; 
    wire core_tval_dmem_addr = core_wb_reg_xcpt ==1'h0; 
    wire core_tval_any_addr = core_tval_dmem_addr | core_wb_reg_cause ==64'h3| core_wb_reg_cause ==64'h1| core_wb_reg_cause ==64'hC| core_wb_reg_cause ==64'h14; 
    wire core_tval_inst = core_wb_reg_cause ==64'h2; 
    wire core_tval_valid = core_wb_xcpt &( core_tval_any_addr | core_tval_inst ); 
  assign  core__GEN_3 = core_wb_xcpt &( core_tval_any_addr & core__csr_io_status_v | core_tval_dmem_addr & core_wb_reg_hls_or_dv ); 
    wire[30:0] core_csr_io_tval_a = core_wb_reg_wdata [63:33]; 
    wire core_csr_io_tval_msb = core_csr_io_tval_a ==31'h0|(& core_csr_io_tval_a ) ?  core_wb_reg_wdata [33]: core_wb_reg_wdata [32]==1'h0; 
  assign  core__GEN_2 = core_tval_valid  ? { core_csr_io_tval_msb , core_wb_reg_wdata [32:0]}:34'h0; 
    wire core_csr_io_htval_htval_valid_imem = core_wb_reg_xcpt & core_wb_reg_cause ==64'h14; 
    wire[33:0] core_csr_io_htval_htval_imem = core_csr_io_htval_htval_valid_imem  ?  core_io_imem_gpa_bits :34'h0; 
    wire core__GEN_122 =( core_csr_io_htval_htval_valid_imem ==1'h0| core_io_imem_gpa_valid )==1'h0; 
    wire core_csr_io_htval_htval_valid_dmem = core_wb_xcpt & core_tval_dmem_addr &(|{ core_io_dmem_s2_xcpt_gf_ld , core_io_dmem_s2_xcpt_gf_st })&(|{ core_io_dmem_s2_xcpt_pf_ld , core_io_dmem_s2_xcpt_pf_st })==1'h0; 
    wire[33:0] core_csr_io_htval_htval_dmem = core_csr_io_htval_htval_valid_dmem  ?  core_io_dmem_s2_gpa :34'h0; 
  assign  core__GEN_1 ={6'h0, core_csr_io_htval_htval_dmem | core_csr_io_htval_htval_imem }; 
  assign  core__wb_reg_inst_31to20 = core_wb_reg_inst [31:20]; 
  assign  core__GEN_0 = core_wb_ctrl_csr &~( core_wb_reg_valid  ? 3'h0:3'h4); 
    wire core__GEN_123 = core_id_ctrl_rxs1 &(| core_id_raddr1 ); 
    wire core__GEN_124 = core_id_ctrl_rxs2 &(| core_id_raddr2 ); 
    wire core__GEN_125 = core_id_ctrl_wxd &(| core_id_waddr ); reg[31:0] core__r ; 
    wire[31:0] core_r ={ core__r [31:1],1'h0}; 
    wire[31:0] core__GEN_126 = core_r &~( core_ll_wen  ? 32'h1<< core_ll_waddr :32'h0); 
    wire core__GEN_127 = core_ll_wen |1'h0; 
    wire[31:0] core__GEN_128 = core_r >> core_id_raddr1 ; 
    wire[31:0] core__GEN_129 = core_r >> core_id_raddr2 ; 
    wire[31:0] core__GEN_130 = core_r >> core_id_waddr ; 
    wire core_id_sboard_hazard = core__GEN_123 & core__GEN_128 [0]&( core_ll_wen & core_ll_waddr == core_id_raddr1 )==1'h0| core__GEN_124 & core__GEN_129 [0]&( core_ll_wen & core_ll_waddr == core_id_raddr2 )==1'h0| core__GEN_125 & core__GEN_130 [0]&( core_ll_wen & core_ll_waddr == core_id_waddr )==1'h0; 
    wire core__GEN_131 = core_wb_set_sboard & core_wb_wen ; 
    wire[31:0] core__GEN_132 = core__GEN_126 |( core__GEN_131  ? 32'h1<< core_wb_waddr :32'h0); 
    wire core__GEN_133 = core__GEN_127 | core__GEN_131 ; 
    wire core_ex_cannot_bypass =(| core_ex_ctrl_csr )| core_ex_ctrl_jalr | core_ex_ctrl_mem | core_ex_ctrl_mul | core_ex_ctrl_div | core_ex_ctrl_fp | core_ex_ctrl_rocc ; 
    wire core_data_hazard_ex = core_ex_ctrl_wxd &( core__GEN_123 & core_id_raddr1 == core_ex_waddr | core__GEN_124 & core_id_raddr2 == core_ex_waddr | core__GEN_125 & core_id_waddr == core_ex_waddr ); 
    wire core_fp_data_hazard_ex = core_id_ctrl_fp & core_ex_ctrl_wfd &( core_io_fpu_dec_ren1 & core_id_raddr1 == core_ex_waddr | core_io_fpu_dec_ren2 & core_id_raddr2 == core_ex_waddr | core_io_fpu_dec_ren3 & core_id_raddr3 == core_ex_waddr | core_io_fpu_dec_wen & core_id_waddr == core_ex_waddr ); 
    wire core_id_ex_hazard = core_ex_reg_valid &( core_data_hazard_ex & core_ex_cannot_bypass | core_fp_data_hazard_ex ); 
    wire core_mem_mem_cmd_bh = core_mem_reg_slow_bypass &1'h1; 
    wire core_mem_cannot_bypass =(| core_mem_ctrl_csr )| core_mem_ctrl_mem & core_mem_mem_cmd_bh | core_mem_ctrl_mul | core_mem_ctrl_div | core_mem_ctrl_fp | core_mem_ctrl_rocc ; 
    wire core_data_hazard_mem = core_mem_ctrl_wxd &( core__GEN_123 & core_id_raddr1 == core_mem_waddr | core__GEN_124 & core_id_raddr2 == core_mem_waddr | core__GEN_125 & core_id_waddr == core_mem_waddr ); 
    wire core_fp_data_hazard_mem = core_id_ctrl_fp & core_mem_ctrl_wfd &( core_io_fpu_dec_ren1 & core_id_raddr1 == core_mem_waddr | core_io_fpu_dec_ren2 & core_id_raddr2 == core_mem_waddr | core_io_fpu_dec_ren3 & core_id_raddr3 == core_mem_waddr | core_io_fpu_dec_wen & core_id_waddr == core_mem_waddr ); 
    wire core_id_mem_hazard = core_mem_reg_valid &( core_data_hazard_mem & core_mem_cannot_bypass | core_fp_data_hazard_mem ); 
  assign  core_id_load_use = core_mem_reg_valid & core_data_hazard_mem & core_mem_ctrl_mem ; 
    wire core_data_hazard_wb = core_wb_ctrl_wxd &( core__GEN_123 & core_id_raddr1 == core_wb_waddr | core__GEN_124 & core_id_raddr2 == core_wb_waddr | core__GEN_125 & core_id_waddr == core_wb_waddr ); 
    wire core_fp_data_hazard_wb = core_id_ctrl_fp & core_wb_ctrl_wfd &( core_io_fpu_dec_ren1 & core_id_raddr1 == core_wb_waddr | core_io_fpu_dec_ren2 & core_id_raddr2 == core_wb_waddr | core_io_fpu_dec_ren3 & core_id_raddr3 == core_wb_waddr | core_io_fpu_dec_wen & core_id_waddr == core_wb_waddr ); 
    wire core_id_wb_hazard = core_wb_reg_valid &( core_data_hazard_wb & core_wb_set_sboard | core_fp_data_hazard_wb ); 
    reg core_dcache_blocked_blocked ; 
    wire core_dcache_blocked = core_dcache_blocked_blocked & core_io_dmem_perf_grant ==1'h0; 
    reg core_rocc_blocked ; 
    wire core__io_rocc_cmd_valid_output ; 
    wire core_ctrl_stalld = core_id_ex_hazard | core_id_mem_hazard | core_id_wb_hazard | core_id_sboard_hazard | core__csr_io_singleStep &( core_ex_reg_valid | core_mem_reg_valid | core_wb_reg_valid )| core_id_csr_en & core__csr_io_decode_0_fp_csr & core_io_fpu_fcsr_rdy ==1'h0| core_id_ctrl_mem & core_dcache_blocked | core_id_ctrl_rocc & core_rocc_blocked | core_id_ctrl_div &(( core__div_io_req_ready | core__div_io_resp_valid & core_wb_wxd ==1'h0)==1'h0| core__GEN_9 )| core_clock_en ==1'h0| core_id_do_fence | core__csr_io_csr_stall | core_id_reg_pause | core_io_traceStall ; 
  assign  core_ctrl_killd = core__ibuf_io_inst_0_valid ==1'h0| core__ibuf_io_inst_0_bits_replay | core_take_pc_mem_wb | core_ctrl_stalld | core__csr_io_interrupt ; 
    wire[33:0] core__io_imem_req_bits_pc_output = core_wb_xcpt | core__csr_io_eret  ?  core__csr_io_evec : core_replay_wb  ?  core_wb_reg_pc : core_mem_npc ; 
    reg core_io_imem_progress_REG ; 
    wire core__io_imem_sfence_valid_output = core_wb_reg_valid & core_wb_reg_sfence ; 
    wire core__io_imem_sfence_bits_rs1_output = core_wb_reg_mem_size [0]; 
    wire core__io_imem_sfence_bits_rs2_output = core_wb_reg_mem_size [1]; 
    wire[32:0] core__io_imem_sfence_bits_addr_output = core_wb_reg_wdata [32:0]; 
    wire core__io_imem_sfence_bits_asid_output = core_wb_reg_rs2 [0]; 
  assign  core__GEN = core_ctrl_stalld ==1'h0; 
    wire[34:0] core__GEN_134 ={1'h0, core_mem_reg_pc }+{33'h0, core_mem_reg_rvc  ? 2'h0:2'h2}; 
    wire[33:0] core__GEN_135 = core__GEN_134 [33:0]; 
    wire[32:0] core__io_imem_btb_update_bits_br_pc_output = core__GEN_135 [32:0]; 
    wire[32:0] core__io_imem_btb_update_bits_pc_output =~(~ core__io_imem_btb_update_bits_br_pc_output |33'h3); 
  assign  core__io_dmem_req_valid_output = core_ex_reg_valid & core_ex_ctrl_mem ; 
    wire[5:0] core_ex_dcache_tag ={ core_ex_waddr , core_ex_ctrl_fp }; 
    wire[30:0] core_io_dmem_req_bits_addr_a = core_ex_rs_0 [63:33]; 
    wire core_io_dmem_req_bits_addr_msb = core_io_dmem_req_bits_addr_a ==31'h0|(& core_io_dmem_req_bits_addr_a ) ?  core__alu_io_adder_out [33]: core__alu_io_adder_out [32]==1'h0; 
  assign  core__io_dmem_req_bits_dv_output = core_ex_reg_hls | core__csr_io_status_dv ; 
  assign  core__io_rocc_cmd_valid_output = core_wb_reg_valid & core_wb_ctrl_rocc & core_replay_wb_common ==1'h0; 
    wire[6:0] core__io_rocc_cmd_bits_inst_WIRE_opcode = core__io_rocc_cmd_bits_inst_WIRE_1 [6:0]; 
    wire[4:0] core__io_rocc_cmd_bits_inst_WIRE_rd = core__io_rocc_cmd_bits_inst_WIRE_1 [11:7]; 
    wire core__io_rocc_cmd_bits_inst_WIRE_xs2 = core__io_rocc_cmd_bits_inst_WIRE_1 [12]; 
    wire core__io_rocc_cmd_bits_inst_WIRE_xs1 = core__io_rocc_cmd_bits_inst_WIRE_1 [13]; 
    wire core__io_rocc_cmd_bits_inst_WIRE_xd = core__io_rocc_cmd_bits_inst_WIRE_1 [14]; 
    wire[4:0] core__io_rocc_cmd_bits_inst_WIRE_rs1 = core__io_rocc_cmd_bits_inst_WIRE_1 [19:15]; 
    wire[4:0] core__io_rocc_cmd_bits_inst_WIRE_rs2 = core__io_rocc_cmd_bits_inst_WIRE_1 [24:20]; 
    wire[6:0] core__io_rocc_cmd_bits_inst_WIRE_funct = core__io_rocc_cmd_bits_inst_WIRE_1 [31:25]; 
    wire core_unpause = core__csr_io_time [4:0]==5'h0| core__csr_io_inhibit_cycle | core_io_dmem_perf_release | core_take_pc_mem_wb ; 
    reg core_icache_blocked_REG ; 
    wire core_icache_blocked =( core_io_imem_resp_valid | core_icache_blocked_REG )==1'h0; 
    wire[63:0] core_coreMonitorBundle_hartid ={63'h0, core_io_hartid }; 
    wire[31:0] core_coreMonitorBundle_timer = core__csr_io_time [31:0]; 
    wire core_coreMonitorBundle_valid = core__csr_io_trace_0_valid & core__csr_io_trace_0_exception ==1'h0; 
    wire[63:0] core_coreMonitorBundle_pc ={ core__csr_io_trace_0_iaddr [33] ? 30'h3FFFFFFF:30'h0, core__csr_io_trace_0_iaddr }; 
    wire core_coreMonitorBundle_wrenx = core_wb_wen & core_wb_set_sboard ==1'h0; 
    wire[4:0] core_coreMonitorBundle_rd0src = core_wb_reg_inst [19:15]; reg[63:0] core_coreMonitorBundle_rd0val_REG ; reg[63:0] core_coreMonitorBundle_rd0val_REG_1 ; 
    wire[63:0] core_coreMonitorBundle_rd0val = core_coreMonitorBundle_rd0val_REG_1 ; 
    wire[4:0] core_coreMonitorBundle_rd1src = core_wb_reg_inst [24:20]; reg[63:0] core_coreMonitorBundle_rd1val_REG ; reg[63:0] core_coreMonitorBundle_rd1val_REG_1 ; 
    wire[63:0] core_coreMonitorBundle_rd1val = core_coreMonitorBundle_rd1val_REG_1 ; 
  always @( posedge  core_clock )
         begin 
             if ( core_reset ==1'h0& core__GEN_122 )
                 begin 
                     if (1)$error("Assertion failed\n    at RocketCore.scala:718 assert(!htval_valid_imem || io.imem.gpa.valid)\n");
                     if (1)$fatal;
                 end 
             if ((1)& core__csr_io_trace_0_valid & core_reset ==1'h0)$fwrite(32'h80000002,"C%d: %d [%d] pc=[%x] W[r%d=%x][%d] R[r%d=%x] R[r%d=%x] inst=[%x] DASM(%x)\n", core_io_hartid , core_coreMonitorBundle_timer , core_coreMonitorBundle_valid , core_coreMonitorBundle_pc , core_wb_ctrl_wxd | core_wb_ctrl_wfd  ?  core_coreMonitorBundle_wrdst :5'h0, core_coreMonitorBundle_wrenx  ?  core_coreMonitorBundle_wrdata :64'h0, core_coreMonitorBundle_wrenx , core_wb_ctrl_rxs1 | core_wb_ctrl_rfs1  ?  core_coreMonitorBundle_rd0src :5'h0, core_wb_ctrl_rxs1 | core_wb_ctrl_rfs1  ?  core_coreMonitorBundle_rd0val :64'h0, core_wb_ctrl_rxs2 | core_wb_ctrl_rfs2  ?  core_coreMonitorBundle_rd1src :5'h0, core_wb_ctrl_rxs2 | core_wb_ctrl_rfs2  ?  core_coreMonitorBundle_rd1val :64'h0, core_coreMonitorBundle_inst , core_coreMonitorBundle_inst );
         end
    wire[63:0] core_xrfWriteBundle_hartid ={63'h0, core_io_hartid }; 
    wire[31:0] core_xrfWriteBundle_timer = core__csr_io_time [31:0]; 
    wire[63:0] core_xrfWriteBundle_pc =64'h0; 
    wire core_xrfWriteBundle_wrenx = core_rf_wen &( core__csr_io_trace_0_valid & core_wb_wen & core_wb_waddr == core_rf_waddr )==1'h0; 
    wire[4:0] core_xrfWriteBundle_rd0src =5'h0; 
    wire[63:0] core_xrfWriteBundle_rd0val =64'h0; 
    wire[4:0] core_xrfWriteBundle_rd1src =5'h0; 
    wire[63:0] core_xrfWriteBundle_rd1val =64'h0; 
    wire[31:0] core_xrfWriteBundle_inst =32'h0;  
    wire core_PlusArgTimeout_clock;
    wire core_PlusArgTimeout_reset;
    wire[31:0] core_PlusArgTimeout_io_count;

    wire[31:0] core_PlusArgTimeout__plusarg_reader_out ;  
    wire core_PlusArgTimeout__GEN = core_PlusArgTimeout_io_count < core_PlusArgTimeout__plusarg_reader_out ==1'h0; 
  always @( posedge  core_PlusArgTimeout_clock )
         begin 
             if ( core_PlusArgTimeout__plusarg_reader_out >32'h0& core_PlusArgTimeout_reset ==1'h0& core_PlusArgTimeout__GEN )
                 begin 
                     if (1)$error("Assertion failed: Timeout exceeded: Kill the emulation after INT rdtime cycles. Off if 0.\n    at PlusArg.scala:64 assert (io.count < max, s\"Timeout exceeded: $docstring\")\n");
                     if (1)$fatal;
                 end 
         end
 
    assign core_PlusArgTimeout_clock = core_clock;
    assign core_PlusArgTimeout_reset = core_reset;
    assign core_PlusArgTimeout_io_count = core__csr_io_time_31to0;
     
  assign  core__csr_io_time_31to0 = core__csr_io_time [31:0]; 
  always @( posedge  core_clock )
         begin 
             if ( core_reset )
                 begin  
                     core_clock_en_reg  <=1'h1; 
                     core_id_reg_fence  <=1'h0; 
                     core__r  <=32'h0;
                 end 
              else 
                 begin 
                     if ( core__GEN_65 )
                         begin 
                             if ( core_id_fence_next ) 
                                 core_id_reg_fence  <=1'h1;
                              else 
                                 if ( core__GEN_59 ) 
                                     core_id_reg_fence  <=1'h0;
                                  else 
                                     begin 
                                     end 
                         end 
                      else 
                         if ( core__GEN_59 ) 
                             core_id_reg_fence  <=1'h0;
                          else 
                             begin 
                             end 
                     if ( core__GEN_133 ) 
                         core__r  <= core__GEN_132 ;
                      else 
                         if ( core__GEN_127 ) 
                             core__r  <= core__GEN_126 ;
                          else 
                             begin 
                             end 
                 end 
         end
  always @( posedge  core_clock )
         begin 
             if ( core_unpause ) 
                 core_id_reg_pause  <=1'h0;
              else 
                 if ( core__GEN_65 )
                     begin 
                         if ( core__GEN_66 ) 
                             core_id_reg_pause  <=1'h1;
                          else 
                             begin 
                             end 
                     end 
                  else 
                     begin 
                     end  
             core_imem_might_request_reg  <= core_ex_pc_valid | core_mem_pc_valid | core__io_ptw_customCSRs_csrs_0_value_output [1];
             if ( core__GEN_65 )
                 begin  
                     core_ex_ctrl_legal  <= core_id_ctrl_legal ; 
                     core_ex_ctrl_fp  <= core_id_ctrl_fp ; 
                     core_ex_ctrl_rocc  <= core_id_ctrl_rocc ; 
                     core_ex_ctrl_branch  <= core_id_ctrl_branch ; 
                     core_ex_ctrl_jal  <= core_id_ctrl_jal ; 
                     core_ex_ctrl_jalr  <= core_id_ctrl_jalr ; 
                     core_ex_ctrl_rxs2  <= core_id_ctrl_rxs2 ; 
                     core_ex_ctrl_rxs1  <= core_id_ctrl_rxs1 ; 
                     core_ex_ctrl_sel_alu2  <= core__GEN_74 ; 
                     core_ex_ctrl_sel_alu1  <= core__GEN_73 ; 
                     core_ex_ctrl_sel_imm  <= core_id_ctrl_sel_imm ; 
                     core_ex_ctrl_alu_dw  <= core__GEN_69 ; 
                     core_ex_ctrl_alu_fn  <= core__GEN_68 ; 
                     core_ex_ctrl_mem  <= core_id_ctrl_mem ; 
                     core_ex_ctrl_mem_cmd  <= core__GEN_79 ; 
                     core_ex_ctrl_rfs1  <= core_id_ctrl_rfs1 ; 
                     core_ex_ctrl_rfs2  <= core_id_ctrl_rfs2 ; 
                     core_ex_ctrl_rfs3  <= core_id_ctrl_rfs3 ; 
                     core_ex_ctrl_wfd  <= core_id_ctrl_wfd ; 
                     core_ex_ctrl_mul  <= core_id_ctrl_mul ; 
                     core_ex_ctrl_div  <= core_id_ctrl_div ; 
                     core_ex_ctrl_wxd  <= core_id_ctrl_wxd ; 
                     core_ex_ctrl_csr  <= core_id_csr ; 
                     core_ex_ctrl_fence_i  <= core_id_ctrl_fence_i ; 
                     core_ex_ctrl_fence  <= core_id_ctrl_fence ; 
                     core_ex_ctrl_amo  <= core_id_ctrl_amo ; 
                     core_ex_ctrl_dp  <= core_id_ctrl_dp ; 
                     core_ex_reg_rvc  <= core__GEN_71 ; 
                     core_ex_reg_flush_pipe  <= core__GEN_75 ; 
                     core_ex_reg_load_use  <= core_id_load_use ; 
                     core_ex_reg_mem_size  <= core__GEN_77 ; 
                     core_ex_reg_hls  <=1'h0; 
                     core_ex_reg_rs_bypass_0  <= core__GEN_84 ; 
                     core_ex_reg_rs_bypass_1  <= core_do_bypass_1 ; 
                     core_ex_reg_rs_lsb_0  <= core__GEN_85 ; 
                     core_ex_reg_rs_lsb_1  <= core__GEN_82 ;
                     if ( core__GEN_83 ) 
                         core_ex_reg_rs_msb_0  <= core__GEN_86 ;
                      else 
                         if ( core__GEN_80 ) 
                             core_ex_reg_rs_msb_0  <= core_id_rs_0 [63:2];
                          else 
                             begin 
                             end 
                     if ( core__GEN_81 ) 
                         core_ex_reg_rs_msb_1  <= core_id_rs_1 [63:2];
                      else 
                         begin 
                         end 
                 end 
              else 
                 begin 
                 end 
             if ( core__GEN_91 ) 
                 core_mem_reg_sfence  <=1'h0;
              else 
                 if ( core_ex_pc_valid )
                     begin  
                         core_mem_ctrl_legal  <= core_ex_ctrl_legal ; 
                         core_mem_ctrl_fp  <= core_ex_ctrl_fp ; 
                         core_mem_ctrl_rocc  <= core_ex_ctrl_rocc ; 
                         core_mem_ctrl_branch  <= core_ex_ctrl_branch ; 
                         core_mem_ctrl_jal  <= core_ex_ctrl_jal ; 
                         core_mem_ctrl_jalr  <= core_ex_ctrl_jalr ; 
                         core_mem_ctrl_rxs2  <= core_ex_ctrl_rxs2 ; 
                         core_mem_ctrl_rxs1  <= core_ex_ctrl_rxs1 ; 
                         core_mem_ctrl_sel_alu2  <= core_ex_ctrl_sel_alu2 ; 
                         core_mem_ctrl_sel_alu1  <= core_ex_ctrl_sel_alu1 ; 
                         core_mem_ctrl_sel_imm  <= core_ex_ctrl_sel_imm ; 
                         core_mem_ctrl_alu_dw  <= core_ex_ctrl_alu_dw ; 
                         core_mem_ctrl_alu_fn  <= core_ex_ctrl_alu_fn ; 
                         core_mem_ctrl_mem  <= core_ex_ctrl_mem ; 
                         core_mem_ctrl_mem_cmd  <= core_ex_ctrl_mem_cmd ; 
                         core_mem_ctrl_rfs1  <= core_ex_ctrl_rfs1 ; 
                         core_mem_ctrl_rfs2  <= core_ex_ctrl_rfs2 ; 
                         core_mem_ctrl_rfs3  <= core_ex_ctrl_rfs3 ; 
                         core_mem_ctrl_wfd  <= core_ex_ctrl_wfd ; 
                         core_mem_ctrl_mul  <= core_ex_ctrl_mul ; 
                         core_mem_ctrl_div  <= core_ex_ctrl_div ; 
                         core_mem_ctrl_wxd  <= core_ex_ctrl_wxd ; 
                         core_mem_ctrl_csr  <= core_ex_ctrl_csr ; 
                         core_mem_ctrl_fence_i  <= core__GEN_101 ; 
                         core_mem_ctrl_fence  <= core_ex_ctrl_fence ; 
                         core_mem_ctrl_amo  <= core_ex_ctrl_amo ; 
                         core_mem_ctrl_dp  <= core_ex_ctrl_dp ; 
                         core_mem_reg_rvc  <= core_ex_reg_rvc ; 
                         core_mem_reg_btb_resp_cfiType  <= core_ex_reg_btb_resp_cfiType ; 
                         core_mem_reg_btb_resp_taken  <= core_ex_reg_btb_resp_taken ; 
                         core_mem_reg_btb_resp_mask  <= core_ex_reg_btb_resp_mask ; 
                         core_mem_reg_btb_resp_bridx  <= core_ex_reg_btb_resp_bridx ; 
                         core_mem_reg_btb_resp_target  <= core_ex_reg_btb_resp_target ; 
                         core_mem_reg_btb_resp_entry  <= core_ex_reg_btb_resp_entry ; 
                         core_mem_reg_btb_resp_bht_history  <= core_ex_reg_btb_resp_bht_history ; 
                         core_mem_reg_btb_resp_bht_value  <= core_ex_reg_btb_resp_bht_value ; 
                         core_mem_reg_flush_pipe  <= core__GEN_102 ; 
                         core_mem_reg_cause  <= core_ex_reg_cause ; 
                         core_mem_reg_slow_bypass  <= core_ex_slow_bypass ; 
                         core_mem_reg_load  <= core__GEN_93 ; 
                         core_mem_reg_store  <= core__GEN_94 ; 
                         core_mem_reg_sfence  <= core_ex_sfence ; 
                         core_mem_reg_pc  <= core_ex_reg_pc ; 
                         core_mem_reg_inst  <= core_ex_reg_inst ; 
                         core_mem_reg_mem_size  <= core_ex_reg_mem_size ; 
                         core_mem_reg_hls_or_dv  <= core__io_dmem_req_bits_dv_output ; 
                         core_mem_reg_raw_inst  <= core_ex_reg_raw_inst ; 
                         core_mem_reg_wdata  <= core__alu_io_out ;
                         if ( core__GEN_95 ) 
                             core_mem_reg_rs2  <= core__GEN_99 ;
                          else 
                             begin 
                             end  
                         core_mem_br_taken  <= core__alu_io_cmp_out ; 
                         core_mem_reg_wphit_0  <= core_ex_reg_wphit_0 ;
                     end 
                  else 
                     begin 
                     end 
             if ( core_mem_pc_valid )
                 begin  
                     core_wb_ctrl_legal  <= core_mem_ctrl_legal ; 
                     core_wb_ctrl_fp  <= core_mem_ctrl_fp ; 
                     core_wb_ctrl_rocc  <= core_mem_ctrl_rocc ; 
                     core_wb_ctrl_branch  <= core_mem_ctrl_branch ; 
                     core_wb_ctrl_jal  <= core_mem_ctrl_jal ; 
                     core_wb_ctrl_jalr  <= core_mem_ctrl_jalr ; 
                     core_wb_ctrl_rxs2  <= core_mem_ctrl_rxs2 ; 
                     core_wb_ctrl_rxs1  <= core_mem_ctrl_rxs1 ; 
                     core_wb_ctrl_sel_alu2  <= core_mem_ctrl_sel_alu2 ; 
                     core_wb_ctrl_sel_alu1  <= core_mem_ctrl_sel_alu1 ; 
                     core_wb_ctrl_sel_imm  <= core_mem_ctrl_sel_imm ; 
                     core_wb_ctrl_alu_dw  <= core_mem_ctrl_alu_dw ; 
                     core_wb_ctrl_alu_fn  <= core_mem_ctrl_alu_fn ; 
                     core_wb_ctrl_mem  <= core_mem_ctrl_mem ; 
                     core_wb_ctrl_mem_cmd  <= core_mem_ctrl_mem_cmd ; 
                     core_wb_ctrl_rfs1  <= core_mem_ctrl_rfs1 ; 
                     core_wb_ctrl_rfs2  <= core_mem_ctrl_rfs2 ; 
                     core_wb_ctrl_rfs3  <= core_mem_ctrl_rfs3 ; 
                     core_wb_ctrl_wfd  <= core_mem_ctrl_wfd ; 
                     core_wb_ctrl_mul  <= core_mem_ctrl_mul ; 
                     core_wb_ctrl_div  <= core_mem_ctrl_div ; 
                     core_wb_ctrl_wxd  <= core_mem_ctrl_wxd ; 
                     core_wb_ctrl_csr  <= core_mem_ctrl_csr ; 
                     core_wb_ctrl_fence_i  <= core_mem_ctrl_fence_i ; 
                     core_wb_ctrl_fence  <= core_mem_ctrl_fence ; 
                     core_wb_ctrl_amo  <= core_mem_ctrl_amo ; 
                     core_wb_ctrl_dp  <= core_mem_ctrl_dp ; 
                     core_wb_reg_cause  <= core_mem_cause ; 
                     core_wb_reg_sfence  <= core_mem_reg_sfence ; 
                     core_wb_reg_pc  <= core_mem_reg_pc ; 
                     core_wb_reg_mem_size  <= core_mem_reg_mem_size ; 
                     core_wb_reg_hls_or_dv  <= core_mem_reg_hls_or_dv ; 
                     core_wb_reg_hfence_v  <= core__GEN_107 ; 
                     core_wb_reg_hfence_g  <= core__GEN_108 ; 
                     core_wb_reg_inst  <= core_mem_reg_inst ; 
                     core_wb_reg_raw_inst  <= core_mem_reg_raw_inst ; 
                     core_wb_reg_wdata  <= core__GEN_105 ;
                     if ( core__GEN_106 ) 
                         core_wb_reg_rs2  <= core_mem_reg_rs2 ;
                      else 
                         begin 
                         end  
                     core_wb_reg_wphit_0  <= core__GEN_109 ;
                 end 
              else 
                 begin 
                 end  
             core_ex_reg_xcpt_interrupt  <= core_take_pc_mem_wb ==1'h0& core__ibuf_io_inst_0_valid & core__csr_io_interrupt ; 
             core_ex_reg_valid  <= core_ctrl_killd ==1'h0;
             if ( core__GEN_87 )
                 begin  
                     core_ex_reg_btb_resp_cfiType  <= core__ibuf_io_btb_resp_cfiType ; 
                     core_ex_reg_btb_resp_taken  <= core__ibuf_io_btb_resp_taken ; 
                     core_ex_reg_btb_resp_mask  <= core__ibuf_io_btb_resp_mask ; 
                     core_ex_reg_btb_resp_bridx  <= core__ibuf_io_btb_resp_bridx ; 
                     core_ex_reg_btb_resp_target  <= core__ibuf_io_btb_resp_target ; 
                     core_ex_reg_btb_resp_entry  <= core__ibuf_io_btb_resp_entry ; 
                     core_ex_reg_btb_resp_bht_history  <= core__ibuf_io_btb_resp_bht_history ; 
                     core_ex_reg_btb_resp_bht_value  <= core__ibuf_io_btb_resp_bht_value ; 
                     core_ex_reg_cause  <= core_id_cause ; 
                     core_ex_reg_pc  <= core__ibuf_io_pc ; 
                     core_ex_reg_inst  <= core__ibuf_io_inst_0_bits_inst_bits ; 
                     core_ex_reg_raw_inst  <= core__ibuf_io_inst_0_bits_raw ; 
                     core_ex_reg_wphit_0  <= core__bpu_io_bpwatch_0_ivalid_0 ;
                 end 
              else 
                 begin 
                 end  
             core_ex_reg_xcpt  <= core_ctrl_killd ==1'h0& core_id_xcpt ; 
             core_ex_reg_replay  <= core_take_pc_mem_wb ==1'h0& core__ibuf_io_inst_0_valid & core__ibuf_io_inst_0_bits_replay ; 
             core_mem_reg_xcpt_interrupt  <= core_take_pc_mem_wb ==1'h0& core_ex_reg_xcpt_interrupt ; 
             core_mem_reg_valid  <= core_ctrl_killx ==1'h0; 
             core_mem_reg_xcpt  <= core_ctrl_killx ==1'h0& core_ex_xcpt ; 
             core_mem_reg_replay  <= core_take_pc_mem_wb ==1'h0& core_replay_ex ; 
             core_wb_reg_valid  <= core_ctrl_killm ==1'h0; 
             core_wb_reg_xcpt  <= core_mem_xcpt & core_take_pc_wb ==1'h0; 
             core_wb_reg_replay  <= core_replay_mem & core_take_pc_wb ==1'h0; 
             core_wb_reg_flush_pipe  <= core_ctrl_killm ==1'h0& core_mem_reg_flush_pipe ; 
             core_div_io_kill_REG  <= core__div_io_req_ready & core__GEN_9 ; 
             core_dcache_blocked_blocked  <= core_io_dmem_req_ready ==1'h0& core_io_dmem_clock_enabled & core_io_dmem_perf_grant ==1'h0&( core_dcache_blocked_blocked | core__io_dmem_req_valid_output | core_io_dmem_s2_nack ); 
             core_rocc_blocked  <= core_wb_xcpt ==1'h0& core_io_rocc_cmd_ready ==1'h0&( core__io_rocc_cmd_valid_output | core_rocc_blocked ); 
             core_io_imem_progress_REG  <= core_wb_reg_valid & core_replay_wb_common ==1'h0; 
             core_icache_blocked_REG  <= core_io_imem_resp_valid ; 
             core_coreMonitorBundle_rd0val_REG  <= core_ex_rs_0 ; 
             core_coreMonitorBundle_rd0val_REG_1  <= core_coreMonitorBundle_rd0val_REG ; 
             core_coreMonitorBundle_rd1val_REG  <= core_ex_rs_1 ; 
             core_coreMonitorBundle_rd1val_REG_1  <= core_coreMonitorBundle_rd1val_REG ;
         end
  assign  core_io_imem_might_request = core_imem_might_request_reg ; 
  assign  core_io_imem_req_valid = core_take_pc_mem_wb ; 
  assign  core_io_imem_req_bits_pc = core__io_imem_req_bits_pc_output ; 
  assign  core_io_imem_req_bits_speculative = core_take_pc_wb ==1'h0; 
  assign  core_io_imem_sfence_valid = core__io_imem_sfence_valid_output ; 
  assign  core_io_imem_sfence_bits_rs1 = core__io_imem_sfence_bits_rs1_output ; 
  assign  core_io_imem_sfence_bits_rs2 = core__io_imem_sfence_bits_rs2_output ; 
  assign  core_io_imem_sfence_bits_addr = core__io_imem_sfence_bits_addr_output ; 
  assign  core_io_imem_sfence_bits_asid = core__io_imem_sfence_bits_asid_output ; 
  assign  core_io_imem_sfence_bits_hv = core__io_imem_sfence_bits_hv_output ; 
  assign  core_io_imem_sfence_bits_hg = core__io_imem_sfence_bits_hg_output ; 
  assign  core_io_imem_btb_update_valid = core_mem_reg_valid & core_take_pc_wb ==1'h0& core_mem_wrong_npc &( core_mem_cfi ==1'h0| core_mem_cfi_taken ); 
  assign  core_io_imem_btb_update_bits_prediction_cfiType = core_mem_reg_btb_resp_cfiType ; 
  assign  core_io_imem_btb_update_bits_prediction_taken = core_mem_reg_btb_resp_taken ; 
  assign  core_io_imem_btb_update_bits_prediction_mask = core_mem_reg_btb_resp_mask ; 
  assign  core_io_imem_btb_update_bits_prediction_bridx = core_mem_reg_btb_resp_bridx ; 
  assign  core_io_imem_btb_update_bits_prediction_target = core_mem_reg_btb_resp_target ; 
  assign  core_io_imem_btb_update_bits_prediction_entry = core_mem_reg_btb_resp_entry ; 
  assign  core_io_imem_btb_update_bits_prediction_bht_history = core_mem_reg_btb_resp_bht_history ; 
  assign  core_io_imem_btb_update_bits_prediction_bht_value = core_mem_reg_btb_resp_bht_value ; 
  assign  core_io_imem_btb_update_bits_pc = core__io_imem_btb_update_bits_pc_output ; 
  assign  core_io_imem_btb_update_bits_target = core__io_imem_req_bits_pc_output [32:0]; 
  assign  core_io_imem_btb_update_bits_taken =1'h0; 
  assign  core_io_imem_btb_update_bits_isValid = core_mem_cfi ; 
  assign  core_io_imem_btb_update_bits_br_pc = core__io_imem_btb_update_bits_br_pc_output ; 
  assign  core_io_imem_btb_update_bits_cfiType =( core_mem_ctrl_jal | core_mem_ctrl_jalr )& core_mem_waddr [0] ? 2'h2: core_mem_ctrl_jalr &5'h1==( core_mem_reg_inst [19:15]&5'h1B) ? 2'h3:{1'h0, core_mem_ctrl_jal | core_mem_ctrl_jalr }; 
  assign  core_io_imem_bht_update_valid = core_mem_reg_valid & core_take_pc_wb ==1'h0; 
  assign  core_io_imem_bht_update_bits_prediction_history = core_mem_reg_btb_resp_bht_history ; 
  assign  core_io_imem_bht_update_bits_prediction_value = core_mem_reg_btb_resp_bht_value ; 
  assign  core_io_imem_bht_update_bits_pc = core__io_imem_btb_update_bits_pc_output ; 
  assign  core_io_imem_bht_update_bits_branch = core_mem_ctrl_branch ; 
  assign  core_io_imem_bht_update_bits_taken = core_mem_br_taken ; 
  assign  core_io_imem_bht_update_bits_mispredict = core_mem_wrong_npc ; 
  assign  core_io_imem_ras_update_valid =1'h0; 
  assign  core_io_imem_ras_update_bits_cfiType =2'h0; 
  assign  core_io_imem_ras_update_bits_returnAddr =33'h0; 
  assign  core_io_imem_flush_icache = core_wb_reg_valid & core_wb_ctrl_fence_i & core_io_dmem_s2_nack ==1'h0; 
  assign  core_io_imem_progress = core_io_imem_progress_REG ; 
  assign  core_io_dmem_req_valid = core__io_dmem_req_valid_output ; 
  assign  core_io_dmem_req_bits_addr ={ core_io_dmem_req_bits_addr_msb , core__alu_io_adder_out [32:0]}; 
  assign  core_io_dmem_req_bits_tag = core_ex_dcache_tag ; 
  assign  core_io_dmem_req_bits_cmd = core_ex_ctrl_mem_cmd ; 
  assign  core_io_dmem_req_bits_size = core_ex_reg_mem_size ; 
  assign  core_io_dmem_req_bits_signed =( core_ex_reg_hls  ?  core_ex_reg_inst [20]: core_ex_reg_inst [14])==1'h0; 
  assign  core_io_dmem_req_bits_dprv = core_ex_reg_hls  ? {1'h0, core__csr_io_hstatus_spvp }: core__csr_io_status_dprv ; 
  assign  core_io_dmem_req_bits_dv = core__io_dmem_req_bits_dv_output ; 
  assign  core_io_dmem_req_bits_phys =1'h0; 
  assign  core_io_dmem_req_bits_no_alloc =1'h0; 
  assign  core_io_dmem_req_bits_no_xcpt =1'h0; 
  assign  core_io_dmem_req_bits_data =64'h0; 
  assign  core_io_dmem_req_bits_mask =8'h0; 
  assign  core_io_dmem_s1_kill = core_killm_common | core_mem_ldst_xcpt | core_fpu_kill_mem ; 
  assign  core_io_dmem_s1_data_data = core_mem_reg_rs2 ; 
  assign  core_io_dmem_s1_data_mask =8'h0; 
  assign  core_io_dmem_s2_kill =1'h0; 
  assign  core_io_dmem_keep_clock_enabled = core__ibuf_io_inst_0_valid & core_id_ctrl_mem & core__csr_io_csr_stall ==1'h0; 
  assign  core_io_ptw_sfence_valid = core__io_imem_sfence_valid_output ; 
  assign  core_io_ptw_sfence_bits_rs1 = core__io_imem_sfence_bits_rs1_output ; 
  assign  core_io_ptw_sfence_bits_rs2 = core__io_imem_sfence_bits_rs2_output ; 
  assign  core_io_ptw_sfence_bits_addr = core__io_imem_sfence_bits_addr_output ; 
  assign  core_io_ptw_sfence_bits_asid = core__io_imem_sfence_bits_asid_output ; 
  assign  core_io_ptw_sfence_bits_hv = core__io_imem_sfence_bits_hv_output ; 
  assign  core_io_ptw_sfence_bits_hg = core__io_imem_sfence_bits_hg_output ; 
  assign  core_io_ptw_status_debug = core__csr_io_status_debug ; 
  assign  core_io_ptw_status_cease = core__csr_io_status_cease ; 
  assign  core_io_ptw_status_wfi = core__csr_io_status_wfi ; 
  assign  core_io_ptw_status_isa = core__csr_io_status_isa ; 
  assign  core_io_ptw_status_dprv = core__csr_io_status_dprv ; 
  assign  core_io_ptw_status_dv = core__csr_io_status_dv ; 
  assign  core_io_ptw_status_prv = core__csr_io_status_prv ; 
  assign  core_io_ptw_status_v = core__csr_io_status_v ; 
  assign  core_io_ptw_status_sd = core__csr_io_status_sd ; 
  assign  core_io_ptw_status_zero2 = core__csr_io_status_zero2 ; 
  assign  core_io_ptw_status_mpv = core__csr_io_status_mpv ; 
  assign  core_io_ptw_status_gva = core__csr_io_status_gva ; 
  assign  core_io_ptw_status_mbe = core__csr_io_status_mbe ; 
  assign  core_io_ptw_status_sbe = core__csr_io_status_sbe ; 
  assign  core_io_ptw_status_sxl = core__csr_io_status_sxl ; 
  assign  core_io_ptw_status_uxl = core__csr_io_status_uxl ; 
  assign  core_io_ptw_status_sd_rv32 = core__csr_io_status_sd_rv32 ; 
  assign  core_io_ptw_status_zero1 = core__csr_io_status_zero1 ; 
  assign  core_io_ptw_status_tsr = core__csr_io_status_tsr ; 
  assign  core_io_ptw_status_tw = core__csr_io_status_tw ; 
  assign  core_io_ptw_status_tvm = core__csr_io_status_tvm ; 
  assign  core_io_ptw_status_mxr = core__csr_io_status_mxr ; 
  assign  core_io_ptw_status_sum = core__csr_io_status_sum ; 
  assign  core_io_ptw_status_mprv = core__csr_io_status_mprv ; 
  assign  core_io_ptw_status_xs = core__csr_io_status_xs ; 
  assign  core_io_ptw_status_fs = core__csr_io_status_fs ; 
  assign  core_io_ptw_status_mpp = core__csr_io_status_mpp ; 
  assign  core_io_ptw_status_vs = core__csr_io_status_vs ; 
  assign  core_io_ptw_status_spp = core__csr_io_status_spp ; 
  assign  core_io_ptw_status_mpie = core__csr_io_status_mpie ; 
  assign  core_io_ptw_status_ube = core__csr_io_status_ube ; 
  assign  core_io_ptw_status_spie = core__csr_io_status_spie ; 
  assign  core_io_ptw_status_upie = core__csr_io_status_upie ; 
  assign  core_io_ptw_status_mie = core__csr_io_status_mie ; 
  assign  core_io_ptw_status_hie = core__csr_io_status_hie ; 
  assign  core_io_ptw_status_sie = core__csr_io_status_sie ; 
  assign  core_io_ptw_status_uie = core__csr_io_status_uie ; 
  assign  core_io_ptw_hstatus_spvp = core__csr_io_hstatus_spvp ; 
  assign  core_io_ptw_customCSRs_csrs_0_value = core__io_ptw_customCSRs_csrs_0_value_output ; 
  assign  core_io_fpu_hartid = core_io_hartid ; 
  assign  core_io_fpu_time ={32'h0, core__csr_io_time [31:0]}; 
  assign  core_io_fpu_inst = core__ibuf_io_inst_0_bits_inst_bits ; 
  assign  core_io_fpu_fromint_data = core_ex_rs_0 ; 
  assign  core_io_fpu_dmem_resp_val = core_dmem_resp_valid & core_dmem_resp_fpu ; 
  assign  core_io_fpu_dmem_resp_type ={1'h0, core_io_dmem_resp_bits_size }; 
  assign  core_io_fpu_dmem_resp_tag = core_dmem_resp_waddr ; 
  assign  core_io_fpu_valid = core_ctrl_killd ==1'h0& core_id_ctrl_fp ; 
  assign  core_io_fpu_killx = core_ctrl_killx ; 
  assign  core_io_fpu_killm = core_killm_common ; 
  assign  core_io_fpu_keep_clock_enabled = core__io_ptw_customCSRs_csrs_0_value_output [2]; 
  assign  core_io_rocc_cmd_valid = core__io_rocc_cmd_valid_output ; 
  assign  core_io_rocc_cmd_bits_inst_funct = core__io_rocc_cmd_bits_inst_WIRE_funct ; 
  assign  core_io_rocc_cmd_bits_inst_rs2 = core__io_rocc_cmd_bits_inst_WIRE_rs2 ; 
  assign  core_io_rocc_cmd_bits_inst_rs1 = core__io_rocc_cmd_bits_inst_WIRE_rs1 ; 
  assign  core_io_rocc_cmd_bits_inst_xd = core__io_rocc_cmd_bits_inst_WIRE_xd ; 
  assign  core_io_rocc_cmd_bits_inst_xs1 = core__io_rocc_cmd_bits_inst_WIRE_xs1 ; 
  assign  core_io_rocc_cmd_bits_inst_xs2 = core__io_rocc_cmd_bits_inst_WIRE_xs2 ; 
  assign  core_io_rocc_cmd_bits_inst_rd = core__io_rocc_cmd_bits_inst_WIRE_rd ; 
  assign  core_io_rocc_cmd_bits_inst_opcode = core__io_rocc_cmd_bits_inst_WIRE_opcode ; 
  assign  core_io_rocc_cmd_bits_rs1 = core_wb_reg_wdata ; 
  assign  core_io_rocc_cmd_bits_rs2 = core_wb_reg_rs2 ; 
  assign  core_io_rocc_cmd_bits_status_debug = core__csr_io_status_debug ; 
  assign  core_io_rocc_cmd_bits_status_cease = core__csr_io_status_cease ; 
  assign  core_io_rocc_cmd_bits_status_wfi = core__csr_io_status_wfi ; 
  assign  core_io_rocc_cmd_bits_status_isa = core__csr_io_status_isa ; 
  assign  core_io_rocc_cmd_bits_status_dprv = core__csr_io_status_dprv ; 
  assign  core_io_rocc_cmd_bits_status_dv = core__csr_io_status_dv ; 
  assign  core_io_rocc_cmd_bits_status_prv = core__csr_io_status_prv ; 
  assign  core_io_rocc_cmd_bits_status_v = core__csr_io_status_v ; 
  assign  core_io_rocc_cmd_bits_status_sd = core__csr_io_status_sd ; 
  assign  core_io_rocc_cmd_bits_status_zero2 = core__csr_io_status_zero2 ; 
  assign  core_io_rocc_cmd_bits_status_mpv = core__csr_io_status_mpv ; 
  assign  core_io_rocc_cmd_bits_status_gva = core__csr_io_status_gva ; 
  assign  core_io_rocc_cmd_bits_status_mbe = core__csr_io_status_mbe ; 
  assign  core_io_rocc_cmd_bits_status_sbe = core__csr_io_status_sbe ; 
  assign  core_io_rocc_cmd_bits_status_sxl = core__csr_io_status_sxl ; 
  assign  core_io_rocc_cmd_bits_status_uxl = core__csr_io_status_uxl ; 
  assign  core_io_rocc_cmd_bits_status_sd_rv32 = core__csr_io_status_sd_rv32 ; 
  assign  core_io_rocc_cmd_bits_status_zero1 = core__csr_io_status_zero1 ; 
  assign  core_io_rocc_cmd_bits_status_tsr = core__csr_io_status_tsr ; 
  assign  core_io_rocc_cmd_bits_status_tw = core__csr_io_status_tw ; 
  assign  core_io_rocc_cmd_bits_status_tvm = core__csr_io_status_tvm ; 
  assign  core_io_rocc_cmd_bits_status_mxr = core__csr_io_status_mxr ; 
  assign  core_io_rocc_cmd_bits_status_sum = core__csr_io_status_sum ; 
  assign  core_io_rocc_cmd_bits_status_mprv = core__csr_io_status_mprv ; 
  assign  core_io_rocc_cmd_bits_status_xs = core__csr_io_status_xs ; 
  assign  core_io_rocc_cmd_bits_status_fs = core__csr_io_status_fs ; 
  assign  core_io_rocc_cmd_bits_status_mpp = core__csr_io_status_mpp ; 
  assign  core_io_rocc_cmd_bits_status_vs = core__csr_io_status_vs ; 
  assign  core_io_rocc_cmd_bits_status_spp = core__csr_io_status_spp ; 
  assign  core_io_rocc_cmd_bits_status_mpie = core__csr_io_status_mpie ; 
  assign  core_io_rocc_cmd_bits_status_ube = core__csr_io_status_ube ; 
  assign  core_io_rocc_cmd_bits_status_spie = core__csr_io_status_spie ; 
  assign  core_io_rocc_cmd_bits_status_upie = core__csr_io_status_upie ; 
  assign  core_io_rocc_cmd_bits_status_mie = core__csr_io_status_mie ; 
  assign  core_io_rocc_cmd_bits_status_hie = core__csr_io_status_hie ; 
  assign  core_io_rocc_cmd_bits_status_sie = core__csr_io_status_sie ; 
  assign  core_io_rocc_cmd_bits_status_uie = core__csr_io_status_uie ; 
  assign  core_io_rocc_resp_ready =1'h0; 
  assign  core_io_rocc_mem_req_ready =1'h0; 
  assign  core_io_rocc_mem_s2_nack =1'h0; 
  assign  core_io_rocc_mem_s2_nack_cause_raw =1'h0; 
  assign  core_io_rocc_mem_s2_uncached =1'h0; 
  assign  core_io_rocc_mem_s2_paddr =32'h0; 
  assign  core_io_rocc_mem_resp_valid =1'h0; 
  assign  core_io_rocc_mem_resp_bits_addr =34'h0; 
  assign  core_io_rocc_mem_resp_bits_tag =6'h0; 
  assign  core_io_rocc_mem_resp_bits_cmd =5'h0; 
  assign  core_io_rocc_mem_resp_bits_size =2'h0; 
  assign  core_io_rocc_mem_resp_bits_signed =1'h0; 
  assign  core_io_rocc_mem_resp_bits_dprv =2'h0; 
  assign  core_io_rocc_mem_resp_bits_dv =1'h0; 
  assign  core_io_rocc_mem_resp_bits_data =64'h0; 
  assign  core_io_rocc_mem_resp_bits_mask =8'h0; 
  assign  core_io_rocc_mem_resp_bits_replay =1'h0; 
  assign  core_io_rocc_mem_resp_bits_has_data =1'h0; 
  assign  core_io_rocc_mem_resp_bits_data_word_bypass =64'h0; 
  assign  core_io_rocc_mem_resp_bits_data_raw =64'h0; 
  assign  core_io_rocc_mem_resp_bits_store_data =64'h0; 
  assign  core_io_rocc_mem_replay_next =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_ma_ld =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_ma_st =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_pf_ld =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_pf_st =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_gf_ld =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_gf_st =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_ae_ld =1'h0; 
  assign  core_io_rocc_mem_s2_xcpt_ae_st =1'h0; 
  assign  core_io_rocc_mem_s2_gpa =34'h0; 
  assign  core_io_rocc_mem_s2_gpa_is_pte =1'h0; 
  assign  core_io_rocc_mem_ordered =1'h0; 
  assign  core_io_rocc_mem_perf_acquire =1'h0; 
  assign  core_io_rocc_mem_perf_release =1'h0; 
  assign  core_io_rocc_mem_perf_grant =1'h0; 
  assign  core_io_rocc_mem_perf_tlbMiss =1'h0; 
  assign  core_io_rocc_mem_perf_blocked =1'h0; 
  assign  core_io_rocc_mem_perf_canAcceptStoreThenLoad =1'h0; 
  assign  core_io_rocc_mem_perf_canAcceptStoreThenRMW =1'h0; 
  assign  core_io_rocc_mem_perf_canAcceptLoadThenLoad =1'h0; 
  assign  core_io_rocc_mem_perf_storeBufferEmptyAfterLoad =1'h0; 
  assign  core_io_rocc_mem_perf_storeBufferEmptyAfterStore =1'h0; 
  assign  core_io_rocc_mem_clock_enabled =1'h0; 
  assign  core_io_rocc_exception = core_wb_xcpt &(| core__csr_io_status_xs ); 
  assign  core_io_trace_insns_0_valid = core__csr_io_trace_0_valid ; 
  assign  core_io_trace_insns_0_iaddr = core__csr_io_trace_0_iaddr ; 
  assign  core_io_trace_insns_0_insn = core__csr_io_trace_0_insn ; 
  assign  core_io_trace_insns_0_priv = core__csr_io_trace_0_priv ; 
  assign  core_io_trace_insns_0_exception = core__csr_io_trace_0_exception ; 
  assign  core_io_trace_time = core__csr_io_time ; 
  assign  core_io_bpwatch_0_valid_0 = core_wb_reg_wphit_0 ; 
  assign  core_io_bpwatch_0_rvalid_0 =1'h0; 
  assign  core_io_bpwatch_0_wvalid_0 =1'h0; 
  assign  core_io_bpwatch_0_ivalid_0 =1'h0; 
  assign  core_io_bpwatch_0_action ={2'h0, core__csr_io_bp_0_control_action }; 
  assign  core_io_cease = core__csr_io_status_cease & core_clock_en_reg ==1'h0; 
  assign  core_io_wfi = core__csr_io_status_wfi ;
    assign core_clock = clock;
    assign core_reset = reset;
    assign core_io_hartid = hartIdSinkNodeIn;
    assign core_io_reset_vector = 32'h0;
    assign core_io_interrupts_debug = intSinkNodeIn_0;
    assign core_io_interrupts_mtip = intSinkNodeIn_2;
    assign core_io_interrupts_msip = intSinkNodeIn_1;
    assign core_io_interrupts_meip = intSinkNodeIn_3;
    assign _core_io_imem_might_request = core_io_imem_might_request;
    assign core_io_imem_clock_enabled = _frontend_io_cpu_clock_enabled;
    assign _core_io_imem_req_valid = core_io_imem_req_valid;
    assign _core_io_imem_req_bits_pc = core_io_imem_req_bits_pc;
    assign _core_io_imem_req_bits_speculative = core_io_imem_req_bits_speculative;
    assign _core_io_imem_sfence_valid = core_io_imem_sfence_valid;
    assign _core_io_imem_sfence_bits_rs1 = core_io_imem_sfence_bits_rs1;
    assign _core_io_imem_sfence_bits_rs2 = core_io_imem_sfence_bits_rs2;
    assign _core_io_imem_sfence_bits_addr = core_io_imem_sfence_bits_addr;
    assign _core_io_imem_sfence_bits_asid = core_io_imem_sfence_bits_asid;
    assign _core_io_imem_sfence_bits_hv = core_io_imem_sfence_bits_hv;
    assign _core_io_imem_sfence_bits_hg = core_io_imem_sfence_bits_hg;
    assign _core_io_imem_resp_ready = core_io_imem_resp_ready;
    assign core_io_imem_resp_valid = _frontend_io_cpu_resp_valid;
    assign core_io_imem_resp_bits_btb_cfiType = _frontend_io_cpu_resp_bits_btb_cfiType;
    assign core_io_imem_resp_bits_btb_taken = _frontend_io_cpu_resp_bits_btb_taken;
    assign core_io_imem_resp_bits_btb_mask = _frontend_io_cpu_resp_bits_btb_mask;
    assign core_io_imem_resp_bits_btb_bridx = _frontend_io_cpu_resp_bits_btb_bridx;
    assign core_io_imem_resp_bits_btb_target = _frontend_io_cpu_resp_bits_btb_target;
    assign core_io_imem_resp_bits_btb_entry = _frontend_io_cpu_resp_bits_btb_entry;
    assign core_io_imem_resp_bits_btb_bht_history = _frontend_io_cpu_resp_bits_btb_bht_history;
    assign core_io_imem_resp_bits_btb_bht_value = _frontend_io_cpu_resp_bits_btb_bht_value;
    assign core_io_imem_resp_bits_pc = _frontend_io_cpu_resp_bits_pc;
    assign core_io_imem_resp_bits_data = _frontend_io_cpu_resp_bits_data;
    assign core_io_imem_resp_bits_mask = _frontend_io_cpu_resp_bits_mask;
    assign core_io_imem_resp_bits_xcpt_pf_inst = _frontend_io_cpu_resp_bits_xcpt_pf_inst;
    assign core_io_imem_resp_bits_xcpt_gf_inst = _frontend_io_cpu_resp_bits_xcpt_gf_inst;
    assign core_io_imem_resp_bits_xcpt_ae_inst = _frontend_io_cpu_resp_bits_xcpt_ae_inst;
    assign core_io_imem_resp_bits_replay = _frontend_io_cpu_resp_bits_replay;
    assign core_io_imem_gpa_valid = _frontend_io_cpu_gpa_valid;
    assign core_io_imem_gpa_bits = _frontend_io_cpu_gpa_bits;
    assign _core_io_imem_btb_update_valid = core_io_imem_btb_update_valid;
    assign _core_io_imem_btb_update_bits_prediction_cfiType = core_io_imem_btb_update_bits_prediction_cfiType;
    assign _core_io_imem_btb_update_bits_prediction_taken = core_io_imem_btb_update_bits_prediction_taken;
    assign _core_io_imem_btb_update_bits_prediction_mask = core_io_imem_btb_update_bits_prediction_mask;
    assign _core_io_imem_btb_update_bits_prediction_bridx = core_io_imem_btb_update_bits_prediction_bridx;
    assign _core_io_imem_btb_update_bits_prediction_target = core_io_imem_btb_update_bits_prediction_target;
    assign _core_io_imem_btb_update_bits_prediction_entry = core_io_imem_btb_update_bits_prediction_entry;
    assign _core_io_imem_btb_update_bits_prediction_bht_history = core_io_imem_btb_update_bits_prediction_bht_history;
    assign _core_io_imem_btb_update_bits_prediction_bht_value = core_io_imem_btb_update_bits_prediction_bht_value;
    assign _core_io_imem_btb_update_bits_pc = core_io_imem_btb_update_bits_pc;
    assign _core_io_imem_btb_update_bits_target = core_io_imem_btb_update_bits_target;
    assign _core_io_imem_btb_update_bits_taken = core_io_imem_btb_update_bits_taken;
    assign _core_io_imem_btb_update_bits_isValid = core_io_imem_btb_update_bits_isValid;
    assign _core_io_imem_btb_update_bits_br_pc = core_io_imem_btb_update_bits_br_pc;
    assign _core_io_imem_btb_update_bits_cfiType = core_io_imem_btb_update_bits_cfiType;
    assign _core_io_imem_bht_update_valid = core_io_imem_bht_update_valid;
    assign _core_io_imem_bht_update_bits_prediction_history = core_io_imem_bht_update_bits_prediction_history;
    assign _core_io_imem_bht_update_bits_prediction_value = core_io_imem_bht_update_bits_prediction_value;
    assign _core_io_imem_bht_update_bits_pc = core_io_imem_bht_update_bits_pc;
    assign _core_io_imem_bht_update_bits_branch = core_io_imem_bht_update_bits_branch;
    assign _core_io_imem_bht_update_bits_taken = core_io_imem_bht_update_bits_taken;
    assign _core_io_imem_bht_update_bits_mispredict = core_io_imem_bht_update_bits_mispredict;
    assign _core_io_imem_ras_update_valid = core_io_imem_ras_update_valid;
    assign _core_io_imem_ras_update_bits_cfiType = core_io_imem_ras_update_bits_cfiType;
    assign _core_io_imem_ras_update_bits_returnAddr = core_io_imem_ras_update_bits_returnAddr;
    assign _core_io_imem_flush_icache = core_io_imem_flush_icache;
    assign core_io_imem_npc = _frontend_io_cpu_npc;
    assign core_io_imem_perf_acquire = _frontend_io_cpu_perf_acquire;
    assign core_io_imem_perf_tlbMiss = _frontend_io_cpu_perf_tlbMiss;
    assign _core_io_imem_progress = core_io_imem_progress;
    assign core_io_dmem_req_ready = _dcacheArb_io_requestor_0_req_ready;
    assign _core_io_dmem_req_valid = core_io_dmem_req_valid;
    assign _core_io_dmem_req_bits_addr = core_io_dmem_req_bits_addr;
    assign _core_io_dmem_req_bits_tag = core_io_dmem_req_bits_tag;
    assign _core_io_dmem_req_bits_cmd = core_io_dmem_req_bits_cmd;
    assign _core_io_dmem_req_bits_size = core_io_dmem_req_bits_size;
    assign _core_io_dmem_req_bits_signed = core_io_dmem_req_bits_signed;
    assign _core_io_dmem_req_bits_dprv = core_io_dmem_req_bits_dprv;
    assign _core_io_dmem_req_bits_dv = core_io_dmem_req_bits_dv;
    assign _core_io_dmem_req_bits_phys = core_io_dmem_req_bits_phys;
    assign _core_io_dmem_req_bits_no_alloc = core_io_dmem_req_bits_no_alloc;
    assign _core_io_dmem_req_bits_no_xcpt = core_io_dmem_req_bits_no_xcpt;
    assign _core_io_dmem_req_bits_data = core_io_dmem_req_bits_data;
    assign _core_io_dmem_req_bits_mask = core_io_dmem_req_bits_mask;
    assign _core_io_dmem_s1_kill = core_io_dmem_s1_kill;
    assign _core_io_dmem_s1_data_data = core_io_dmem_s1_data_data;
    assign _core_io_dmem_s1_data_mask = core_io_dmem_s1_data_mask;
    assign core_io_dmem_s2_nack = _dcacheArb_io_requestor_0_s2_nack;
    assign core_io_dmem_s2_nack_cause_raw = _dcacheArb_io_requestor_0_s2_nack_cause_raw;
    assign _core_io_dmem_s2_kill = core_io_dmem_s2_kill;
    assign core_io_dmem_s2_uncached = _dcacheArb_io_requestor_0_s2_uncached;
    assign core_io_dmem_s2_paddr = _dcacheArb_io_requestor_0_s2_paddr;
    assign core_io_dmem_resp_valid = _dcacheArb_io_requestor_0_resp_valid;
    assign core_io_dmem_resp_bits_addr = _dcacheArb_io_requestor_0_resp_bits_addr;
    assign core_io_dmem_resp_bits_tag = _dcacheArb_io_requestor_0_resp_bits_tag;
    assign core_io_dmem_resp_bits_cmd = _dcacheArb_io_requestor_0_resp_bits_cmd;
    assign core_io_dmem_resp_bits_size = _dcacheArb_io_requestor_0_resp_bits_size;
    assign core_io_dmem_resp_bits_signed = _dcacheArb_io_requestor_0_resp_bits_signed;
    assign core_io_dmem_resp_bits_dprv = _dcacheArb_io_requestor_0_resp_bits_dprv;
    assign core_io_dmem_resp_bits_dv = _dcacheArb_io_requestor_0_resp_bits_dv;
    assign core_io_dmem_resp_bits_data = _dcacheArb_io_requestor_0_resp_bits_data;
    assign core_io_dmem_resp_bits_mask = _dcacheArb_io_requestor_0_resp_bits_mask;
    assign core_io_dmem_resp_bits_replay = _dcacheArb_io_requestor_0_resp_bits_replay;
    assign core_io_dmem_resp_bits_has_data = _dcacheArb_io_requestor_0_resp_bits_has_data;
    assign core_io_dmem_resp_bits_data_word_bypass = _dcacheArb_io_requestor_0_resp_bits_data_word_bypass;
    assign core_io_dmem_resp_bits_data_raw = _dcacheArb_io_requestor_0_resp_bits_data_raw;
    assign core_io_dmem_resp_bits_store_data = _dcacheArb_io_requestor_0_resp_bits_store_data;
    assign core_io_dmem_replay_next = _dcacheArb_io_requestor_0_replay_next;
    assign core_io_dmem_s2_xcpt_ma_ld = _dcacheArb_io_requestor_0_s2_xcpt_ma_ld;
    assign core_io_dmem_s2_xcpt_ma_st = _dcacheArb_io_requestor_0_s2_xcpt_ma_st;
    assign core_io_dmem_s2_xcpt_pf_ld = _dcacheArb_io_requestor_0_s2_xcpt_pf_ld;
    assign core_io_dmem_s2_xcpt_pf_st = _dcacheArb_io_requestor_0_s2_xcpt_pf_st;
    assign core_io_dmem_s2_xcpt_gf_ld = _dcacheArb_io_requestor_0_s2_xcpt_gf_ld;
    assign core_io_dmem_s2_xcpt_gf_st = _dcacheArb_io_requestor_0_s2_xcpt_gf_st;
    assign core_io_dmem_s2_xcpt_ae_ld = _dcacheArb_io_requestor_0_s2_xcpt_ae_ld;
    assign core_io_dmem_s2_xcpt_ae_st = _dcacheArb_io_requestor_0_s2_xcpt_ae_st;
    assign core_io_dmem_s2_gpa = _dcacheArb_io_requestor_0_s2_gpa;
    assign core_io_dmem_s2_gpa_is_pte = _dcacheArb_io_requestor_0_s2_gpa_is_pte;
    assign core_io_dmem_ordered = _dcacheArb_io_requestor_0_ordered;
    assign core_io_dmem_perf_acquire = _dcacheArb_io_requestor_0_perf_acquire;
    assign core_io_dmem_perf_release = _dcacheArb_io_requestor_0_perf_release;
    assign core_io_dmem_perf_grant = _dcacheArb_io_requestor_0_perf_grant;
    assign core_io_dmem_perf_tlbMiss = _dcacheArb_io_requestor_0_perf_tlbMiss;
    assign core_io_dmem_perf_blocked = _dcacheArb_io_requestor_0_perf_blocked;
    assign core_io_dmem_perf_canAcceptStoreThenLoad = _dcacheArb_io_requestor_0_perf_canAcceptStoreThenLoad;
    assign core_io_dmem_perf_canAcceptStoreThenRMW = _dcacheArb_io_requestor_0_perf_canAcceptStoreThenRMW;
    assign core_io_dmem_perf_canAcceptLoadThenLoad = _dcacheArb_io_requestor_0_perf_canAcceptLoadThenLoad;
    assign core_io_dmem_perf_storeBufferEmptyAfterLoad = _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterLoad;
    assign core_io_dmem_perf_storeBufferEmptyAfterStore = _dcacheArb_io_requestor_0_perf_storeBufferEmptyAfterStore;
    assign _core_io_dmem_keep_clock_enabled = core_io_dmem_keep_clock_enabled;
    assign core_io_dmem_clock_enabled = _dcacheArb_io_requestor_0_clock_enabled;
    assign _core_io_ptw_ptbr_mode = core_io_ptw_ptbr_mode;
    assign _core_io_ptw_ptbr_asid = core_io_ptw_ptbr_asid;
    assign _core_io_ptw_ptbr_ppn = core_io_ptw_ptbr_ppn;
    assign _core_io_ptw_hgatp_mode = core_io_ptw_hgatp_mode;
    assign _core_io_ptw_hgatp_asid = core_io_ptw_hgatp_asid;
    assign _core_io_ptw_hgatp_ppn = core_io_ptw_hgatp_ppn;
    assign _core_io_ptw_vsatp_mode = core_io_ptw_vsatp_mode;
    assign _core_io_ptw_vsatp_asid = core_io_ptw_vsatp_asid;
    assign _core_io_ptw_vsatp_ppn = core_io_ptw_vsatp_ppn;
    assign _core_io_ptw_sfence_valid = core_io_ptw_sfence_valid;
    assign _core_io_ptw_sfence_bits_rs1 = core_io_ptw_sfence_bits_rs1;
    assign _core_io_ptw_sfence_bits_rs2 = core_io_ptw_sfence_bits_rs2;
    assign _core_io_ptw_sfence_bits_addr = core_io_ptw_sfence_bits_addr;
    assign _core_io_ptw_sfence_bits_asid = core_io_ptw_sfence_bits_asid;
    assign _core_io_ptw_sfence_bits_hv = core_io_ptw_sfence_bits_hv;
    assign _core_io_ptw_sfence_bits_hg = core_io_ptw_sfence_bits_hg;
    assign _core_io_ptw_status_debug = core_io_ptw_status_debug;
    assign _core_io_ptw_status_cease = core_io_ptw_status_cease;
    assign _core_io_ptw_status_wfi = core_io_ptw_status_wfi;
    assign _core_io_ptw_status_isa = core_io_ptw_status_isa;
    assign _core_io_ptw_status_dprv = core_io_ptw_status_dprv;
    assign _core_io_ptw_status_dv = core_io_ptw_status_dv;
    assign _core_io_ptw_status_prv = core_io_ptw_status_prv;
    assign _core_io_ptw_status_v = core_io_ptw_status_v;
    assign _core_io_ptw_status_sd = core_io_ptw_status_sd;
    assign _core_io_ptw_status_zero2 = core_io_ptw_status_zero2;
    assign _core_io_ptw_status_mpv = core_io_ptw_status_mpv;
    assign _core_io_ptw_status_gva = core_io_ptw_status_gva;
    assign _core_io_ptw_status_mbe = core_io_ptw_status_mbe;
    assign _core_io_ptw_status_sbe = core_io_ptw_status_sbe;
    assign _core_io_ptw_status_sxl = core_io_ptw_status_sxl;
    assign _core_io_ptw_status_uxl = core_io_ptw_status_uxl;
    assign _core_io_ptw_status_sd_rv32 = core_io_ptw_status_sd_rv32;
    assign _core_io_ptw_status_zero1 = core_io_ptw_status_zero1;
    assign _core_io_ptw_status_tsr = core_io_ptw_status_tsr;
    assign _core_io_ptw_status_tw = core_io_ptw_status_tw;
    assign _core_io_ptw_status_tvm = core_io_ptw_status_tvm;
    assign _core_io_ptw_status_mxr = core_io_ptw_status_mxr;
    assign _core_io_ptw_status_sum = core_io_ptw_status_sum;
    assign _core_io_ptw_status_mprv = core_io_ptw_status_mprv;
    assign _core_io_ptw_status_xs = core_io_ptw_status_xs;
    assign _core_io_ptw_status_fs = core_io_ptw_status_fs;
    assign _core_io_ptw_status_mpp = core_io_ptw_status_mpp;
    assign _core_io_ptw_status_vs = core_io_ptw_status_vs;
    assign _core_io_ptw_status_spp = core_io_ptw_status_spp;
    assign _core_io_ptw_status_mpie = core_io_ptw_status_mpie;
    assign _core_io_ptw_status_ube = core_io_ptw_status_ube;
    assign _core_io_ptw_status_spie = core_io_ptw_status_spie;
    assign _core_io_ptw_status_upie = core_io_ptw_status_upie;
    assign _core_io_ptw_status_mie = core_io_ptw_status_mie;
    assign _core_io_ptw_status_hie = core_io_ptw_status_hie;
    assign _core_io_ptw_status_sie = core_io_ptw_status_sie;
    assign _core_io_ptw_status_uie = core_io_ptw_status_uie;
    assign _core_io_ptw_hstatus_zero6 = core_io_ptw_hstatus_zero6;
    assign _core_io_ptw_hstatus_vsxl = core_io_ptw_hstatus_vsxl;
    assign _core_io_ptw_hstatus_zero5 = core_io_ptw_hstatus_zero5;
    assign _core_io_ptw_hstatus_vtsr = core_io_ptw_hstatus_vtsr;
    assign _core_io_ptw_hstatus_vtw = core_io_ptw_hstatus_vtw;
    assign _core_io_ptw_hstatus_vtvm = core_io_ptw_hstatus_vtvm;
    assign _core_io_ptw_hstatus_zero3 = core_io_ptw_hstatus_zero3;
    assign _core_io_ptw_hstatus_vgein = core_io_ptw_hstatus_vgein;
    assign _core_io_ptw_hstatus_zero2 = core_io_ptw_hstatus_zero2;
    assign _core_io_ptw_hstatus_hu = core_io_ptw_hstatus_hu;
    assign _core_io_ptw_hstatus_spvp = core_io_ptw_hstatus_spvp;
    assign _core_io_ptw_hstatus_spv = core_io_ptw_hstatus_spv;
    assign _core_io_ptw_hstatus_gva = core_io_ptw_hstatus_gva;
    assign _core_io_ptw_hstatus_vsbe = core_io_ptw_hstatus_vsbe;
    assign _core_io_ptw_hstatus_zero1 = core_io_ptw_hstatus_zero1;
    assign _core_io_ptw_gstatus_debug = core_io_ptw_gstatus_debug;
    assign _core_io_ptw_gstatus_cease = core_io_ptw_gstatus_cease;
    assign _core_io_ptw_gstatus_wfi = core_io_ptw_gstatus_wfi;
    assign _core_io_ptw_gstatus_isa = core_io_ptw_gstatus_isa;
    assign _core_io_ptw_gstatus_dprv = core_io_ptw_gstatus_dprv;
    assign _core_io_ptw_gstatus_dv = core_io_ptw_gstatus_dv;
    assign _core_io_ptw_gstatus_prv = core_io_ptw_gstatus_prv;
    assign _core_io_ptw_gstatus_v = core_io_ptw_gstatus_v;
    assign _core_io_ptw_gstatus_sd = core_io_ptw_gstatus_sd;
    assign _core_io_ptw_gstatus_zero2 = core_io_ptw_gstatus_zero2;
    assign _core_io_ptw_gstatus_mpv = core_io_ptw_gstatus_mpv;
    assign _core_io_ptw_gstatus_gva = core_io_ptw_gstatus_gva;
    assign _core_io_ptw_gstatus_mbe = core_io_ptw_gstatus_mbe;
    assign _core_io_ptw_gstatus_sbe = core_io_ptw_gstatus_sbe;
    assign _core_io_ptw_gstatus_sxl = core_io_ptw_gstatus_sxl;
    assign _core_io_ptw_gstatus_uxl = core_io_ptw_gstatus_uxl;
    assign _core_io_ptw_gstatus_sd_rv32 = core_io_ptw_gstatus_sd_rv32;
    assign _core_io_ptw_gstatus_zero1 = core_io_ptw_gstatus_zero1;
    assign _core_io_ptw_gstatus_tsr = core_io_ptw_gstatus_tsr;
    assign _core_io_ptw_gstatus_tw = core_io_ptw_gstatus_tw;
    assign _core_io_ptw_gstatus_tvm = core_io_ptw_gstatus_tvm;
    assign _core_io_ptw_gstatus_mxr = core_io_ptw_gstatus_mxr;
    assign _core_io_ptw_gstatus_sum = core_io_ptw_gstatus_sum;
    assign _core_io_ptw_gstatus_mprv = core_io_ptw_gstatus_mprv;
    assign _core_io_ptw_gstatus_xs = core_io_ptw_gstatus_xs;
    assign _core_io_ptw_gstatus_fs = core_io_ptw_gstatus_fs;
    assign _core_io_ptw_gstatus_mpp = core_io_ptw_gstatus_mpp;
    assign _core_io_ptw_gstatus_vs = core_io_ptw_gstatus_vs;
    assign _core_io_ptw_gstatus_spp = core_io_ptw_gstatus_spp;
    assign _core_io_ptw_gstatus_mpie = core_io_ptw_gstatus_mpie;
    assign _core_io_ptw_gstatus_ube = core_io_ptw_gstatus_ube;
    assign _core_io_ptw_gstatus_spie = core_io_ptw_gstatus_spie;
    assign _core_io_ptw_gstatus_upie = core_io_ptw_gstatus_upie;
    assign _core_io_ptw_gstatus_mie = core_io_ptw_gstatus_mie;
    assign _core_io_ptw_gstatus_hie = core_io_ptw_gstatus_hie;
    assign _core_io_ptw_gstatus_sie = core_io_ptw_gstatus_sie;
    assign _core_io_ptw_gstatus_uie = core_io_ptw_gstatus_uie;
    assign _core_io_ptw_pmp_0_cfg_l = core_io_ptw_pmp_0_cfg_l;
    assign _core_io_ptw_pmp_0_cfg_res = core_io_ptw_pmp_0_cfg_res;
    assign _core_io_ptw_pmp_0_cfg_a = core_io_ptw_pmp_0_cfg_a;
    assign _core_io_ptw_pmp_0_cfg_x = core_io_ptw_pmp_0_cfg_x;
    assign _core_io_ptw_pmp_0_cfg_w = core_io_ptw_pmp_0_cfg_w;
    assign _core_io_ptw_pmp_0_cfg_r = core_io_ptw_pmp_0_cfg_r;
    assign _core_io_ptw_pmp_0_addr = core_io_ptw_pmp_0_addr;
    assign _core_io_ptw_pmp_0_mask = core_io_ptw_pmp_0_mask;
    assign _core_io_ptw_pmp_1_cfg_l = core_io_ptw_pmp_1_cfg_l;
    assign _core_io_ptw_pmp_1_cfg_res = core_io_ptw_pmp_1_cfg_res;
    assign _core_io_ptw_pmp_1_cfg_a = core_io_ptw_pmp_1_cfg_a;
    assign _core_io_ptw_pmp_1_cfg_x = core_io_ptw_pmp_1_cfg_x;
    assign _core_io_ptw_pmp_1_cfg_w = core_io_ptw_pmp_1_cfg_w;
    assign _core_io_ptw_pmp_1_cfg_r = core_io_ptw_pmp_1_cfg_r;
    assign _core_io_ptw_pmp_1_addr = core_io_ptw_pmp_1_addr;
    assign _core_io_ptw_pmp_1_mask = core_io_ptw_pmp_1_mask;
    assign _core_io_ptw_pmp_2_cfg_l = core_io_ptw_pmp_2_cfg_l;
    assign _core_io_ptw_pmp_2_cfg_res = core_io_ptw_pmp_2_cfg_res;
    assign _core_io_ptw_pmp_2_cfg_a = core_io_ptw_pmp_2_cfg_a;
    assign _core_io_ptw_pmp_2_cfg_x = core_io_ptw_pmp_2_cfg_x;
    assign _core_io_ptw_pmp_2_cfg_w = core_io_ptw_pmp_2_cfg_w;
    assign _core_io_ptw_pmp_2_cfg_r = core_io_ptw_pmp_2_cfg_r;
    assign _core_io_ptw_pmp_2_addr = core_io_ptw_pmp_2_addr;
    assign _core_io_ptw_pmp_2_mask = core_io_ptw_pmp_2_mask;
    assign _core_io_ptw_pmp_3_cfg_l = core_io_ptw_pmp_3_cfg_l;
    assign _core_io_ptw_pmp_3_cfg_res = core_io_ptw_pmp_3_cfg_res;
    assign _core_io_ptw_pmp_3_cfg_a = core_io_ptw_pmp_3_cfg_a;
    assign _core_io_ptw_pmp_3_cfg_x = core_io_ptw_pmp_3_cfg_x;
    assign _core_io_ptw_pmp_3_cfg_w = core_io_ptw_pmp_3_cfg_w;
    assign _core_io_ptw_pmp_3_cfg_r = core_io_ptw_pmp_3_cfg_r;
    assign _core_io_ptw_pmp_3_addr = core_io_ptw_pmp_3_addr;
    assign _core_io_ptw_pmp_3_mask = core_io_ptw_pmp_3_mask;
    assign _core_io_ptw_pmp_4_cfg_l = core_io_ptw_pmp_4_cfg_l;
    assign _core_io_ptw_pmp_4_cfg_res = core_io_ptw_pmp_4_cfg_res;
    assign _core_io_ptw_pmp_4_cfg_a = core_io_ptw_pmp_4_cfg_a;
    assign _core_io_ptw_pmp_4_cfg_x = core_io_ptw_pmp_4_cfg_x;
    assign _core_io_ptw_pmp_4_cfg_w = core_io_ptw_pmp_4_cfg_w;
    assign _core_io_ptw_pmp_4_cfg_r = core_io_ptw_pmp_4_cfg_r;
    assign _core_io_ptw_pmp_4_addr = core_io_ptw_pmp_4_addr;
    assign _core_io_ptw_pmp_4_mask = core_io_ptw_pmp_4_mask;
    assign _core_io_ptw_pmp_5_cfg_l = core_io_ptw_pmp_5_cfg_l;
    assign _core_io_ptw_pmp_5_cfg_res = core_io_ptw_pmp_5_cfg_res;
    assign _core_io_ptw_pmp_5_cfg_a = core_io_ptw_pmp_5_cfg_a;
    assign _core_io_ptw_pmp_5_cfg_x = core_io_ptw_pmp_5_cfg_x;
    assign _core_io_ptw_pmp_5_cfg_w = core_io_ptw_pmp_5_cfg_w;
    assign _core_io_ptw_pmp_5_cfg_r = core_io_ptw_pmp_5_cfg_r;
    assign _core_io_ptw_pmp_5_addr = core_io_ptw_pmp_5_addr;
    assign _core_io_ptw_pmp_5_mask = core_io_ptw_pmp_5_mask;
    assign _core_io_ptw_pmp_6_cfg_l = core_io_ptw_pmp_6_cfg_l;
    assign _core_io_ptw_pmp_6_cfg_res = core_io_ptw_pmp_6_cfg_res;
    assign _core_io_ptw_pmp_6_cfg_a = core_io_ptw_pmp_6_cfg_a;
    assign _core_io_ptw_pmp_6_cfg_x = core_io_ptw_pmp_6_cfg_x;
    assign _core_io_ptw_pmp_6_cfg_w = core_io_ptw_pmp_6_cfg_w;
    assign _core_io_ptw_pmp_6_cfg_r = core_io_ptw_pmp_6_cfg_r;
    assign _core_io_ptw_pmp_6_addr = core_io_ptw_pmp_6_addr;
    assign _core_io_ptw_pmp_6_mask = core_io_ptw_pmp_6_mask;
    assign _core_io_ptw_pmp_7_cfg_l = core_io_ptw_pmp_7_cfg_l;
    assign _core_io_ptw_pmp_7_cfg_res = core_io_ptw_pmp_7_cfg_res;
    assign _core_io_ptw_pmp_7_cfg_a = core_io_ptw_pmp_7_cfg_a;
    assign _core_io_ptw_pmp_7_cfg_x = core_io_ptw_pmp_7_cfg_x;
    assign _core_io_ptw_pmp_7_cfg_w = core_io_ptw_pmp_7_cfg_w;
    assign _core_io_ptw_pmp_7_cfg_r = core_io_ptw_pmp_7_cfg_r;
    assign _core_io_ptw_pmp_7_addr = core_io_ptw_pmp_7_addr;
    assign _core_io_ptw_pmp_7_mask = core_io_ptw_pmp_7_mask;
    assign core_io_ptw_perf_l2miss = _ptw_io_dpath_perf_l2miss;
    assign core_io_ptw_perf_l2hit = _ptw_io_dpath_perf_l2hit;
    assign core_io_ptw_perf_pte_miss = _ptw_io_dpath_perf_pte_miss;
    assign core_io_ptw_perf_pte_hit = _ptw_io_dpath_perf_pte_hit;
    assign _core_io_ptw_customCSRs_csrs_0_ren = core_io_ptw_customCSRs_csrs_0_ren;
    assign _core_io_ptw_customCSRs_csrs_0_wen = core_io_ptw_customCSRs_csrs_0_wen;
    assign _core_io_ptw_customCSRs_csrs_0_wdata = core_io_ptw_customCSRs_csrs_0_wdata;
    assign _core_io_ptw_customCSRs_csrs_0_value = core_io_ptw_customCSRs_csrs_0_value;
    assign core_io_ptw_customCSRs_csrs_0_stall = _ptw_io_dpath_customCSRs_csrs_0_stall;
    assign core_io_ptw_customCSRs_csrs_0_set = _ptw_io_dpath_customCSRs_csrs_0_set;
    assign core_io_ptw_customCSRs_csrs_0_sdata = _ptw_io_dpath_customCSRs_csrs_0_sdata;
    assign _core_io_ptw_customCSRs_csrs_1_ren = core_io_ptw_customCSRs_csrs_1_ren;
    assign _core_io_ptw_customCSRs_csrs_1_wen = core_io_ptw_customCSRs_csrs_1_wen;
    assign _core_io_ptw_customCSRs_csrs_1_wdata = core_io_ptw_customCSRs_csrs_1_wdata;
    assign _core_io_ptw_customCSRs_csrs_1_value = core_io_ptw_customCSRs_csrs_1_value;
    assign core_io_ptw_customCSRs_csrs_1_stall = _ptw_io_dpath_customCSRs_csrs_1_stall;
    assign core_io_ptw_customCSRs_csrs_1_set = _ptw_io_dpath_customCSRs_csrs_1_set;
    assign core_io_ptw_customCSRs_csrs_1_sdata = _ptw_io_dpath_customCSRs_csrs_1_sdata;
    assign _core_io_ptw_customCSRs_csrs_2_ren = core_io_ptw_customCSRs_csrs_2_ren;
    assign _core_io_ptw_customCSRs_csrs_2_wen = core_io_ptw_customCSRs_csrs_2_wen;
    assign _core_io_ptw_customCSRs_csrs_2_wdata = core_io_ptw_customCSRs_csrs_2_wdata;
    assign _core_io_ptw_customCSRs_csrs_2_value = core_io_ptw_customCSRs_csrs_2_value;
    assign core_io_ptw_customCSRs_csrs_2_stall = _ptw_io_dpath_customCSRs_csrs_2_stall;
    assign core_io_ptw_customCSRs_csrs_2_set = _ptw_io_dpath_customCSRs_csrs_2_set;
    assign core_io_ptw_customCSRs_csrs_2_sdata = _ptw_io_dpath_customCSRs_csrs_2_sdata;
    assign _core_io_ptw_customCSRs_csrs_3_ren = core_io_ptw_customCSRs_csrs_3_ren;
    assign _core_io_ptw_customCSRs_csrs_3_wen = core_io_ptw_customCSRs_csrs_3_wen;
    assign _core_io_ptw_customCSRs_csrs_3_wdata = core_io_ptw_customCSRs_csrs_3_wdata;
    assign _core_io_ptw_customCSRs_csrs_3_value = core_io_ptw_customCSRs_csrs_3_value;
    assign core_io_ptw_customCSRs_csrs_3_stall = _ptw_io_dpath_customCSRs_csrs_3_stall;
    assign core_io_ptw_customCSRs_csrs_3_set = _ptw_io_dpath_customCSRs_csrs_3_set;
    assign core_io_ptw_customCSRs_csrs_3_sdata = _ptw_io_dpath_customCSRs_csrs_3_sdata;
    assign core_io_ptw_clock_enabled = _ptw_io_dpath_clock_enabled;
    assign core_io_fpu_fcsr_flags_valid = 1'h0;
    assign core_io_fpu_fcsr_flags_bits = 5'h0;
    assign core_io_fpu_toint_data = 64'h0;
    assign core_io_fpu_fcsr_rdy = 1'h0;
    assign core_io_fpu_nack_mem = 1'h0;
    assign core_io_fpu_illegal_rm = 1'h0;
    assign core_io_fpu_dec_ldst = 1'h0;
    assign core_io_fpu_dec_wen = 1'h0;
    assign core_io_fpu_dec_ren1 = 1'h0;
    assign core_io_fpu_dec_ren2 = 1'h0;
    assign core_io_fpu_dec_ren3 = 1'h0;
    assign core_io_fpu_dec_swap12 = 1'h0;
    assign core_io_fpu_dec_swap23 = 1'h0;
    assign core_io_fpu_dec_typeTagIn = 2'h0;
    assign core_io_fpu_dec_typeTagOut = 2'h0;
    assign core_io_fpu_dec_fromint = 1'h0;
    assign core_io_fpu_dec_toint = 1'h0;
    assign core_io_fpu_dec_fastpipe = 1'h0;
    assign core_io_fpu_dec_fma = 1'h0;
    assign core_io_fpu_dec_div = 1'h0;
    assign core_io_fpu_dec_sqrt = 1'h0;
    assign core_io_fpu_dec_wflags = 1'h0;
    assign core_io_fpu_sboard_set = 1'h0;
    assign core_io_fpu_sboard_clr = 1'h0;
    assign core_io_fpu_sboard_clra = 5'h0;
    assign core_io_rocc_cmd_ready = 1'h0;
    assign core_io_rocc_resp_valid = 1'h0;
    assign core_io_rocc_resp_bits_rd = 5'h0;
    assign core_io_rocc_resp_bits_data = 64'h0;
    assign core_io_rocc_mem_req_valid = 1'h0;
    assign core_io_rocc_mem_req_bits_addr = 34'h0;
    assign core_io_rocc_mem_req_bits_tag = 6'h0;
    assign core_io_rocc_mem_req_bits_cmd = 5'h0;
    assign core_io_rocc_mem_req_bits_size = 2'h0;
    assign core_io_rocc_mem_req_bits_signed = 1'h0;
    assign core_io_rocc_mem_req_bits_dprv = 2'h0;
    assign core_io_rocc_mem_req_bits_dv = 1'h0;
    assign core_io_rocc_mem_req_bits_phys = 1'h0;
    assign core_io_rocc_mem_req_bits_no_alloc = 1'h0;
    assign core_io_rocc_mem_req_bits_no_xcpt = 1'h0;
    assign core_io_rocc_mem_req_bits_data = 64'h0;
    assign core_io_rocc_mem_req_bits_mask = 8'h0;
    assign core_io_rocc_mem_s1_kill = 1'h0;
    assign core_io_rocc_mem_s1_data_data = 64'h0;
    assign core_io_rocc_mem_s1_data_mask = 8'h0;
    assign core_io_rocc_mem_s2_kill = 1'h0;
    assign core_io_rocc_mem_keep_clock_enabled = 1'h0;
    assign core_io_rocc_busy = 1'h0;
    assign core_io_rocc_interrupt = 1'h0;
    assign traceSourceNodeOut_insns_0_valid = core_io_trace_insns_0_valid;
    assign traceSourceNodeOut_insns_0_iaddr = core_io_trace_insns_0_iaddr;
    assign traceSourceNodeOut_insns_0_insn = core_io_trace_insns_0_insn;
    assign traceSourceNodeOut_insns_0_priv = core_io_trace_insns_0_priv;
    assign traceSourceNodeOut_insns_0_exception = core_io_trace_insns_0_exception;
    assign traceSourceNodeOut_insns_0_interrupt = core_io_trace_insns_0_interrupt;
    assign traceSourceNodeOut_insns_0_cause = core_io_trace_insns_0_cause;
    assign traceSourceNodeOut_insns_0_tval = core_io_trace_insns_0_tval;
    assign traceSourceNodeOut_time = core_io_trace_time;
    assign bpwatchSourceNodeOut_0_valid_0 = core_io_bpwatch_0_valid_0;
    assign bpwatchSourceNodeOut_0_rvalid_0 = core_io_bpwatch_0_rvalid_0;
    assign bpwatchSourceNodeOut_0_wvalid_0 = core_io_bpwatch_0_wvalid_0;
    assign bpwatchSourceNodeOut_0_ivalid_0 = core_io_bpwatch_0_ivalid_0;
    assign bpwatchSourceNodeOut_0_action = core_io_bpwatch_0_action;
    assign _core_io_wfi = core_io_wfi;
    assign core_io_traceStall = traceAuxSinkNodeIn_stall;
    
  reg         wfiNodeOut_0_REG;	// src/main/scala/tile/Interrupts.scala:126:36
  wire        wfiNodeOut_0 = wfiNodeOut_0_REG;	// src/main/scala/diplomacy/Nodes.scala:1205:17, src/main/scala/tile/Interrupts.scala:126:36
  always @(posedge clock) begin
    if (reset)
      wfiNodeOut_0_REG <= 1'h0;	// src/main/scala/tile/BaseTile.scala:295:16, src/main/scala/tile/Interrupts.scala:126:36
    else
      wfiNodeOut_0_REG <= _core_io_wfi;	// src/main/scala/tile/Interrupts.scala:126:36, src/main/scala/tile/RocketTile.scala:127:20
  end // always @(posedge)
  assign auto_buffer_out_a_valid = buffer_auto_out_a_valid;
  assign auto_buffer_out_a_bits_opcode = buffer_auto_out_a_bits_opcode;
  assign auto_buffer_out_a_bits_param = buffer_auto_out_a_bits_param;
  assign auto_buffer_out_a_bits_size = buffer_auto_out_a_bits_size;
  assign auto_buffer_out_a_bits_source = buffer_auto_out_a_bits_source;
  assign auto_buffer_out_a_bits_address = buffer_auto_out_a_bits_address;
  assign auto_buffer_out_a_bits_user_amba_prot_bufferable =
    buffer_auto_out_a_bits_user_amba_prot_bufferable;
  assign auto_buffer_out_a_bits_user_amba_prot_modifiable =
    buffer_auto_out_a_bits_user_amba_prot_modifiable;
  assign auto_buffer_out_a_bits_user_amba_prot_readalloc =
    buffer_auto_out_a_bits_user_amba_prot_readalloc;
  assign auto_buffer_out_a_bits_user_amba_prot_writealloc =
    buffer_auto_out_a_bits_user_amba_prot_writealloc;
  assign auto_buffer_out_a_bits_user_amba_prot_privileged =
    buffer_auto_out_a_bits_user_amba_prot_privileged;
  assign auto_buffer_out_a_bits_user_amba_prot_secure =
    buffer_auto_out_a_bits_user_amba_prot_secure;
  assign auto_buffer_out_a_bits_user_amba_prot_fetch =
    buffer_auto_out_a_bits_user_amba_prot_fetch;
  assign auto_buffer_out_a_bits_mask = buffer_auto_out_a_bits_mask;
  assign auto_buffer_out_a_bits_data = buffer_auto_out_a_bits_data;
  assign auto_buffer_out_a_bits_corrupt = buffer_auto_out_a_bits_corrupt;
  assign auto_buffer_out_b_ready = buffer_auto_out_b_ready;
  assign auto_buffer_out_c_valid = buffer_auto_out_c_valid;
  assign auto_buffer_out_c_bits_opcode = buffer_auto_out_c_bits_opcode;
  assign auto_buffer_out_c_bits_param = buffer_auto_out_c_bits_param;
  assign auto_buffer_out_c_bits_size = buffer_auto_out_c_bits_size;
  assign auto_buffer_out_c_bits_source = buffer_auto_out_c_bits_source;
  assign auto_buffer_out_c_bits_address = buffer_auto_out_c_bits_address;
  assign auto_buffer_out_c_bits_user_amba_prot_bufferable =
    buffer_auto_out_c_bits_user_amba_prot_bufferable;
  assign auto_buffer_out_c_bits_user_amba_prot_modifiable =
    buffer_auto_out_c_bits_user_amba_prot_modifiable;
  assign auto_buffer_out_c_bits_user_amba_prot_readalloc =
    buffer_auto_out_c_bits_user_amba_prot_readalloc;
  assign auto_buffer_out_c_bits_user_amba_prot_writealloc =
    buffer_auto_out_c_bits_user_amba_prot_writealloc;
  assign auto_buffer_out_c_bits_user_amba_prot_privileged =
    buffer_auto_out_c_bits_user_amba_prot_privileged;
  assign auto_buffer_out_c_bits_user_amba_prot_secure =
    buffer_auto_out_c_bits_user_amba_prot_secure;
  assign auto_buffer_out_c_bits_user_amba_prot_fetch =
    buffer_auto_out_c_bits_user_amba_prot_fetch;
  assign auto_buffer_out_c_bits_data = buffer_auto_out_c_bits_data;
  assign auto_buffer_out_c_bits_corrupt = buffer_auto_out_c_bits_corrupt;
  assign auto_buffer_out_d_ready = buffer_auto_out_d_ready;
  assign auto_buffer_out_e_valid = buffer_auto_out_e_valid;
  assign auto_buffer_out_e_bits_sink = buffer_auto_out_e_bits_sink;
  assign auto_broadcast_out_insns_0_valid = broadcast_3_auto_out_insns_0_valid;
  assign auto_broadcast_out_insns_0_iaddr = broadcast_3_auto_out_insns_0_iaddr;
  assign auto_broadcast_out_insns_0_insn = broadcast_3_auto_out_insns_0_insn;
  assign auto_broadcast_out_insns_0_priv = broadcast_3_auto_out_insns_0_priv;
  assign auto_broadcast_out_insns_0_exception = broadcast_3_auto_out_insns_0_exception;
  assign auto_broadcast_out_insns_0_interrupt = broadcast_3_auto_out_insns_0_interrupt;
  assign auto_broadcast_out_insns_0_cause = broadcast_3_auto_out_insns_0_cause;
  assign auto_broadcast_out_insns_0_tval = broadcast_3_auto_out_insns_0_tval;
  assign auto_broadcast_out_time = broadcast_3_auto_out_time;
  assign auto_wfi_out_0 = wfiNodeOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_cease_out_0 = ceaseNodeOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_halt_out_0 = haltNodeOut_0;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_group_0_iretire =
    traceCoreSourceNodeOut_group_0_iretire;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_group_0_iaddr = traceCoreSourceNodeOut_group_0_iaddr;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_group_0_itype = traceCoreSourceNodeOut_group_0_itype;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_group_0_ilastsize =
    traceCoreSourceNodeOut_group_0_ilastsize;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_priv = traceCoreSourceNodeOut_priv;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_tval = traceCoreSourceNodeOut_tval;	// src/main/scala/diplomacy/Nodes.scala:1205:17
  assign auto_trace_core_source_out_cause = traceCoreSourceNodeOut_cause;	// src/main/scala/diplomacy/Nodes.scala:1205:17
endmodule